module top (n0, n1, n2, n3, n4);
    input n0, n1;
    input [63:0] n2;
    input [7:0] n3;
    output [31:0] n4;
    wire n0, n1;
    wire [63:0] n2;
    wire [7:0] n3;
    wire [31:0] n4;
    wire [7:0] n5;
    wire [31:0] n6;
    wire [15:0] n7;
    wire [15:0] n8;
    wire [7:0] n9;
    wire [3:0] n10;
    wire [15:0] n11;
    wire [7:0] n12;
    wire [15:0] n13;
    wire [7:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426;
    or g0(n322 ,n282 ,n291);
    nor g1(n411 ,n340 ,n342);
    nand g2(n401 ,n14[7] ,n400);
    not g3(n100 ,n303);
    dff g4(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n173), .Q(n11[7]));
    not g5(n102 ,n302);
    not g6(n324 ,n7[8]);
    nand g7(n355 ,n14[2] ,n354);
    nand g8(n23 ,n18 ,n16);
    buf g9(n4[26], n4[31]);
    nor g10(n18 ,n11[7] ,n11[6]);
    xnor g11(n425 ,n14[2] ,n353);
    buf g12(n4[16], n4[31]);
    buf g13(n4[30], n4[31]);
    nand g14(n282 ,n5[3] ,n294);
    nor g15(n158 ,n322 ,n137);
    xnor g16(n299 ,n11[2] ,n53);
    nand g17(n131 ,n11[0] ,n107);
    dff g18(.RN(n363), .SN(1'b1), .CK(n0), .D(n424), .Q(n14[3]));
    nor g19(n52 ,n11[1] ,n11[0]);
    nor g20(n419 ,n328 ,n326);
    buf g21(n4[25], n4[31]);
    xnor g22(n4[12] ,n293 ,n6[12]);
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n129), .Q(n8[5]));
    nand g24(n211 ,n319 ,n189);
    nor g25(n146 ,n117 ,n84);
    xnor g26(n4[15] ,n293 ,n6[15]);
    buf g27(n4[24], n4[31]);
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n170), .Q(n11[3]));
    not g29(n337 ,n336);
    not g30(n90 ,n8[3]);
    nand g31(n206 ,n314 ,n189);
    nand g32(n210 ,n318 ,n189);
    or g33(n239 ,n13[15] ,n228);
    xnor g34(n416 ,n7[4] ,n331);
    nand g35(n76 ,n11[14] ,n75);
    xnor g36(n408 ,n7[12] ,n345);
    nor g37(n302 ,n59 ,n61);
    not g38(n328 ,n327);
    nand g39(n225 ,n191 ,n219);
    nand g40(n144 ,n10[1] ,n321);
    xnor g41(n309 ,n11[12] ,n71);
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n138), .Q(n8[0]));
    buf g43(n4[28], n4[31]);
    nor g44(n168 ,n101 ,n133);
    nor g45(n359 ,n14[5] ,n358);
    not g46(n354 ,n353);
    xnor g47(n4[14] ,n293 ,n6[14]);
    nor g48(n44 ,n37 ,n43);
    nor g49(n17 ,n11[1] ,n11[0]);
    nor g50(n149 ,n116 ,n84);
    not g51(n68 ,n67);
    xnor g52(n7[6] ,n2[22] ,n83);
    xnor g53(n421 ,n14[6] ,n360);
    or g54(n243 ,n13[6] ,n228);
    xnor g55(n319 ,n12[2] ,n39);
    xnor g56(n4[9] ,n293 ,n6[9]);
    nor g57(n306 ,n66 ,n68);
    not g58(n91 ,n299);
    nand g59(n387 ,n1 ,n7[9]);
    nor g60(n58 ,n49 ,n57);
    nor g61(n147 ,n111 ,n84);
    not g62(n363 ,n1);
    nand g63(n48 ,n12[6] ,n47);
    not g64(n40 ,n39);
    dff g65(.RN(n363), .SN(1'b1), .CK(n0), .D(n420), .Q(n14[7]));
    xnor g66(n7[3] ,n2[19] ,n79);
    xor g67(n7[13] ,n2[29] ,n2[13]);
    dff g68(.RN(n375), .SN(n391), .CK(n0), .D(n415), .Q(n13[5]));
    nand g69(n270 ,n238 ,n255);
    nand g70(n213 ,n135 ,n194);
    nor g71(n162 ,n93 ,n133);
    not g72(n296 ,n5[5]);
    or g73(n377 ,n363 ,n7[3]);
    dff g74(.RN(n363), .SN(1'b1), .CK(n0), .D(n423), .Q(n14[4]));
    nor g75(n407 ,n347 ,n349);
    xnor g76(n78 ,n2[4] ,n3[4]);
    nand g77(n41 ,n12[2] ,n40);
    dff g78(.RN(n377), .SN(n393), .CK(n0), .D(n417), .Q(n13[3]));
    xnor g79(n413 ,n7[7] ,n336);
    nand g80(n381 ,n1 ,n7[15]);
    not g81(n349 ,n348);
    dff g82(.RN(n378), .SN(n396), .CK(n0), .D(n418), .Q(n13[2]));
    nor g83(n426 ,n354 ,n352);
    nand g84(n390 ,n1 ,n7[6]);
    nor g85(n320 ,n40 ,n38);
    nand g86(n55 ,n11[2] ,n54);
    nor g87(n151 ,n110 ,n84);
    nand g88(n142 ,n8[0] ,n10[0]);
    dff g89(.RN(n369), .SN(n386), .CK(n0), .D(n410), .Q(n13[10]));
    nand g90(n271 ,n234 ,n256);
    nand g91(n207 ,n315 ,n189);
    nor g92(n284 ,n297 ,n5[0]);
    not g93(n75 ,n74);
    dff g94(.RN(n371), .SN(n388), .CK(n0), .D(n412), .Q(n13[8]));
    nand g95(n266 ,n239 ,n251);
    not g96(n228 ,n229);
    nor g97(n28 ,n15 ,n27);
    xnor g98(n7[4] ,n2[20] ,n78);
    nand g99(n403 ,n14[4] ,n402);
    nand g100(n62 ,n11[6] ,n61);
    nand g101(n291 ,n5[1] ,n289);
    not g102(n344 ,n343);
    nand g103(n133 ,n1 ,n3[0]);
    nand g104(n203 ,n12[2] ,n190);
    not g105(n179 ,n178);
    nand g106(n353 ,n14[1] ,n14[0]);
    nand g107(n399 ,n14[6] ,n14[5]);
    not g108(n118 ,n5[3]);
    or g109(n237 ,n13[12] ,n228);
    or g110(n248 ,n13[1] ,n228);
    or g111(n236 ,n13[13] ,n228);
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n149), .Q(n5[2]));
    nand g113(n145 ,n9[2] ,n10[1]);
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n222), .Q(n12[1]));
    dff g115(.RN(n380), .SN(n395), .CK(n0), .D(n7[0]), .Q(n13[0]));
    nor g116(n230 ,n153 ,n229);
    nand g117(n33 ,n12[1] ,n12[0]);
    xnor g118(n417 ,n7[3] ,n329);
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n217), .Q(n12[6]));
    or g120(n375 ,n363 ,n7[5]);
    not g121(n202 ,n201);
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n140), .Q(n5[4]));
    not g123(n325 ,n7[12]);
    nand g124(n278 ,n247 ,n263);
    not g125(n109 ,n12[0]);
    xnor g126(n308 ,n11[11] ,n69);
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n168), .Q(n11[14]));
    not g128(n47 ,n46);
    not g129(n15 ,n11[12]);
    not g130(n99 ,n308);
    nor g131(n232 ,n84 ,n225);
    not g132(n51 ,n11[12]);
    buf g133(n4[23], n4[31]);
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n174), .Q(n11[9]));
    nand g135(n341 ,n7[9] ,n339);
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n169), .Q(n11[11]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n231), .Q(n10[1]));
    not g138(n96 ,n307);
    nor g139(n45 ,n12[5] ,n44);
    not g140(n84 ,n1);
    nand g141(n331 ,n7[3] ,n330);
    nor g142(n400 ,n398 ,n397);
    not g143(n361 ,n360);
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n157), .Q(n11[0]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n132), .Q(n9[0]));
    nand g146(n250 ,n13[8] ,n240);
    nor g147(n161 ,n96 ,n133);
    nand g148(n221 ,n195 ,n209);
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n223), .Q(n12[2]));
    nand g150(n223 ,n203 ,n211);
    not g151(n113 ,n8[4]);
    nand g152(n274 ,n242 ,n265);
    or g153(n235 ,n13[14] ,n228);
    xnor g154(n4[6] ,n293 ,n6[6]);
    or g155(n241 ,n13[8] ,n228);
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n164), .Q(n11[15]));
    not g157(n88 ,n8[5]);
    nand g158(n386 ,n1 ,n7[10]);
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n226), .Q(n10[0]));
    nand g160(n391 ,n1 ,n7[5]);
    nor g161(n333 ,n7[5] ,n332);
    nor g162(n59 ,n11[5] ,n58);
    nand g163(n264 ,n13[6] ,n240);
    nand g164(n176 ,n142 ,n131);
    xnor g165(n315 ,n12[6] ,n46);
    xnor g166(n81 ,n2[1] ,n3[1]);
    nand g167(n268 ,n236 ,n253);
    nand g168(n184 ,n107 ,n181);
    nand g169(n60 ,n11[5] ,n58);
    nand g170(n212 ,n320 ,n189);
    xor g171(n7[14] ,n2[30] ,n2[14]);
    xnor g172(n4[0] ,n293 ,n6[0]);
    dff g173(.RN(n365), .SN(n384), .CK(n0), .D(n408), .Q(n13[12]));
    not g174(n364 ,n14[0]);
    not g175(n104 ,n312);
    nor g176(n66 ,n11[9] ,n65);
    not g177(n54 ,n53);
    nand g178(n397 ,n14[1] ,n14[0]);
    nor g179(n123 ,n119 ,n8[0]);
    dff g180(.RN(n373), .SN(n390), .CK(n0), .D(n414), .Q(n13[6]));
    nor g181(n166 ,n91 ,n133);
    not g182(n56 ,n55);
    nor g183(n192 ,n184 ,n187);
    nor g184(n173 ,n95 ,n133);
    xnor g185(n414 ,n7[6] ,n334);
    nand g186(n262 ,n13[1] ,n240);
    nand g187(n362 ,n14[6] ,n361);
    xnor g188(n4[4] ,n293 ,n6[4]);
    nor g189(n128 ,n88 ,n84);
    nor g190(n189 ,n84 ,n178);
    nand g191(n329 ,n7[2] ,n328);
    nand g192(n261 ,n13[3] ,n240);
    not g193(n297 ,n313);
    not g194(n112 ,n5[4]);
    dff g195(.RN(n363), .SN(1'b1), .CK(n0), .D(n422), .Q(n14[5]));
    xor g196(n7[8] ,n2[24] ,n2[8]);
    xnor g197(n405 ,n7[15] ,n350);
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n175), .Q(n11[5]));
    nand g199(n385 ,n1 ,n7[11]);
    not g200(n93 ,n305);
    nor g201(n148 ,n114 ,n84);
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n130), .Q(n8[2]));
    nand g203(n256 ,n13[10] ,n240);
    not g204(n85 ,n9[0]);
    nand g205(n200 ,n12[3] ,n190);
    not g206(n106 ,n310);
    nor g207(n125 ,n90 ,n84);
    xnor g208(n301 ,n11[4] ,n57);
    nand g209(n46 ,n12[5] ,n44);
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n139), .Q(n9[1]));
    nand g211(n181 ,n3[0] ,n134);
    buf g212(n4[22], n4[31]);
    xnor g213(n418 ,n7[2] ,n327);
    not g214(n95 ,n304);
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n160), .Q(n11[12]));
    nor g216(n127 ,n86 ,n84);
    xnor g217(n286 ,n11[0] ,n12[0]);
    not g218(n103 ,n300);
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n150), .Q(n5[5]));
    nor g220(n141 ,n115 ,n84);
    nand g221(n199 ,n12[1] ,n190);
    buf g222(n4[17], n4[31]);
    or g223(n249 ,n13[4] ,n228);
    nor g224(n130 ,n119 ,n84);
    nand g225(n53 ,n11[1] ,n11[0]);
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n127), .Q(n9[3]));
    nand g227(n253 ,n13[13] ,n240);
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n166), .Q(n11[2]));
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n278), .Q(n6[2]));
    buf g230(n4[20], n4[31]);
    nor g231(n177 ,n122 ,n121);
    xnor g232(n290 ,n286 ,n8[0]);
    not g233(n105 ,n301);
    or g234(n215 ,n191 ,n201);
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n268), .Q(n6[13]));
    buf g236(n4[27], n4[31]);
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n258), .Q(n6[0]));
    nand g238(n279 ,n248 ,n262);
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n270), .Q(n6[11]));
    nor g240(n422 ,n359 ,n361);
    dff g241(.RN(n366), .SN(n382), .CK(n0), .D(n406), .Q(n13[14]));
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n273), .Q(n6[12]));
    xnor g243(n4[5] ,n293 ,n6[5]);
    nor g244(n16 ,n11[5] ,n11[4]);
    not g245(n49 ,n11[4]);
    nor g246(n29 ,n11[13] ,n28);
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n154), .Q(n5[0]));
    or g248(n31 ,n12[5] ,n12[4]);
    nor g249(n73 ,n11[13] ,n72);
    nor g250(n240 ,n84 ,n229);
    nand g251(n383 ,n1 ,n7[13]);
    buf g252(n4[19], n4[31]);
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n224), .Q(n12[3]));
    nor g254(n310 ,n73 ,n75);
    nand g255(n204 ,n12[0] ,n190);
    dff g256(.RN(n372), .SN(n381), .CK(n0), .D(n405), .Q(n13[15]));
    or g257(n380 ,n363 ,n7[0]);
    nand g258(n122 ,n8[5] ,n113);
    nor g259(n129 ,n113 ,n84);
    xnor g260(n406 ,n7[14] ,n348);
    nand g261(n188 ,n136 ,n177);
    nand g262(n272 ,n245 ,n257);
    nand g263(n252 ,n13[14] ,n240);
    not g264(n37 ,n12[4]);
    nand g265(n224 ,n200 ,n210);
    nand g266(n281 ,n5[7] ,n295);
    nand g267(n255 ,n13[11] ,n240);
    xnor g268(n303 ,n11[6] ,n60);
    nand g269(n69 ,n11[10] ,n68);
    nor g270(n124 ,n90 ,n8[2]);
    not g271(n101 ,n311);
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n275), .Q(n6[6]));
    nand g273(n193 ,n109 ,n189);
    not g274(n342 ,n341);
    not g275(n295 ,n5[6]);
    nor g276(n160 ,n94 ,n133);
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n151), .Q(n5[6]));
    nor g278(n289 ,n281 ,n288);
    xnor g279(n7[1] ,n81 ,n2[17]);
    or g280(n365 ,n363 ,n7[12]);
    nand g281(n327 ,n7[1] ,n404);
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n271), .Q(n6[10]));
    or g283(n371 ,n363 ,n7[8]);
    nand g284(n343 ,n7[10] ,n342);
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n165), .Q(n11[4]));
    xnor g286(n4[7] ,n293 ,n6[7]);
    or g287(n247 ,n13[2] ,n228);
    or g288(n234 ,n13[10] ,n228);
    nand g289(n67 ,n11[9] ,n65);
    nor g290(n150 ,n112 ,n84);
    nand g291(n36 ,n12[3] ,n35);
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n272), .Q(n6[9]));
    xnor g293(n312 ,n76 ,n11[15]);
    nand g294(n334 ,n7[5] ,n332);
    nand g295(n208 ,n316 ,n189);
    dff g296(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n269), .Q(n6[8]));
    xnor g297(n7[5] ,n80 ,n2[21]);
    nand g298(n71 ,n11[11] ,n70);
    nand g299(n276 ,n244 ,n259);
    nor g300(n139 ,n85 ,n84);
    dff g301(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n220), .Q(n12[5]));
    nor g302(n352 ,n14[1] ,n14[0]);
    dff g303(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n147), .Q(n5[1]));
    nor g304(n283 ,n296 ,n5[4]);
    nor g305(n167 ,n97 ,n133);
    not g306(n63 ,n62);
    nor g307(n332 ,n323 ,n331);
    xnor g308(n83 ,n2[6] ,n3[6]);
    nor g309(n340 ,n7[9] ,n339);
    nand g310(n396 ,n1 ,n7[2]);
    or g311(n376 ,n363 ,n7[4]);
    nand g312(n153 ,n1 ,n13[0]);
    dff g313(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n172), .Q(n11[13]));
    nand g314(n57 ,n11[3] ,n56);
    nand g315(n275 ,n243 ,n264);
    nand g316(n194 ,n185 ,n183);
    xnor g317(n307 ,n11[10] ,n67);
    nand g318(n26 ,n17 ,n25);
    xnor g319(n285 ,n2[0] ,n3[0]);
    nand g320(n388 ,n1 ,n7[8]);
    nand g321(n345 ,n7[11] ,n344);
    not g322(n111 ,n5[0]);
    nor g323(n164 ,n104 ,n133);
    xnor g324(n79 ,n2[3] ,n3[3]);
    nand g325(n321 ,n21 ,n29);
    xnor g326(n410 ,n7[10] ,n341);
    not g327(n294 ,n5[2]);
    nand g328(n43 ,n12[3] ,n42);
    nand g329(n209 ,n317 ,n189);
    dff g330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n146), .Q(n8[7]));
    or g331(n20 ,n11[3] ,n11[2]);
    nand g332(n121 ,n8[7] ,n117);
    xor g333(n7[9] ,n2[25] ,n2[9]);
    or g334(n370 ,n363 ,n7[9]);
    or g335(n32 ,n12[7] ,n12[6]);
    not g336(n154 ,n153);
    nand g337(n382 ,n1 ,n7[14]);
    dff g338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n221), .Q(n12[4]));
    xnor g339(n4[3] ,n293 ,n6[3]);
    nor g340(n65 ,n50 ,n64);
    nand g341(n74 ,n11[13] ,n72);
    or g342(n378 ,n363 ,n7[2]);
    not g343(n30 ,n12[2]);
    xnor g344(n4[8] ,n293 ,n6[8]);
    or g345(n238 ,n13[11] ,n228);
    xnor g346(n82 ,n2[2] ,n3[2]);
    nand g347(n197 ,n12[7] ,n190);
    nand g348(n198 ,n12[6] ,n190);
    nand g349(n251 ,n13[15] ,n240);
    nand g350(n277 ,n246 ,n261);
    or g351(n369 ,n363 ,n7[10]);
    xnor g352(n317 ,n12[4] ,n43);
    nand g353(n64 ,n11[7] ,n63);
    nor g354(n126 ,n87 ,n84);
    nor g355(n136 ,n107 ,n10[1]);
    xnor g356(n409 ,n7[11] ,n343);
    nor g357(n233 ,n13[0] ,n228);
    nand g358(n273 ,n237 ,n254);
    dff g359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n274), .Q(n6[7]));
    not g360(n89 ,n9[1]);
    nand g361(n205 ,n9[0] ,n189);
    nor g362(n358 ,n351 ,n357);
    nand g363(n393 ,n1 ,n7[3]);
    not g364(n116 ,n5[1]);
    not g365(n219 ,n218);
    nand g366(n143 ,n9[0] ,n9[1]);
    nand g367(n263 ,n13[2] ,n240);
    buf g368(n4[21], n4[31]);
    nor g369(n347 ,n7[13] ,n346);
    nor g370(n187 ,n145 ,n171);
    nand g371(n348 ,n7[13] ,n346);
    nand g372(n196 ,n12[5] ,n190);
    nand g373(n214 ,n204 ,n193);
    nor g374(n346 ,n325 ,n345);
    dff g375(.RN(n363), .SN(1'b1), .CK(n0), .D(n421), .Q(n14[6]));
    or g376(n242 ,n13[7] ,n228);
    or g377(n258 ,n233 ,n230);
    xnor g378(n304 ,n11[7] ,n62);
    nand g379(n357 ,n14[3] ,n356);
    nor g380(n163 ,n100 ,n133);
    nor g381(n21 ,n11[15] ,n11[14]);
    dff g382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n167), .Q(n11[1]));
    not g383(n351 ,n14[4]);
    xnor g384(n318 ,n12[3] ,n41);
    nand g385(n338 ,n7[7] ,n337);
    xnor g386(n305 ,n11[8] ,n64);
    nor g387(n140 ,n118 ,n84);
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n120), .Q(n9[2]));
    xor g389(n7[11] ,n2[27] ,n2[11]);
    nand g390(n336 ,n7[6] ,n335);
    not g391(n132 ,n133);
    nor g392(n72 ,n51 ,n71);
    xnor g393(n293 ,n292 ,n290);
    dff g394(.RN(n374), .SN(n389), .CK(n0), .D(n413), .Q(n13[7]));
    not g395(n87 ,n8[2]);
    xnor g396(n412 ,n7[8] ,n338);
    nand g397(n350 ,n7[14] ,n349);
    not g398(n70 ,n69);
    xnor g399(n4[13] ,n293 ,n6[13]);
    or g400(n245 ,n13[9] ,n228);
    not g401(n114 ,n5[2]);
    nor g402(n27 ,n20 ,n26);
    not g403(n94 ,n309);
    dff g404(.RN(n363), .SN(1'b1), .CK(n0), .D(n425), .Q(n14[2]));
    not g405(n117 ,n8[6]);
    not g406(n402 ,n401);
    nor g407(n174 ,n98 ,n133);
    nand g408(n191 ,n135 ,n159);
    xnor g409(n7[2] ,n2[18] ,n82);
    dff g410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n267), .Q(n6[14]));
    nand g411(n218 ,n186 ,n202);
    dff g412(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n126), .Q(n8[3]));
    xnor g413(n424 ,n14[3] ,n355);
    nand g414(n389 ,n1 ,n7[7]);
    dff g415(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n161), .Q(n11[10]));
    nand g416(n288 ,n284 ,n283);
    nor g417(n135 ,n84 ,n10[2]);
    xnor g418(n311 ,n11[14] ,n74);
    nand g419(n280 ,n249 ,n260);
    not g420(n97 ,n298);
    dff g421(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n141), .Q(n5[7]));
    or g422(n373 ,n363 ,n7[6]);
    not g423(n50 ,n11[8]);
    or g424(n367 ,n363 ,n7[13]);
    nor g425(n339 ,n324 ,n338);
    nor g426(n157 ,n11[0] ,n133);
    nor g427(n34 ,n32 ,n31);
    xnor g428(n4[11] ,n293 ,n6[11]);
    nor g429(n415 ,n333 ,n335);
    nor g430(n165 ,n105 ,n133);
    nand g431(n180 ,n322 ,n134);
    xnor g432(n4[1] ,n293 ,n6[1]);
    xnor g433(n77 ,n2[7] ,n3[7]);
    nand g434(n156 ,n123 ,n124);
    nor g435(n25 ,n24 ,n23);
    dff g436(.RN(n367), .SN(n383), .CK(n0), .D(n407), .Q(n13[13]));
    or g437(n244 ,n13[5] ,n228);
    or g438(n159 ,n107 ,n144);
    dff g439(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n128), .Q(n8[6]));
    xnor g440(n314 ,n12[7] ,n48);
    dff g441(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n216), .Q(n12[7]));
    not g442(n107 ,n10[0]);
    dff g443(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n232), .Q(n10[2]));
    nor g444(n175 ,n102 ,n133);
    dff g445(.RN(n376), .SN(n392), .CK(n0), .D(n416), .Q(n13[4]));
    not g446(n108 ,n8[0]);
    not g447(n115 ,n5[6]);
    dff g448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n214), .Q(n12[0]));
    not g449(n356 ,n355);
    dff g450(.RN(n363), .SN(1'b1), .CK(n0), .D(n426), .Q(n14[1]));
    buf g451(n4[18], n4[31]);
    xnor g452(n4[2] ,n293 ,n6[2]);
    xnor g453(n4[10] ,n293 ,n6[10]);
    nand g454(n254 ,n13[12] ,n240);
    dff g455(.RN(n379), .SN(n394), .CK(n0), .D(n419), .Q(n13[1]));
    nor g456(n138 ,n84 ,n92);
    not g457(n155 ,n143);
    or g458(n366 ,n363 ,n7[14]);
    dff g459(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n148), .Q(n5[3]));
    nor g460(n22 ,n11[11] ,n11[10]);
    dff g461(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n125), .Q(n8[4]));
    not g462(n42 ,n41);
    nor g463(n190 ,n84 ,n179);
    nor g464(n227 ,n10[1] ,n218);
    xor g465(n292 ,n287 ,n322);
    nand g466(n35 ,n30 ,n33);
    nor g467(n120 ,n89 ,n84);
    nor g468(n169 ,n99 ,n133);
    xnor g469(n7[7] ,n2[23] ,n77);
    xor g470(n7[10] ,n2[26] ,n2[10]);
    nor g471(n201 ,n156 ,n188);
    not g472(n86 ,n9[2]);
    xnor g473(n423 ,n14[4] ,n357);
    nand g474(n360 ,n14[5] ,n358);
    nor g475(n183 ,n158 ,n182);
    nand g476(n222 ,n199 ,n212);
    nor g477(n226 ,n192 ,n215);
    nor g478(n231 ,n191 ,n227);
    nor g479(n170 ,n103 ,n133);
    nor g480(n152 ,n108 ,n84);
    buf g481(n4[29], n4[31]);
    nor g482(n134 ,n10[0] ,n10[1]);
    xnor g483(n420 ,n362 ,n14[7]);
    not g484(n92 ,n2[0]);
    xor g485(n7[12] ,n2[28] ,n2[12]);
    not g486(n137 ,n136);
    not g487(n330 ,n329);
    nand g488(n265 ,n13[7] ,n240);
    nor g489(n38 ,n12[1] ,n12[0]);
    dff g490(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n279), .Q(n6[1]));
    dff g491(.RN(n368), .SN(n385), .CK(n0), .D(n409), .Q(n13[11]));
    dff g492(.RN(n370), .SN(n387), .CK(n0), .D(n411), .Q(n13[9]));
    nand g493(n195 ,n12[4] ,n190);
    nor g494(n316 ,n45 ,n47);
    or g495(n368 ,n363 ,n7[11]);
    not g496(n61 ,n60);
    dff g497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n152), .Q(n8[1]));
    nand g498(n178 ,n10[2] ,n134);
    nand g499(n269 ,n241 ,n250);
    nand g500(n216 ,n197 ,n206);
    nor g501(n19 ,n11[9] ,n11[8]);
    nand g502(n185 ,n10[1] ,n176);
    nor g503(n298 ,n54 ,n52);
    nand g504(n259 ,n13[5] ,n240);
    nand g505(n394 ,n1 ,n7[1]);
    not g506(n119 ,n8[1]);
    not g507(n98 ,n306);
    or g508(n372 ,n363 ,n7[15]);
    xnor g509(n7[0] ,n2[16] ,n285);
    dff g510(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n277), .Q(n6[3]));
    dff g511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n229), .Q(n6[16]));
    nand g512(n395 ,n1 ,n7[0]);
    nand g513(n257 ,n13[9] ,n240);
    nand g514(n171 ,n9[3] ,n155);
    xnor g515(n4[31] ,n6[16] ,n293);
    not g516(n182 ,n181);
    or g517(n246 ,n13[3] ,n228);
    nand g518(n39 ,n12[1] ,n12[0]);
    not g519(n110 ,n5[5]);
    or g520(n379 ,n363 ,n7[1]);
    nand g521(n229 ,n205 ,n213);
    nand g522(n186 ,n10[2] ,n180);
    xnor g523(n287 ,n9[0] ,n10[0]);
    not g524(n335 ,n334);
    dff g525(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n162), .Q(n11[8]));
    nand g526(n260 ,n13[4] ,n240);
    nand g527(n24 ,n22 ,n19);
    dff g528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n280), .Q(n6[4]));
    nand g529(n392 ,n1 ,n7[4]);
    nand g530(n384 ,n1 ,n7[12]);
    xor g531(n7[15] ,n2[31] ,n2[15]);
    nand g532(n313 ,n36 ,n34);
    dff g533(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n276), .Q(n6[5]));
    dff g534(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n266), .Q(n6[15]));
    xnor g535(n300 ,n11[3] ,n55);
    nor g536(n326 ,n7[1] ,n404);
    dff g537(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n163), .Q(n11[6]));
    nand g538(n267 ,n235 ,n252);
    nand g539(n217 ,n198 ,n207);
    nor g540(n172 ,n106 ,n133);
    xnor g541(n80 ,n2[5] ,n3[5]);
    nand g542(n220 ,n196 ,n208);
    not g543(n323 ,n7[4]);
    nor g544(n404 ,n399 ,n403);
    or g545(n374 ,n363 ,n7[7]);
    nand g546(n398 ,n14[3] ,n14[2]);
    dff g547(.RN(n363), .SN(1'b1), .CK(n0), .D(n364), .Q(n14[0]));
endmodule
