module top (n0, n1, n4, n5, n2, n3, n6, n7, n12, n14, n15, n8, n9, n10, n11, n13);
    input n0, n1, n2, n3;
    input [7:0] n4, n5;
    output [2:0] n6, n7, n8, n9, n10, n11;
    output [7:0] n12, n13;
    output n14, n15;
    wire n0, n1, n2, n3;
    wire [7:0] n4, n5;
    wire [2:0] n6, n7, n8, n9, n10, n11;
    wire [7:0] n12, n13;
    wire n14, n15;
    wire [31:0] n16;
    wire n17, n18, n19, n20, n21, n22, n23, n24;
    wire n25, n26, n27, n28, n29, n30, n31, n32;
    wire n33, n34, n35, n36, n37, n38, n39, n40;
    wire n41, n42, n43, n44, n45, n46, n47, n48;
    wire n49, n50, n51, n52, n53, n54, n55, n56;
    wire n57, n58, n59, n60, n61, n62, n63, n64;
    wire n65, n66, n67, n68, n69, n70, n71, n72;
    wire n73, n74, n75, n76, n77, n78, n79, n80;
    wire n81, n82, n83, n84, n85, n86, n87, n88;
    wire n89, n90, n91, n92, n93, n94, n95, n96;
    wire n97, n98, n99, n100, n101, n102, n103, n104;
    wire n105, n106, n107, n108, n109, n110, n111, n112;
    wire n113, n114, n115, n116, n117, n118, n119, n120;
    wire n121, n122, n123, n124, n125, n126, n127, n128;
    wire n129, n130, n131, n132, n133, n134, n135, n136;
    wire n137, n138, n139, n140, n141, n142, n143, n144;
    wire n145, n146, n147, n148, n149, n150, n151, n152;
    wire n153, n154, n155, n156, n157, n158, n159, n160;
    wire n161, n162, n163, n164, n165, n166, n167, n168;
    wire n169, n170, n171, n172, n173, n174, n175, n176;
    wire n177, n178, n179, n180, n181, n182, n183, n184;
    wire n185, n186, n187, n188, n189, n190, n191, n192;
    wire n193, n194, n195, n196, n197, n198, n199, n200;
    wire n201, n202, n203, n204, n205, n206, n207, n208;
    wire n209, n210, n211, n212, n213;
    dff g0(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n92), .Q(n13[1]));
    not g1(n45 ,n3);
    nand g2(n139 ,n127 ,n129);
    nand g3(n126 ,n4[4] ,n107);
    nand g4(n163 ,n206 ,n142);
    nor g5(n84 ,n42 ,n37);
    nor g6(n199 ,n122 ,n195);
    not g7(n30 ,n29);
    dff g8(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n103), .Q(n12[6]));
    dff g9(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n141), .Q(n14));
    not g10(n109 ,n108);
    nor g11(n178 ,n37 ,n147);
    nand g12(n73 ,n6[1] ,n6[2]);
    nor g13(n88 ,n54 ,n37);
    nor g14(n141 ,n60 ,n135);
    nand g15(n61 ,n7[2] ,n37);
    nand g16(n58 ,n7[0] ,n37);
    nand g17(n63 ,n6[2] ,n1);
    nand g18(n150 ,n50 ,n142);
    nor g19(n101 ,n69 ,n67);
    not g20(n40 ,n4[3]);
    nand g21(n165 ,n209 ,n142);
    nand g22(n111 ,n6[1] ,n68);
    nor g23(n90 ,n51 ,n37);
    nor g24(n130 ,n45 ,n98);
    nor g25(n86 ,n37 ,n40);
    nor g26(n175 ,n3 ,n171);
    not g27(n124 ,n123);
    nor g28(n94 ,n41 ,n37);
    nand g29(n203 ,n61 ,n201);
    nor g30(n117 ,n79 ,n106);
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n91), .Q(n13[2]));
    nand g32(n162 ,n207 ,n142);
    nand g33(n75 ,n6[2] ,n48);
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n86), .Q(n13[3]));
    nand g35(n156 ,n16[3] ,n146);
    nor g36(n147 ,n117 ,n144);
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n96), .Q(n13[5]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n85), .Q(n11[0]));
    nor g39(n83 ,n55 ,n37);
    nand g40(n169 ,n210 ,n142);
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n101), .Q(n12[2]));
    or g42(n148 ,n138 ,n143);
    nor g43(n102 ,n65 ,n75);
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n184), .Q(n16[1]));
    xnor g45(n211 ,n16[8] ,n34);
    nand g46(n118 ,n47 ,n108);
    nor g47(n125 ,n37 ,n109);
    nor g48(n187 ,n63 ,n186);
    xnor g49(n208 ,n16[5] ,n29);
    not g50(n105 ,n104);
    nand g51(n145 ,n213 ,n136);
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n180), .Q(n16[5]));
    nand g53(n160 ,n212 ,n142);
    nor g54(n119 ,n37 ,n105);
    nand g55(n172 ,n153 ,n169);
    nand g56(n19 ,n16[9] ,n16[8]);
    not g57(n46 ,n4[2]);
    nand g58(n143 ,n128 ,n137);
    or g59(n100 ,n73 ,n77);
    not g60(n66 ,n65);
    nor g61(n134 ,n5[2] ,n116);
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n66), .Q(n8[0]));
    not g63(n50 ,n16[0]);
    not g64(n22 ,n16[2]);
    xnor g65(n205 ,n16[2] ,n24);
    nand g66(n198 ,n62 ,n192);
    nor g67(n115 ,n59 ,n97);
    not g68(n136 ,n135);
    nor g69(n59 ,n38 ,n5[5]);
    nor g70(n103 ,n73 ,n65);
    nand g71(n69 ,n6[1] ,n1);
    nand g72(n174 ,n164 ,n150);
    nand g73(n138 ,n1 ,n129);
    nor g74(n85 ,n43 ,n37);
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n174), .Q(n16[0]));
    nand g76(n164 ,n16[0] ,n146);
    not g77(n44 ,n4[0]);
    nand g78(n127 ,n4[1] ,n104);
    nand g79(n196 ,n189 ,n191);
    nor g80(n173 ,n133 ,n149);
    nor g81(n210 ,n33 ,n35);
    nand g82(n176 ,n151 ,n160);
    nand g83(n190 ,n100 ,n186);
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n175), .Q(n15));
    not g85(n38 ,n6[0]);
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n99), .Q(n12[3]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n183), .Q(n16[2]));
    nor g88(n213 ,n18 ,n21);
    nand g89(n149 ,n121 ,n140);
    nor g90(n206 ,n26 ,n28);
    nand g91(n18 ,n16[6] ,n16[5]);
    nand g92(n106 ,n6[2] ,n71);
    not g93(n76 ,n75);
    nand g94(n62 ,n7[1] ,n37);
    nor g95(n93 ,n37 ,n44);
    nand g96(n95 ,n15 ,n1);
    nand g97(n180 ,n159 ,n161);
    not g98(n53 ,n10[1]);
    nor g99(n60 ,n14 ,n213);
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n90), .Q(n13[4]));
    nor g101(n133 ,n5[0] ,n118);
    xnor g102(n207 ,n16[4] ,n27);
    nand g103(n129 ,n5[0] ,n108);
    nand g104(n177 ,n152 ,n168);
    nor g105(n79 ,n4[5] ,n4[4]);
    nand g106(n182 ,n156 ,n163);
    nand g107(n67 ,n6[0] ,n49);
    nand g108(n166 ,n204 ,n142);
    buf g109(n153 ,n145);
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n179), .Q(n16[6]));
    nor g111(n91 ,n37 ,n46);
    nor g112(n71 ,n6[0] ,n6[1]);
    nand g113(n170 ,n205 ,n142);
    nor g114(n135 ,n110 ,n125);
    nor g115(n20 ,n19 ,n17);
    nor g116(n142 ,n213 ,n135);
    buf g117(n13[6], n8[0]);
    nand g118(n200 ,n58 ,n197);
    not g119(n43 ,n10[0]);
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n196), .Q(n6[0]));
    not g121(n52 ,n8[2]);
    not g122(n48 ,n6[1]);
    nand g123(n161 ,n208 ,n142);
    not g124(n107 ,n106);
    buf g125(n12[7], 1'b0);
    xnor g126(n209 ,n16[6] ,n31);
    nor g127(n17 ,n16[4] ,n16[3]);
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n83), .Q(n11[2]));
    nand g129(n65 ,n6[0] ,n1);
    or g130(n116 ,n4[3] ,n111);
    not g131(n55 ,n10[2]);
    buf g132(n154 ,n145);
    nand g133(n167 ,n95 ,n145);
    buf g134(n152 ,n145);
    not g135(n47 ,n5[1]);
    nor g136(n140 ,n134 ,n120);
    nor g137(n77 ,n6[0] ,n5[3]);
    not g138(n72 ,n71);
    not g139(n193 ,n192);
    nand g140(n179 ,n154 ,n165);
    xnor g141(n212 ,n16[9] ,n36);
    not g142(n54 ,n8[0]);
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n84), .Q(n10[1]));
    nand g144(n36 ,n16[8] ,n35);
    or g145(n122 ,n37 ,n113);
    nor g146(n192 ,n178 ,n188);
    nor g147(n97 ,n5[4] ,n78);
    not g148(n64 ,n63);
    nand g149(n74 ,n6[1] ,n38);
    not g150(n146 ,n145);
    xor g151(n204 ,n16[1] ,n16[0]);
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n177), .Q(n16[8]));
    nand g153(n27 ,n16[3] ,n25);
    nand g154(n31 ,n16[5] ,n30);
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n94), .Q(n10[2]));
    not g156(n37 ,n1);
    nor g157(n201 ,n187 ,n199);
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n202), .Q(n6[2]));
    not g159(n202 ,n201);
    nand g160(n123 ,n39 ,n104);
    nor g161(n92 ,n37 ,n39);
    not g162(n42 ,n9[1]);
    nor g163(n33 ,n16[7] ,n32);
    not g164(n41 ,n9[2]);
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n70), .Q(n8[1]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n89), .Q(n9[1]));
    not g167(n197 ,n196);
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n182), .Q(n16[3]));
    nor g169(n81 ,n57 ,n37);
    nor g170(n110 ,n63 ,n74);
    nand g171(n184 ,n158 ,n166);
    nand g172(n183 ,n157 ,n170);
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n82), .Q(n11[1]));
    not g174(n68 ,n67);
    nor g175(n186 ,n132 ,n185);
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n88), .Q(n9[0]));
    nand g177(n98 ,n6[0] ,n76);
    nand g178(n181 ,n155 ,n162);
    nor g179(n194 ,n139 ,n190);
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n203), .Q(n7[2]));
    nand g181(n21 ,n16[7] ,n20);
    nand g182(n29 ,n16[4] ,n28);
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n200), .Q(n7[0]));
    not g184(n80 ,n79);
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n93), .Q(n13[0]));
    buf g186(n151 ,n145);
    not g187(n56 ,n8[1]);
    nor g188(n188 ,n69 ,n186);
    nor g189(n87 ,n52 ,n37);
    or g190(n189 ,n65 ,n186);
    nand g191(n168 ,n211 ,n142);
    nand g192(n24 ,n16[1] ,n16[0]);
    nand g193(n157 ,n16[2] ,n146);
    not g194(n114 ,n113);
    nor g195(n113 ,n6[2] ,n72);
    not g196(n171 ,n167);
    nor g197(n99 ,n63 ,n72);
    or g198(n144 ,n130 ,n139);
    nor g199(n104 ,n6[2] ,n74);
    nand g200(n195 ,n126 ,n194);
    not g201(n112 ,n111);
    nand g202(n128 ,n4[3] ,n112);
    buf g203(n13[7], n8[1]);
    not g204(n49 ,n6[2]);
    nand g205(n34 ,n16[7] ,n32);
    not g206(n70 ,n69);
    dff g207(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n176), .Q(n16[9]));
    not g208(n96 ,n95);
    or g209(n191 ,n148 ,n190);
    nor g210(n32 ,n23 ,n31);
    nand g211(n155 ,n16[4] ,n146);
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n193), .Q(n6[1]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n110), .Q(n12[5]));
    nor g214(n120 ,n80 ,n106);
    not g215(n51 ,n14);
    not g216(n28 ,n27);
    not g217(n35 ,n34);
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n81), .Q(n10[0]));
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n119), .Q(n12[1]));
    nand g220(n185 ,n131 ,n173);
    not g221(n57 ,n9[0]);
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n125), .Q(n12[0]));
    or g223(n131 ,n73 ,n115);
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n172), .Q(n16[7]));
    nor g225(n26 ,n16[3] ,n25);
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n181), .Q(n16[4]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n87), .Q(n9[2]));
    nand g228(n158 ,n16[1] ,n146);
    not g229(n78 ,n77);
    or g230(n121 ,n4[0] ,n114);
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n198), .Q(n7[1]));
    nor g232(n82 ,n53 ,n37);
    nor g233(n132 ,n4[2] ,n123);
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n102), .Q(n12[4]));
    not g235(n39 ,n4[1]);
    not g236(n23 ,n16[6]);
    nor g237(n89 ,n56 ,n37);
    nor g238(n25 ,n22 ,n24);
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n64), .Q(n8[2]));
    nor g240(n137 ,n130 ,n124);
    buf g241(n159 ,n145);
    nor g242(n108 ,n6[1] ,n67);
endmodule
