module top (n0, n1, n2);
    input n0, n1;
    output n2;
    wire n0, n1;
    wire n2;
    wire [31:0] n3;
    wire [31:0] n4;
    wire [7:0] n5;
    wire n6, n7, n8, n9, n10, n11, n12, n13;
    wire n14, n15, n16, n17, n18, n19, n20, n21;
    wire n22, n23, n24, n25, n26, n27, n28, n29;
    wire n30, n31, n32, n33, n34, n35, n36, n37;
    wire n38, n39, n40, n41, n42, n43, n44, n45;
    wire n46, n47, n48, n49, n50, n51, n52, n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171, n172, n173;
    wire n174, n175, n176, n177, n178, n179, n180, n181;
    wire n182, n183, n184, n185, n186, n187, n188, n189;
    wire n190, n191, n192, n193, n194, n195, n196, n197;
    wire n198, n199, n200, n201, n202, n203, n204, n205;
    wire n206, n207, n208, n209, n210, n211, n212, n213;
    wire n214, n215, n216, n217, n218, n219, n220, n221;
    wire n222, n223, n224, n225, n226, n227, n228, n229;
    wire n230, n231, n232, n233, n234, n235, n236, n237;
    wire n238, n239, n240, n241, n242, n243, n244, n245;
    wire n246, n247, n248, n249, n250, n251, n252, n253;
    wire n254, n255, n256, n257, n258, n259, n260, n261;
    wire n262, n263, n264, n265, n266, n267, n268, n269;
    wire n270, n271, n272, n273, n274, n275, n276, n277;
    wire n278, n279, n280, n281, n282, n283, n284, n285;
    nor g0(n198 ,n168 ,n178);
    nand g1(n68 ,n3[2] ,n67);
    xnor g2(n247 ,n4[16] ,n36);
    dff g3(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n180), .Q(n269));
    nand g4(n42 ,n4[19] ,n41);
    nand g5(n14 ,n4[4] ,n13);
    nand g6(n226 ,n207 ,n206);
    nor g7(n117 ,n102 ,n3[2]);
    xnor g8(n260 ,n54 ,n4[26]);
    xnor g9(n241 ,n24 ,n4[10]);
    nand g10(n224 ,n265 ,n222);
    dff g11(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n205), .Q(n4[3]));
    nand g12(n30 ,n4[12] ,n29);
    nand g13(n223 ,n266 ,n222);
    nand g14(n123 ,n106 ,n104);
    dff g15(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n198), .Q(n4[9]));
    nand g16(n218 ,n3[2] ,n179);
    nand g17(n58 ,n4[27] ,n57);
    nor g18(n208 ,n160 ,n178);
    not g19(n146 ,n256);
    or g20(n174 ,n268 ,n259);
    nor g21(n179 ,n269 ,n176);
    not g22(n41 ,n40);
    nor g23(n215 ,n146 ,n178);
    nand g24(n39 ,n4[16] ,n37);
    nor g25(n285 ,n284 ,n283);
    not g26(n152 ,n245);
    nand g27(n66 ,n3[1] ,n3[0]);
    nor g28(n135 ,n117 ,n132);
    xnor g29(n244 ,n30 ,n4[13]);
    dff g30(.RN(n270), .SN(1'b1), .CK(n0), .D(n4[0]), .Q(n5[0]));
    or g31(n268 ,n4[31] ,n142);
    nor g32(n104 ,n4[16] ,n4[15]);
    nand g33(n141 ,n128 ,n140);
    nand g34(n18 ,n4[6] ,n17);
    nor g35(n110 ,n4[20] ,n4[19]);
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n212), .Q(n4[27]));
    nor g37(n187 ,n171 ,n178);
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n191), .Q(n4[15]));
    nor g39(n200 ,n164 ,n178);
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n189), .Q(n4[17]));
    nand g41(n32 ,n4[13] ,n31);
    nor g42(n78 ,n4[26] ,n4[25]);
    not g43(n47 ,n46);
    xnor g44(n261 ,n56 ,n4[27]);
    nand g45(n22 ,n4[8] ,n21);
    nor g46(n188 ,n148 ,n178);
    not g47(n149 ,n251);
    nand g48(n122 ,n105 ,n111);
    nor g49(n271 ,n5[4] ,n5[6]);
    nand g50(n20 ,n4[7] ,n19);
    nand g51(n221 ,n267 ,n182);
    nand g52(n178 ,n174 ,n175);
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n226), .Q(n2));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n185), .Q(n4[21]));
    nand g55(n16 ,n4[5] ,n15);
    not g56(n171 ,n250);
    dff g57(.RN(n270), .SN(1'b1), .CK(n0), .D(n4[5]), .Q(n5[5]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n193), .Q(n4[13]));
    nor g59(n109 ,n4[6] ,n4[5]);
    not g60(n177 ,n178);
    nor g61(n129 ,n4[4] ,n124);
    nand g62(n9 ,n4[17] ,n4[16]);
    nor g63(n120 ,n4[12] ,n4[11]);
    or g64(n137 ,n115 ,n136);
    not g65(n57 ,n56);
    or g66(n132 ,n116 ,n130);
    not g67(n67 ,n66);
    not g68(n153 ,n254);
    not g69(n25 ,n24);
    nand g70(n206 ,n268 ,n177);
    not g71(n157 ,n244);
    not g72(n172 ,n241);
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n214), .Q(n4[23]));
    nand g74(n181 ,n269 ,n175);
    nand g75(n56 ,n4[26] ,n55);
    nor g76(n205 ,n158 ,n178);
    nand g77(n231 ,n219 ,n225);
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n186), .Q(n4[20]));
    xnor g79(n234 ,n4[3] ,n10);
    not g80(n43 ,n42);
    not g81(n160 ,n258);
    xnor g82(n246 ,n34 ,n4[15]);
    nor g83(n142 ,n138 ,n141);
    not g84(n33 ,n32);
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n220), .Q(n4[28]));
    nand g86(n12 ,n4[3] ,n11);
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n208), .Q(n4[31]));
    not g88(n45 ,n44);
    nand g89(n133 ,n109 ,n129);
    nand g90(n60 ,n4[28] ,n59);
    nand g91(n48 ,n4[22] ,n47);
    not g92(n63 ,n62);
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n202), .Q(n4[4]));
    nand g94(n24 ,n4[9] ,n23);
    xnor g95(n243 ,n28 ,n4[12]);
    nor g96(n278 ,n4[5] ,n4[3]);
    not g97(n154 ,n253);
    not g98(n222 ,n221);
    nor g99(n213 ,n156 ,n178);
    nand g100(n40 ,n4[18] ,n38);
    not g101(n168 ,n240);
    nor g102(n91 ,n85 ,n84);
    not g103(n165 ,n236);
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n203), .Q(n4[2]));
    nand g105(n119 ,n3[1] ,n101);
    nand g106(n64 ,n4[30] ,n63);
    not g107(n31 ,n30);
    nor g108(n197 ,n145 ,n178);
    nor g109(n116 ,n101 ,n3[1]);
    nor g110(n190 ,n166 ,n178);
    nor g111(n194 ,n169 ,n178);
    not g112(n100 ,n4[3]);
    xnor g113(n233 ,n4[2] ,n7);
    nand g114(n126 ,n113 ,n120);
    xnor g115(n266 ,n68 ,n3[3]);
    or g116(n139 ,n122 ,n137);
    nor g117(n107 ,n4[8] ,n4[7]);
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n201), .Q(n4[5]));
    or g119(n99 ,n3[2] ,n3[1]);
    xnor g120(n245 ,n32 ,n4[14]);
    not g121(n170 ,n232);
    nor g122(n105 ,n4[30] ,n4[29]);
    xor g123(n232 ,n4[1] ,n4[0]);
    not g124(n29 ,n28);
    nor g125(n184 ,n154 ,n178);
    nor g126(n192 ,n152 ,n178);
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n200), .Q(n4[6]));
    dff g128(.RN(n270), .SN(1'b1), .CK(n0), .D(n4[4]), .Q(n5[4]));
    not g129(n148 ,n249);
    not g130(n11 ,n10);
    buf g131(n259 ,n98);
    nor g132(n72 ,n4[18] ,n4[17]);
    xnor g133(n240 ,n22 ,n4[9]);
    dff g134(.RN(n270), .SN(1'b1), .CK(n0), .D(n4[6]), .Q(n5[6]));
    xnor g135(n253 ,n46 ,n4[22]);
    nor g136(n111 ,n4[28] ,n4[27]);
    nand g137(n7 ,n4[1] ,n4[0]);
    nand g138(n219 ,n3[1] ,n179);
    nor g139(n113 ,n4[14] ,n4[13]);
    nor g140(n128 ,n123 ,n126);
    xnor g141(n257 ,n62 ,n4[30]);
    nor g142(n191 ,n143 ,n178);
    nand g143(n112 ,n3[2] ,n102);
    xnor g144(n237 ,n4[6] ,n16);
    not g145(n159 ,n233);
    not g146(n51 ,n50);
    not g147(n151 ,n255);
    not g148(n19 ,n18);
    nor g149(n264 ,n67 ,n65);
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n199), .Q(n4[8]));
    not g151(n161 ,n263);
    dff g152(.RN(n270), .SN(1'b1), .CK(n0), .D(n4[7]), .Q(n5[7]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n194), .Q(n4[12]));
    nor g154(n77 ,n4[8] ,n4[7]);
    not g155(n164 ,n237);
    nand g156(n36 ,n4[15] ,n35);
    not g157(n182 ,n181);
    xnor g158(n238 ,n4[7] ,n18);
    xnor g159(n250 ,n40 ,n4[19]);
    xnor g160(n262 ,n58 ,n4[28]);
    nand g161(n136 ,n114 ,n134);
    nor g162(n203 ,n159 ,n178);
    nand g163(n50 ,n4[23] ,n49);
    nor g164(n220 ,n150 ,n178);
    nor g165(n210 ,n161 ,n178);
    not g166(n155 ,n239);
    or g167(n227 ,n3[0] ,n221);
    nor g168(n214 ,n153 ,n178);
    nor g169(n202 ,n162 ,n178);
    nor g170(n189 ,n173 ,n178);
    nor g171(n130 ,n3[0] ,n127);
    xnor g172(n256 ,n52 ,n4[25]);
    nor g173(n38 ,n9 ,n36);
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n231), .Q(n3[1]));
    not g175(n156 ,n260);
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n197), .Q(n4[7]));
    nand g177(n52 ,n4[24] ,n51);
    nor g178(n280 ,n277 ,n276);
    not g179(n8 ,n7);
    not g180(n145 ,n238);
    xnor g181(n258 ,n64 ,n4[31]);
    nor g182(n81 ,n4[12] ,n4[11]);
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n195), .Q(n4[11]));
    nor g184(n98 ,n93 ,n97);
    nand g185(n28 ,n4[11] ,n27);
    not g186(n53 ,n52);
    nand g187(n46 ,n4[21] ,n45);
    nand g188(n207 ,n2 ,n178);
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n192), .Q(n4[14]));
    not g190(n169 ,n243);
    nand g191(n267 ,n3[3] ,n99);
    xnor g192(n252 ,n44 ,n4[21]);
    xnor g193(n239 ,n20 ,n4[8]);
    not g194(n150 ,n262);
    nor g195(n75 ,n4[14] ,n4[13]);
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n228), .Q(n3[0]));
    nand g197(n10 ,n4[2] ,n8);
    nor g198(n186 ,n149 ,n178);
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n183), .Q(n4[0]));
    nor g200(n83 ,n4[6] ,n4[5]);
    nor g201(n103 ,n4[22] ,n4[21]);
    nor g202(n140 ,n133 ,n139);
    nand g203(n125 ,n103 ,n110);
    or g204(n97 ,n96 ,n95);
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n184), .Q(n4[22]));
    nor g206(n115 ,n100 ,n3[3]);
    nor g207(n273 ,n4[7] ,n4[1]);
    nor g208(n70 ,n4[24] ,n4[23]);
    nand g209(n121 ,n118 ,n112);
    nor g210(n199 ,n155 ,n178);
    not g211(n69 ,n4[3]);
    xor g212(n249 ,n4[18] ,n38);
    nand g213(n44 ,n4[20] ,n43);
    nor g214(n82 ,n4[30] ,n4[29]);
    nand g215(n89 ,n82 ,n80);
    nand g216(n284 ,n279 ,n280);
    not g217(n166 ,n247);
    nand g218(n34 ,n4[14] ,n33);
    nor g219(n90 ,n69 ,n76);
    xnor g220(n248 ,n39 ,n4[17]);
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n229), .Q(n3[3]));
    nand g222(n26 ,n4[10] ,n25);
    nor g223(n195 ,n167 ,n178);
    nand g224(n276 ,n4[2] ,n4[0]);
    nor g225(n196 ,n172 ,n178);
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n213), .Q(n4[26]));
    not g227(n147 ,n252);
    nand g228(n62 ,n4[29] ,n61);
    nor g229(n180 ,n174 ,n176);
    nand g230(n281 ,n272 ,n271);
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n187), .Q(n4[19]));
    nor g232(n74 ,n4[22] ,n4[21]);
    not g233(n15 ,n14);
    not g234(n167 ,n242);
    not g235(n270 ,n1);
    nor g236(n92 ,n89 ,n87);
    not g237(n173 ,n248);
    nand g238(n124 ,n108 ,n107);
    nand g239(n230 ,n218 ,n224);
    dff g240(.RN(n270), .SN(1'b1), .CK(n0), .D(n4[3]), .Q(n5[3]));
    not g241(n61 ,n60);
    nand g242(n211 ,n3[0] ,n179);
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n209), .Q(n4[30]));
    nor g244(n216 ,n151 ,n178);
    nor g245(n65 ,n3[1] ,n3[0]);
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n230), .Q(n3[2]));
    nand g247(n84 ,n72 ,n71);
    nor g248(n209 ,n144 ,n178);
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n204), .Q(n4[1]));
    not g250(n59 ,n58);
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n216), .Q(n4[24]));
    nand g252(n275 ,n5[1] ,n5[3]);
    nand g253(n54 ,n4[25] ,n53);
    not g254(n144 ,n257);
    nor g255(n114 ,n4[26] ,n4[23]);
    nand g256(n96 ,n83 ,n94);
    or g257(n283 ,n281 ,n282);
    dff g258(.RN(n270), .SN(1'b1), .CK(n0), .D(n285), .Q(n6));
    nor g259(n106 ,n4[18] ,n4[17]);
    nand g260(n282 ,n278 ,n273);
    xnor g261(n255 ,n50 ,n4[24]);
    nand g262(n225 ,n264 ,n222);
    nor g263(n272 ,n5[0] ,n5[2]);
    nor g264(n71 ,n4[16] ,n4[15]);
    xnor g265(n254 ,n48 ,n4[23]);
    nor g266(n212 ,n163 ,n178);
    not g267(n13 ,n12);
    nor g268(n204 ,n170 ,n178);
    or g269(n93 ,n88 ,n86);
    not g270(n176 ,n175);
    xnor g271(n242 ,n26 ,n4[11]);
    not g272(n143 ,n246);
    not g273(n49 ,n48);
    nor g274(n73 ,n4[10] ,n4[9]);
    nand g275(n87 ,n78 ,n70);
    nand g276(n229 ,n217 ,n223);
    nor g277(n79 ,n4[20] ,n4[19]);
    xnor g278(n235 ,n4[4] ,n12);
    nor g279(n76 ,n4[2] ,n4[1]);
    nor g280(n175 ,n1 ,n6);
    nor g281(n108 ,n4[10] ,n4[9]);
    xnor g282(n251 ,n42 ,n4[20]);
    nand g283(n217 ,n3[3] ,n179);
    not g284(n101 ,n4[1]);
    not g285(n55 ,n54);
    nand g286(n95 ,n92 ,n91);
    nand g287(n118 ,n3[3] ,n100);
    dff g288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n210), .Q(n4[29]));
    nand g289(n88 ,n75 ,n81);
    nand g290(n85 ,n74 ,n79);
    not g291(n102 ,n4[2]);
    dff g292(.RN(n270), .SN(1'b1), .CK(n0), .D(n4[1]), .Q(n5[1]));
    not g293(n37 ,n36);
    not g294(n162 ,n235);
    xnor g295(n265 ,n3[2] ,n66);
    not g296(n35 ,n34);
    nor g297(n193 ,n157 ,n178);
    nand g298(n274 ,n5[5] ,n5[7]);
    xnor g299(n263 ,n60 ,n4[29]);
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n190), .Q(n4[16]));
    nand g301(n228 ,n211 ,n227);
    or g302(n131 ,n4[24] ,n125);
    nand g303(n86 ,n73 ,n77);
    not g304(n17 ,n16);
    dff g305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n196), .Q(n4[10]));
    nor g306(n201 ,n165 ,n178);
    nor g307(n185 ,n147 ,n178);
    nor g308(n183 ,n4[0] ,n178);
    not g309(n23 ,n22);
    nor g310(n279 ,n275 ,n274);
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n188), .Q(n4[18]));
    not g312(n27 ,n26);
    dff g313(.RN(n270), .SN(1'b1), .CK(n0), .D(n4[2]), .Q(n5[2]));
    not g314(n21 ,n20);
    nand g315(n277 ,n4[6] ,n4[4]);
    nor g316(n134 ,n4[25] ,n131);
    not g317(n163 ,n261);
    dff g318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n215), .Q(n4[25]));
    nor g319(n80 ,n4[28] ,n4[27]);
    nor g320(n138 ,n121 ,n135);
    nor g321(n94 ,n4[4] ,n90);
    not g322(n158 ,n234);
    xnor g323(n236 ,n4[5] ,n14);
    nand g324(n127 ,n4[0] ,n119);
endmodule
