module top (n0, n1, n3, n5, n6, n7, n4, n2, n8, n9, n10, n11, n12, n14, n13);
    input n0, n1, n2;
    input [1:0] n3, n4;
    input [15:0] n5;
    input [31:0] n6;
    input [3:0] n7;
    output [31:0] n8;
    output n9, n10;
    output [3:0] n11;
    output [7:0] n12, n13;
    output [15:0] n14;
    wire n0, n1, n2;
    wire [1:0] n3, n4;
    wire [15:0] n5;
    wire [31:0] n6;
    wire [3:0] n7;
    wire [31:0] n8;
    wire n9, n10;
    wire [3:0] n11;
    wire [7:0] n12, n13;
    wire [15:0] n14;
    wire [3:0] n15;
    wire [1:0] n16;
    wire [15:0] n17;
    wire [3:0] n18;
    wire [2:0] n19;
    wire [31:0] n20;
    wire n21, n22, n23, n24, n25, n26, n27, n28;
    wire n29, n30, n31, n32, n33, n34, n35, n36;
    wire n37, n38, n39, n40, n41, n42, n43, n44;
    wire n45, n46, n47, n48, n49, n50, n51, n52;
    wire n53, n54, n55, n56, n57, n58, n59, n60;
    wire n61, n62, n63, n64, n65, n66, n67, n68;
    wire n69, n70, n71, n72, n73, n74, n75, n76;
    wire n77, n78, n79, n80, n81, n82, n83, n84;
    wire n85, n86, n87, n88, n89, n90, n91, n92;
    wire n93, n94, n95, n96, n97, n98, n99, n100;
    wire n101, n102, n103, n104, n105, n106, n107, n108;
    wire n109, n110, n111, n112, n113, n114, n115, n116;
    wire n117, n118, n119, n120, n121, n122, n123, n124;
    wire n125, n126, n127, n128, n129, n130, n131, n132;
    wire n133, n134, n135, n136, n137, n138, n139, n140;
    wire n141, n142, n143, n144, n145, n146, n147, n148;
    wire n149, n150, n151, n152, n153, n154, n155, n156;
    wire n157, n158, n159, n160, n161, n162, n163, n164;
    wire n165, n166, n167, n168, n169, n170, n171, n172;
    wire n173, n174, n175, n176, n177, n178, n179, n180;
    wire n181, n182, n183, n184, n185, n186, n187, n188;
    wire n189, n190, n191, n192, n193, n194, n195, n196;
    wire n197, n198, n199, n200, n201, n202, n203, n204;
    wire n205, n206, n207, n208, n209, n210, n211, n212;
    wire n213, n214, n215, n216, n217, n218, n219, n220;
    wire n221, n222, n223, n224, n225, n226, n227, n228;
    wire n229, n230, n231, n232, n233, n234, n235, n236;
    wire n237, n238, n239, n240, n241, n242, n243, n244;
    wire n245, n246, n247, n248, n249, n250, n251, n252;
    wire n253, n254, n255, n256, n257, n258, n259, n260;
    wire n261, n262, n263, n264, n265, n266, n267, n268;
    wire n269, n270, n271, n272, n273, n274, n275, n276;
    wire n277, n278, n279, n280, n281, n282, n283, n284;
    wire n285, n286, n287, n288, n289, n290, n291, n292;
    wire n293, n294, n295, n296, n297, n298, n299, n300;
    wire n301, n302, n303, n304, n305, n306, n307, n308;
    wire n309, n310, n311, n312, n313, n314, n315, n316;
    wire n317, n318, n319, n320, n321, n322, n323, n324;
    wire n325, n326, n327, n328, n329, n330, n331, n332;
    wire n333, n334, n335, n336, n337, n338, n339, n340;
    wire n341, n342, n343, n344, n345, n346, n347, n348;
    wire n349, n350, n351, n352, n353, n354, n355, n356;
    wire n357, n358, n359, n360, n361, n362, n363, n364;
    wire n365, n366, n367, n368, n369, n370, n371, n372;
    wire n373, n374, n375, n376, n377, n378, n379, n380;
    wire n381, n382, n383, n384, n385, n386, n387, n388;
    wire n389, n390, n391, n392, n393, n394, n395, n396;
    wire n397, n398, n399, n400, n401;
    nand g0(n278 ,n8[14] ,n201);
    nand g1(n63 ,n14[10] ,n62);
    nand g2(n116 ,n19[1] ,n88);
    nor g3(n388 ,n67 ,n69);
    dff g4(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n363), .Q(n11[0]));
    nand g5(n277 ,n8[15] ,n201);
    dff g6(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n298), .Q(n16[1]));
    nand g7(n322 ,n165 ,n218);
    dff g8(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n133), .Q(n20[5]));
    nand g9(n68 ,n14[13] ,n66);
    nand g10(n54 ,n14[5] ,n52);
    xnor g11(n386 ,n14[15] ,n70);
    dff g12(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n308), .Q(n14[8]));
    nand g13(n109 ,n379 ,n83);
    nand g14(n237 ,n399 ,n153);
    not g15(n111 ,n110);
    nand g16(n305 ,n190 ,n228);
    nor g17(n103 ,n20[0] ,n82);
    dff g18(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n120), .Q(n20[9]));
    buf g19(n8[21], 1'b0);
    nor g20(n59 ,n44 ,n58);
    nand g21(n313 ,n199 ,n236);
    dff g22(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n372), .Q(n19[1]));
    nand g23(n146 ,n5[6] ,n111);
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n313), .Q(n14[3]));
    dff g25(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n294), .Q(n17[0]));
    nor g26(n283 ,n18[1] ,n206);
    nand g27(n211 ,n11[2] ,n155);
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n353), .Q(n8[2]));
    nor g29(n92 ,n72 ,n71);
    not g30(n64 ,n63);
    xnor g31(n377 ,n20[2] ,n30);
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n315), .Q(n14[1]));
    nand g33(n106 ,n373 ,n102);
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n128), .Q(n20[2]));
    nor g35(n139 ,n75 ,n115);
    buf g36(n8[30], 1'b0);
    nand g37(n294 ,n148 ,n183);
    nand g38(n208 ,n14[1] ,n154);
    nand g39(n254 ,n17[4] ,n200);
    nand g40(n210 ,n11[3] ,n155);
    nand g41(n221 ,n17[12] ,n151);
    not g42(n129 ,n123);
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n340), .Q(n8[15]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n129), .Q(n20[7]));
    nor g45(n284 ,n204 ,n202);
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n349), .Q(n8[6]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n323), .Q(n17[14]));
    nand g48(n357 ,n19[1] ,n328);
    buf g49(n8[29], 1'b0);
    buf g50(n8[22], 1'b0);
    not g51(n128 ,n122);
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n345), .Q(n8[10]));
    buf g53(n13[0], 1'b0);
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n320), .Q(n18[1]));
    nor g55(n174 ,n104 ,n158);
    nor g56(n358 ,n375 ,n285);
    nand g57(n225 ,n387 ,n153);
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n93), .Q(n13[4]));
    nand g59(n245 ,n17[14] ,n200);
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n269), .Q(n17[8]));
    nand g61(n259 ,n18[3] ,n200);
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n325), .Q(n17[12]));
    nand g63(n27 ,n20[7] ,n26);
    nand g64(n272 ,n8[19] ,n201);
    nand g65(n61 ,n14[9] ,n59);
    nand g66(n352 ,n295 ,n259);
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n312), .Q(n14[4]));
    nand g68(n263 ,n17[5] ,n200);
    nor g69(n154 ,n71 ,n117);
    buf g70(n8[27], 1'b0);
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n92), .Q(n13[5]));
    nand g72(n164 ,n7[0] ,n111);
    nand g73(n183 ,n17[0] ,n151);
    nand g74(n307 ,n192 ,n230);
    buf g75(n12[2], 1'b0);
    nand g76(n273 ,n8[18] ,n201);
    nor g77(n93 ,n76 ,n71);
    xnor g78(n399 ,n14[2] ,n47);
    nand g79(n217 ,n18[0] ,n151);
    nand g80(n316 ,n8[9] ,n201);
    nand g81(n37 ,n20[5] ,n36);
    not g82(n329 ,n328);
    xnor g83(n374 ,n15[1] ,n15[0]);
    xnor g84(n384 ,n20[9] ,n42);
    nor g85(n104 ,n10 ,n86);
    or g86(n204 ,n71 ,n137);
    nand g87(n171 ,n73 ,n153);
    nand g88(n318 ,n161 ,n214);
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n85), .Q(n13[6]));
    nand g90(n222 ,n17[11] ,n151);
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n351), .Q(n8[4]));
    not g92(n121 ,n109);
    nand g93(n332 ,n90 ,n283);
    nand g94(n186 ,n14[14] ,n154);
    nand g95(n163 ,n7[1] ,n111);
    nand g96(n240 ,n385 ,n134);
    not g97(n45 ,n14[12]);
    or g98(n135 ,n98 ,n114);
    nand g99(n195 ,n14[6] ,n154);
    nor g100(n39 ,n20[7] ,n38);
    nand g101(n95 ,n11[1] ,n1);
    nand g102(n168 ,n5[11] ,n111);
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n270), .Q(n17[7]));
    nand g104(n261 ,n18[1] ,n200);
    nand g105(n166 ,n5[14] ,n111);
    buf g106(n12[1], 1'b0);
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n336), .Q(n8[19]));
    nand g108(n51 ,n14[3] ,n50);
    nand g109(n292 ,n8[5] ,n201);
    nand g110(n47 ,n14[1] ,n14[0]);
    nand g111(n269 ,n144 ,n178);
    not g112(n73 ,n14[0]);
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n268), .Q(n17[9]));
    nand g114(n342 ,n279 ,n266);
    nand g115(n142 ,n5[10] ,n111);
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n318), .Q(n18[3]));
    nand g117(n325 ,n170 ,n221);
    nand g118(n98 ,n11[0] ,n1);
    nand g119(n194 ,n14[7] ,n154);
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n324), .Q(n17[13]));
    not g121(n133 ,n127);
    nand g122(n362 ,n210 ,n360);
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n244), .Q(n14[0]));
    nand g124(n223 ,n14[2] ,n154);
    nand g125(n265 ,n110 ,n240);
    not g126(n41 ,n40);
    nand g127(n35 ,n20[4] ,n34);
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n304), .Q(n14[12]));
    nand g129(n165 ,n5[15] ,n111);
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n346), .Q(n8[9]));
    nor g131(n134 ,n2 ,n112);
    not g132(n62 ,n61);
    not g133(n207 ,n206);
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n352), .Q(n8[3]));
    nand g135(n282 ,n8[11] ,n201);
    xnor g136(n381 ,n20[6] ,n37);
    nand g137(n192 ,n14[9] ,n154);
    or g138(n79 ,n15[0] ,n15[2]);
    nand g139(n303 ,n150 ,n188);
    nand g140(n238 ,n400 ,n153);
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n314), .Q(n14[2]));
    nand g142(n370 ,n211 ,n331);
    nor g143(n392 ,n60 ,n62);
    nand g144(n178 ,n17[8] ,n151);
    nand g145(n209 ,n14[0] ,n154);
    nand g146(n291 ,n8[8] ,n201);
    nand g147(n24 ,n20[6] ,n20[5]);
    nand g148(n295 ,n8[3] ,n201);
    nand g149(n334 ,n15[1] ,n242);
    xnor g150(n390 ,n14[11] ,n63);
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n342), .Q(n8[13]));
    nor g152(n94 ,n76 ,n16[1]);
    nand g153(n321 ,n164 ,n217);
    not g154(n82 ,n83);
    nand g155(n112 ,n89 ,n88);
    nand g156(n231 ,n393 ,n153);
    nand g157(n250 ,n17[8] ,n200);
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n321), .Q(n18[0]));
    nand g159(n327 ,n8[10] ,n201);
    not g160(n36 ,n35);
    nand g161(n70 ,n14[14] ,n69);
    not g162(n48 ,n47);
    nand g163(n141 ,n2 ,n113);
    nand g164(n220 ,n17[13] ,n151);
    xnor g165(n393 ,n14[8] ,n58);
    not g166(n75 ,n19[2]);
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n96), .Q(n13[3]));
    or g168(n360 ,n100 ,n330);
    nand g169(n233 ,n395 ,n153);
    xnor g170(n398 ,n14[3] ,n49);
    nand g171(n336 ,n272 ,n257);
    nand g172(n180 ,n17[6] ,n151);
    nand g173(n333 ,n141 ,n286);
    nand g174(n315 ,n208 ,n238);
    nand g175(n248 ,n17[10] ,n200);
    nand g176(n348 ,n289 ,n253);
    nand g177(n236 ,n398 ,n153);
    not g178(n85 ,n84);
    nand g179(n320 ,n163 ,n216);
    nand g180(n196 ,n14[5] ,n154);
    nand g181(n247 ,n17[11] ,n200);
    nand g182(n123 ,n382 ,n83);
    xnor g183(n389 ,n14[12] ,n65);
    nand g184(n355 ,n299 ,n262);
    nand g185(n145 ,n5[7] ,n111);
    nand g186(n317 ,n159 ,n198);
    nand g187(n125 ,n381 ,n83);
    nand g188(n301 ,n186 ,n225);
    not g189(n157 ,n156);
    nand g190(n158 ,n1 ,n112);
    nand g191(n300 ,n185 ,n224);
    nand g192(n127 ,n380 ,n83);
    nand g193(n276 ,n8[16] ,n201);
    nand g194(n122 ,n377 ,n83);
    not g195(n131 ,n125);
    nand g196(n270 ,n145 ,n179);
    buf g197(n8[26], 1'b0);
    xor g198(n361 ,n202 ,n15[0]);
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n303), .Q(n16[0]));
    nand g200(n49 ,n14[2] ,n48);
    xnor g201(n395 ,n14[6] ,n54);
    nand g202(n147 ,n5[4] ,n111);
    nand g203(n216 ,n18[1] ,n151);
    nand g204(n323 ,n166 ,n219);
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n130), .Q(n20[8]));
    nor g206(n86 ,n19[1] ,n19[2]);
    nand g207(n124 ,n383 ,n83);
    nor g208(n151 ,n71 ,n111);
    nand g209(n302 ,n187 ,n226);
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n362), .Q(n11[3]));
    nand g211(n274 ,n146 ,n180);
    nand g212(n30 ,n20[1] ,n20[0]);
    not g213(n28 ,n20[2]);
    nand g214(n310 ,n195 ,n233);
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n370), .Q(n11[2]));
    nand g216(n319 ,n162 ,n215);
    nand g217(n364 ,n334 ,n356);
    nor g218(n21 ,n15[1] ,n15[0]);
    nand g219(n255 ,n17[2] ,n200);
    nand g220(n234 ,n396 ,n153);
    nand g221(n256 ,n17[1] ,n200);
    nand g222(n150 ,n3[0] ,n111);
    nand g223(n206 ,n78 ,n153);
    nand g224(n252 ,n17[6] ,n200);
    nor g225(n23 ,n20[4] ,n20[3]);
    buf g226(n8[28], 1'b0);
    nor g227(n173 ,n115 ,n157);
    nand g228(n299 ,n8[0] ,n201);
    nand g229(n214 ,n18[3] ,n151);
    xnor g230(n383 ,n20[8] ,n40);
    nand g231(n239 ,n17[10] ,n151);
    buf g232(n8[23], 1'b0);
    nand g233(n314 ,n223 ,n237);
    nand g234(n337 ,n273 ,n245);
    nand g235(n312 ,n197 ,n235);
    nor g236(n90 ,n18[0] ,n18[3]);
    nor g237(n115 ,n15[1] ,n79);
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n348), .Q(n8[7]));
    or g239(n401 ,n15[0] ,n22);
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n311), .Q(n14[5]));
    nand g241(n235 ,n397 ,n153);
    nand g242(n202 ,n106 ,n138);
    nand g243(n345 ,n327 ,n252);
    nand g244(n363 ,n135 ,n332);
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n341), .Q(n8[14]));
    buf g246(n137 ,n115);
    nor g247(n32 ,n20[3] ,n31);
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n319), .Q(n18[2]));
    nand g249(n330 ,n18[1] ,n207);
    not g250(n96 ,n95);
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n354), .Q(n8[1]));
    nand g252(n287 ,n169 ,n189);
    nand g253(n266 ,n17[9] ,n200);
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n343), .Q(n8[12]));
    nand g255(n341 ,n278 ,n248);
    nor g256(n396 ,n53 ,n55);
    nand g257(n184 ,n16[1] ,n151);
    nand g258(n229 ,n391 ,n153);
    or g259(n172 ,n105 ,n158);
    nand g260(n226 ,n388 ,n153);
    nand g261(n365 ,n136 ,n359);
    not g262(n130 ,n124);
    not g263(n44 ,n14[8]);
    nand g264(n143 ,n5[1] ,n111);
    dff g265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n347), .Q(n8[8]));
    nand g266(n350 ,n292 ,n256);
    buf g267(n12[3], 1'b0);
    nor g268(n385 ,n24 ,n27);
    not g269(n117 ,n116);
    nand g270(n213 ,n14[12] ,n154);
    dff g271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n300), .Q(n14[15]));
    or g272(n372 ,n265 ,n366);
    buf g273(n13[1], 1'b0);
    nand g274(n280 ,n160 ,n212);
    nand g275(n193 ,n14[8] ,n154);
    nor g276(n83 ,n71 ,n385);
    nand g277(n177 ,n17[9] ,n151);
    xnor g278(n397 ,n14[4] ,n51);
    nor g279(n156 ,n84 ,n118);
    nand g280(n246 ,n17[12] ,n200);
    dff g281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n350), .Q(n8[5]));
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n307), .Q(n14[9]));
    nand g283(n102 ,n19[0] ,n19[2]);
    nand g284(n354 ,n297 ,n261);
    nand g285(n251 ,n17[7] ,n200);
    nand g286(n296 ,n8[2] ,n201);
    not g287(n77 ,n18[3]);
    nand g288(n253 ,n17[3] ,n200);
    nand g289(n343 ,n281 ,n250);
    dff g290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n306), .Q(n14[10]));
    nand g291(n289 ,n8[7] ,n201);
    not g292(n120 ,n108);
    nor g293(n38 ,n29 ,n37);
    dff g294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n371), .Q(n15[2]));
    nor g295(n67 ,n14[13] ,n66);
    not g296(n91 ,n90);
    nand g297(n197 ,n14[4] ,n154);
    dff g298(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n364), .Q(n15[1]));
    nand g299(n264 ,n175 ,n240);
    nand g300(n351 ,n293 ,n258);
    nand g301(n190 ,n14[11] ,n154);
    nand g302(n218 ,n17[15] ,n151);
    or g303(n136 ,n95 ,n114);
    dff g304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n333), .Q(n19[0]));
    buf g305(n12[6], 1'b0);
    nand g306(n290 ,n8[6] ,n201);
    nand g307(n25 ,n20[9] ,n20[8]);
    nor g308(n335 ,n329 ,n264);
    nor g309(n89 ,n71 ,n19[1]);
    nand g310(n144 ,n5[8] ,n111);
    not g311(n43 ,n14[4]);
    dff g312(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n326), .Q(n17[11]));
    nand g313(n65 ,n14[11] ,n64);
    nor g314(n382 ,n39 ,n41);
    dff g315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n305), .Q(n14[11]));
    xnor g316(n394 ,n14[7] ,n56);
    nand g317(n268 ,n140 ,n177);
    not g318(n285 ,n284);
    nand g319(n199 ,n14[3] ,n154);
    nand g320(n308 ,n193 ,n231);
    not g321(n78 ,n18[2]);
    buf g322(n8[31], 1'b0);
    nor g323(n31 ,n28 ,n30);
    nor g324(n60 ,n14[9] ,n59);
    nand g325(n324 ,n167 ,n220);
    nand g326(n257 ,n17[15] ,n200);
    nand g327(n306 ,n191 ,n229);
    xnor g328(n391 ,n14[10] ,n61);
    nand g329(n297 ,n8[1] ,n201);
    not g330(n373 ,n401);
    nand g331(n100 ,n18[0] ,n77);
    dff g332(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n280), .Q(n17[5]));
    dff g333(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n288), .Q(n17[1]));
    nor g334(n138 ,n88 ,n118);
    nand g335(n219 ,n17[14] ,n151);
    nand g336(n227 ,n389 ,n153);
    dff g337(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n121), .Q(n20[4]));
    nand g338(n347 ,n291 ,n254);
    not g339(n200 ,n201);
    nand g340(n175 ,n89 ,n139);
    nand g341(n267 ,n142 ,n239);
    nand g342(n340 ,n277 ,n247);
    nand g343(n179 ,n17[7] ,n151);
    xor g344(n375 ,n15[2] ,n21);
    nand g345(n84 ,n19[0] ,n1);
    nand g346(n140 ,n5[9] ,n111);
    nor g347(n242 ,n71 ,n203);
    buf g348(n12[4], 1'b0);
    nand g349(n311 ,n196 ,n234);
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n274), .Q(n17[6]));
    or g351(n331 ,n91 ,n330);
    xnor g352(n379 ,n20[4] ,n33);
    nand g353(n170 ,n5[12] ,n111);
    not g354(n99 ,n98);
    dff g355(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n369), .Q(n19[2]));
    nand g356(n288 ,n143 ,n182);
    nand g357(n304 ,n213 ,n227);
    or g358(n368 ,n241 ,n358);
    nand g359(n97 ,n19[1] ,n19[2]);
    nand g360(n126 ,n376 ,n83);
    dff g361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n367), .Q(n15[0]));
    not g362(n87 ,n86);
    nor g363(n46 ,n14[1] ,n14[0]);
    nor g364(n114 ,n19[0] ,n97);
    nand g365(n118 ,n97 ,n87);
    nand g366(n359 ,n101 ,n283);
    buf g367(n12[0], 1'b0);
    nand g368(n249 ,n17[13] ,n200);
    nor g369(n366 ,n357 ,n286);
    nand g370(n176 ,n94 ,n153);
    nand g371(n148 ,n5[0] ,n111);
    dff g372(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n267), .Q(n17[10]));
    nand g373(n33 ,n20[3] ,n31);
    nand g374(n182 ,n17[1] ,n151);
    nand g375(n258 ,n17[0] ,n200);
    nand g376(n160 ,n5[5] ,n111);
    nor g377(n367 ,n204 ,n361);
    nor g378(n153 ,n71 ,n116);
    nand g379(n230 ,n392 ,n153);
    nand g380(n275 ,n8[17] ,n201);
    dff g381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n338), .Q(n8[17]));
    not g382(n76 ,n16[0]);
    buf g383(n8[25], 1'b0);
    dff g384(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n301), .Q(n14[14]));
    not g385(n132 ,n126);
    dff g386(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n103), .Q(n20[0]));
    buf g387(n8[20], 1'b0);
    nand g388(n293 ,n8[4] ,n201);
    nor g389(n378 ,n32 ,n34);
    nand g390(n232 ,n394 ,n153);
    not g391(n34 ,n33);
    dff g392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n344), .Q(n8[11]));
    buf g393(n12[7], 1'b0);
    dff g394(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n271), .Q(n17[4]));
    nand g395(n107 ,n378 ,n83);
    buf g396(n12[5], 1'b0);
    nor g397(n52 ,n43 ,n51);
    not g398(n119 ,n107);
    nor g399(n155 ,n71 ,n114);
    xor g400(n376 ,n20[1] ,n20[0]);
    or g401(n22 ,n15[2] ,n15[1]);
    nor g402(n371 ,n71 ,n368);
    not g403(n203 ,n202);
    nor g404(n88 ,n19[0] ,n19[2]);
    not g405(n55 ,n54);
    nand g406(n356 ,n374 ,n284);
    dff g407(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n309), .Q(n14[7]));
    nand g408(n328 ,n16[1] ,n205);
    nand g409(n326 ,n168 ,n222);
    dff g410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n310), .Q(n14[6]));
    not g411(n72 ,n16[1]);
    nand g412(n262 ,n18[0] ,n200);
    not g413(n71 ,n1);
    nor g414(n26 ,n25 ,n23);
    dff g415(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n317), .Q(n17[3]));
    xnor g416(n380 ,n20[5] ,n35);
    dff g417(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n80), .Q(n13[7]));
    not g418(n69 ,n68);
    not g419(n57 ,n56);
    dff g420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n337), .Q(n8[18]));
    not g421(n29 ,n20[6]);
    nand g422(n344 ,n282 ,n251);
    not g423(n152 ,n153);
    nand g424(n201 ,n19[1] ,n156);
    nand g425(n353 ,n296 ,n260);
    nand g426(n161 ,n7[3] ,n111);
    nand g427(n188 ,n16[0] ,n151);
    nand g428(n191 ,n14[10] ,n154);
    dff g429(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n322), .Q(n17[15]));
    xnor g430(n387 ,n14[14] ,n68);
    not g431(n50 ,n49);
    nand g432(n279 ,n8[13] ,n201);
    nand g433(n159 ,n5[3] ,n111);
    nor g434(n205 ,n16[0] ,n152);
    dff g435(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n339), .Q(n8[16]));
    nor g436(n286 ,n205 ,n173);
    dff g437(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n243), .Q(n9));
    nor g438(n105 ,n9 ,n81);
    nor g439(n81 ,n19[0] ,n19[1]);
    nand g440(n40 ,n20[7] ,n38);
    dff g441(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n119), .Q(n20[3]));
    nand g442(n58 ,n14[7] ,n57);
    nand g443(n185 ,n14[15] ,n154);
    nand g444(n349 ,n290 ,n255);
    dff g445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n302), .Q(n14[13]));
    nand g446(n298 ,n149 ,n184);
    nand g447(n243 ,n201 ,n172);
    nor g448(n66 ,n45 ,n65);
    dff g449(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n131), .Q(n20[6]));
    nand g450(n339 ,n276 ,n246);
    nand g451(n42 ,n20[8] ,n41);
    nand g452(n212 ,n17[5] ,n151);
    nand g453(n189 ,n17[2] ,n151);
    nand g454(n338 ,n275 ,n249);
    nand g455(n56 ,n14[6] ,n55);
    nand g456(n369 ,n176 ,n335);
    nand g457(n187 ,n14[13] ,n154);
    not g458(n113 ,n112);
    nand g459(n167 ,n5[13] ,n111);
    nand g460(n108 ,n384 ,n83);
    dff g461(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n365), .Q(n11[1]));
    not g462(n101 ,n100);
    dff g463(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n99), .Q(n13[2]));
    nand g464(n309 ,n194 ,n232);
    nand g465(n181 ,n17[4] ,n151);
    nand g466(n271 ,n147 ,n181);
    dff g467(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n174), .Q(n10));
    dff g468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n287), .Q(n17[2]));
    nor g469(n80 ,n74 ,n71);
    nand g470(n162 ,n7[2] ,n111);
    nand g471(n110 ,n85 ,n86);
    nand g472(n169 ,n5[2] ,n111);
    not g473(n74 ,n19[1]);
    nand g474(n346 ,n316 ,n263);
    dff g475(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n132), .Q(n20[1]));
    nand g476(n149 ,n3[1] ,n111);
    dff g477(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n355), .Q(n8[0]));
    nand g478(n281 ,n8[12] ,n201);
    nand g479(n244 ,n209 ,n171);
    nand g480(n224 ,n386 ,n153);
    nor g481(n241 ,n15[2] ,n203);
    nor g482(n400 ,n48 ,n46);
    nand g483(n260 ,n18[2] ,n200);
    nor g484(n53 ,n14[5] ,n52);
    nand g485(n215 ,n18[2] ,n151);
    nand g486(n198 ,n17[3] ,n151);
    nand g487(n228 ,n390 ,n153);
    buf g488(n8[24], 1'b0);
endmodule
