module top (n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12);
    input n0, n1, n2, n3;
    input [1:0] n4, n5;
    output n6, n7;
    output [6:0] n8, n9;
    output [3:0] n10, n11, n12;
    wire n0, n1, n2, n3;
    wire [1:0] n4, n5;
    wire n6, n7;
    wire [6:0] n8, n9;
    wire [3:0] n10, n11, n12;
    wire [2:0] n13;
    wire [15:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66;
    nand g0(n45 ,n4[0] ,n38);
    not g1(n10[0] ,n46);
    xnor g2(n10[2] ,n61 ,n59);
    not g3(n11[0] ,n20);
    nand g4(n14[5] ,n43 ,n66);
    nand g5(n41 ,n5[1] ,n37);
    nand g6(n62 ,n54 ,n57);
    nand g7(n47 ,n4[1] ,n38);
    buf g8(n12[1], 1'b0);
    dff g9(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n27), .Q(n13[0]));
    nand g10(n64 ,n57 ,n63);
    not g11(n25 ,n24);
    nand g12(n48 ,n32 ,n39);
    nor g13(n23 ,n22 ,n6);
    buf g14(n12[3], 1'b0);
    nand g15(n57 ,n33 ,n53);
    nor g16(n61 ,n56 ,n58);
    buf g17(n8[2], 1'b0);
    nor g18(n16 ,n10[3] ,n10[2]);
    not g19(n11[1] ,n21);
    nand g20(n30 ,n5[1] ,n2);
    buf g21(n8[3], n8[6]);
    nor g22(n27 ,n1 ,n26);
    buf g23(n8[5], n8[6]);
    buf g24(n11[3], 1'b0);
    buf g25(n8[0], n8[6]);
    not g26(n22 ,n13[0]);
    nand g27(n50 ,n41 ,n45);
    buf g28(n9[2], n8[6]);
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n23), .Q(n6));
    nand g30(n63 ,n55 ,n60);
    or g31(n43 ,n32 ,n39);
    nand g32(n52 ,n40 ,n47);
    buf g33(n9[6], 1'b0);
    nand g34(n21 ,n14[5] ,n19);
    or g35(n60 ,n58 ,n59);
    nand g36(n44 ,n5[1] ,n38);
    xnor g37(n10[1] ,n34 ,n51);
    nor g38(n15 ,n10[1] ,n10[0]);
    not g39(n37 ,n36);
    buf g40(n12[0], 1'b0);
    buf g41(n9[0], n8[6]);
    nand g42(n39 ,n4[1] ,n37);
    nand g43(n66 ,n48 ,n65);
    or g44(n54 ,n33 ,n53);
    not g45(n31 ,n30);
    buf g46(n11[2], 1'b0);
    buf g47(n8[4], n8[6]);
    buf g48(n9[1], n8[6]);
    nand g49(n36 ,n3 ,n13[0]);
    nor g50(n18 ,n10[3] ,n10[2]);
    nand g51(n55 ,n31 ,n50);
    not g52(n35 ,n34);
    nand g53(n49 ,n48 ,n43);
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n13[0]), .Q(n8[6]));
    nand g55(n34 ,n5[0] ,n2);
    nand g56(n32 ,n4[1] ,n2);
    not g57(n53 ,n52);
    nor g58(n29 ,n3 ,n13[0]);
    nand g59(n19 ,n18 ,n17);
    nand g60(n46 ,n5[0] ,n38);
    buf g61(n9[5], n8[6]);
    nand g62(n20 ,n14[4] ,n19);
    nor g63(n26 ,n13[0] ,n25);
    buf g64(n9[4], n8[6]);
    buf g65(n7, 1'b0);
    nand g66(n42 ,n5[0] ,n37);
    nand g67(n59 ,n35 ,n51);
    nand g68(n40 ,n4[0] ,n37);
    nand g69(n33 ,n4[0] ,n2);
    nor g70(n38 ,n37 ,n29);
    nand g71(n24 ,n2 ,n28);
    nand g72(n65 ,n54 ,n64);
    nor g73(n17 ,n10[1] ,n10[0]);
    buf g74(n8[1], 1'b0);
    buf g75(n9[3], 1'b0);
    not g76(n56 ,n55);
    nor g77(n58 ,n31 ,n50);
    xnor g78(n10[3] ,n62 ,n63);
    nand g79(n28 ,n16 ,n15);
    xnor g80(n14[4] ,n49 ,n65);
    nand g81(n51 ,n42 ,n44);
    buf g82(n12[2], 1'b0);
endmodule
