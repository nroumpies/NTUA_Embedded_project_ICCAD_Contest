module top (n0, n1, n2, n6, n3, n7, n5, n12, n4, n8, n9, n10, n11, n13, n14, n15, n16);
    input n0, n1, n2, n3, n4;
    input [7:0] n5;
    output n6, n7, n8, n9, n10, n11;
    output [7:0] n12, n13, n14, n15;
    output [15:0] n16;
    wire n0, n1, n2, n3, n4;
    wire [7:0] n5;
    wire n6, n7, n8, n9, n10, n11;
    wire [7:0] n12, n13, n14, n15;
    wire [15:0] n16;
    wire [2:0] n17;
    wire [2:0] n18;
    wire [4:0] n19;
    wire [15:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [7:0] n23;
    wire [7:0] n24;
    wire [7:0] n25;
    wire [7:0] n26;
    wire [7:0] n27;
    wire [7:0] n28;
    wire [7:0] n29;
    wire [7:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [7:0] n36;
    wire [3:0] n37;
    wire [3:0] n38;
    wire [7:0] n39;
    wire [15:0] n40;
    wire [2:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [7:0] n44;
    wire [7:0] n45;
    wire [7:0] n46;
    wire [7:0] n47;
    wire [7:0] n48;
    wire [7:0] n49;
    wire [7:0] n50;
    wire [7:0] n51;
    wire [7:0] n52;
    wire [7:0] n53;
    wire [7:0] n54;
    wire [7:0] n55;
    wire [7:0] n56;
    wire [7:0] n57;
    wire [4:0] n58;
    wire [3:0] n59;
    wire [3:0] n60;
    wire [7:0] n61;
    wire [2:0] n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
    wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
    wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
    wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
    wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
    wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
    wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
    wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
    wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
    wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
    wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
    wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
    wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
    wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
    wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
    wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
    wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
    wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
    wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
    wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
    wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
    wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
    wire n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742;
    wire n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750;
    wire n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758;
    wire n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766;
    wire n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774;
    wire n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782;
    wire n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790;
    wire n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798;
    wire n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806;
    wire n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814;
    wire n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822;
    wire n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
    wire n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838;
    wire n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846;
    wire n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854;
    wire n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
    wire n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870;
    wire n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878;
    wire n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886;
    wire n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894;
    wire n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902;
    wire n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910;
    wire n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918;
    wire n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
    wire n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934;
    wire n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
    wire n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950;
    wire n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958;
    wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
    wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974;
    wire n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982;
    wire n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990;
    wire n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998;
    wire n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
    wire n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014;
    wire n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022;
    wire n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;
    wire n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038;
    wire n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046;
    wire n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054;
    wire n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062;
    wire n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070;
    wire n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078;
    wire n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086;
    wire n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094;
    wire n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102;
    wire n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110;
    wire n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118;
    wire n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126;
    wire n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134;
    wire n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142;
    wire n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150;
    wire n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158;
    wire n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166;
    wire n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174;
    wire n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182;
    wire n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190;
    wire n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198;
    wire n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206;
    wire n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214;
    wire n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222;
    wire n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230;
    wire n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238;
    wire n2239, n2240, n2241, n2242, n2243, n2244;
    nand g0(n1785 ,n26[3] ,n1475);
    nand g1(n869 ,n20[8] ,n585);
    nand g2(n1966 ,n844 ,n1780);
    nand g3(n1878 ,n1544 ,n1565);
    dff g4(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2127), .Q(n12[1]));
    nand g5(n1575 ,n46[5] ,n1374);
    nand g6(n158 ,n41[1] ,n41[0]);
    not g7(n118 ,n117);
    nand g8(n106 ,n20[8] ,n20[7]);
    nand g9(n806 ,n5[3] ,n554);
    nand g10(n1859 ,n34[5] ,n1473);
    nand g11(n150 ,n40[5] ,n149);
    nand g12(n1523 ,n57[6] ,n1362);
    not g13(n700 ,n681);
    nand g14(n1014 ,n651 ,n523);
    nor g15(n1511 ,n193 ,n1390);
    nand g16(n1633 ,n39[7] ,n1472);
    nand g17(n2121 ,n1120 ,n2100);
    nand g18(n2058 ,n1898 ,n1645);
    nand g19(n1124 ,n41[0] ,n890);
    nand g20(n2066 ,n1760 ,n1695);
    nand g21(n1529 ,n2209 ,n1385);
    dff g22(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1205), .Q(n45[6]));
    or g23(n1947 ,n1885 ,n1884);
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1968), .Q(n27[6]));
    nand g25(n664 ,n34[3] ,n426);
    nand g26(n474 ,n61[0] ,n383);
    nor g27(n76 ,n19[3] ,n71);
    nand g28(n1182 ,n1023 ,n731);
    nor g29(n890 ,n193 ,n488);
    not g30(n597 ,n507);
    nand g31(n1705 ,n39[1] ,n1471);
    nand g32(n356 ,n2 ,n303);
    nand g33(n881 ,n20[11] ,n585);
    buf g34(n15[2], 1'b0);
    nand g35(n1261 ,n19[3] ,n886);
    not g36(n1578 ,n1516);
    nand g37(n829 ,n5[4] ,n576);
    nand g38(n1438 ,n42[4] ,n1376);
    nand g39(n1026 ,n53[3] ,n560);
    nor g40(n2149 ,n1937 ,n2147);
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1963), .Q(n20[2]));
    nand g42(n1584 ,n33[4] ,n1486);
    nand g43(n973 ,n43[3] ,n562);
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1972), .Q(n27[3]));
    nand g45(n1517 ,n43[6] ,n1363);
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2007), .Q(n23[0]));
    nand g47(n1325 ,n1240 ,n1239);
    not g48(n1387 ,n1318);
    nand g49(n633 ,n26[7] ,n431);
    not g50(n1474 ,n1475);
    nand g51(n935 ,n47[3] ,n566);
    nand g52(n2020 ,n1734 ,n1663);
    nand g53(n1299 ,n941 ,n746);
    nor g54(n2105 ,n1927 ,n1926);
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1268), .Q(n46[3]));
    nand g56(n153 ,n40[7] ,n151);
    nand g57(n905 ,n52[2] ,n572);
    nor g58(n145 ,n40[3] ,n144);
    nand g59(n1418 ,n55[2] ,n1370);
    xnor g60(n2214 ,n20[8] ,n177);
    nand g61(n1166 ,n845 ,n810);
    nand g62(n910 ,n51[7] ,n570);
    nand g63(n789 ,n5[2] ,n565);
    nand g64(n1634 ,n39[6] ,n1472);
    nor g65(n165 ,n20[1] ,n20[0]);
    nand g66(n669 ,n25[3] ,n476);
    nor g67(n1589 ,n1058 ,n1567);
    nand g68(n132 ,n58[1] ,n58[0]);
    nand g69(n1988 ,n1793 ,n1602);
    nand g70(n945 ,n46[3] ,n568);
    nand g71(n965 ,n688 ,n627);
    nand g72(n1801 ,n24[3] ,n1479);
    nand g73(n1020 ,n656 ,n524);
    nand g74(n1834 ,n1514 ,n1154);
    nand g75(n1156 ,n918 ,n722);
    nand g76(n1515 ,n57[2] ,n1362);
    nor g77(n1335 ,n209 ,n1311);
    nand g78(n1339 ,n62[0] ,n1194);
    nand g79(n325 ,n194 ,n257);
    or g80(n2180 ,n19[4] ,n17[0]);
    nand g81(n880 ,n20[2] ,n585);
    nand g82(n1173 ,n852 ,n816);
    nor g83(n2184 ,n2180 ,n2183);
    nand g84(n326 ,n41[2] ,n281);
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1998), .Q(n24[1]));
    nand g86(n1855 ,n34[6] ,n1473);
    nand g87(n1838 ,n1519 ,n1417);
    nand g88(n924 ,n50[1] ,n574);
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2051), .Q(n33[0]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2053), .Q(n32[6]));
    nor g91(n1326 ,n193 ,n1313);
    nand g92(n1272 ,n1070 ,n785);
    nor g93(n1351 ,n1104 ,n1108);
    nand g94(n1073 ,n56[5] ,n575);
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1582), .Q(n17[1]));
    nand g96(n1301 ,n1060 ,n794);
    nand g97(n852 ,n48[7] ,n563);
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1216), .Q(n44[3]));
    or g99(n1936 ,n1850 ,n1849);
    nand g100(n1290 ,n866 ,n831);
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1146), .Q(n52[2]));
    nand g102(n816 ,n5[7] ,n564);
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2083), .Q(n20[8]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1224), .Q(n43[3]));
    xnor g105(n2195 ,n37[3] ,n162);
    nor g106(n1245 ,n192 ,n1082);
    nand g107(n1653 ,n39[0] ,n1472);
    nor g108(n373 ,n195 ,n327);
    nand g109(n1663 ,n39[7] ,n1467);
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1266), .Q(n53[2]));
    xnor g111(n2211 ,n20[2] ,n166);
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1994), .Q(n24[5]));
    nor g113(n377 ,n218 ,n328);
    nand g114(n505 ,n30[1] ,n425);
    not g115(n231 ,n41[0]);
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n286), .Q(n16[3]));
    nand g117(n1613 ,n39[6] ,n1480);
    nand g118(n1614 ,n39[5] ,n1480);
    xnor g119(n2204 ,n20[10] ,n180);
    nand g120(n1495 ,n266 ,n1384);
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2012), .Q(n22[3]));
    nand g122(n1522 ,n47[4] ,n1371);
    nand g123(n1870 ,n1500 ,n1400);
    nand g124(n996 ,n462 ,n645);
    nand g125(n1919 ,n31[7] ,n1490);
    not g126(n477 ,n478);
    nand g127(n1297 ,n1066 ,n720);
    nand g128(n478 ,n2236 ,n395);
    nand g129(n1986 ,n1792 ,n1600);
    not g130(n1391 ,n1323);
    nand g131(n1221 ,n970 ,n759);
    nand g132(n1566 ,n55[6] ,n1370);
    nand g133(n653 ,n26[0] ,n431);
    nand g134(n2002 ,n1807 ,n1614);
    nand g135(n1155 ,n916 ,n723);
    nand g136(n1746 ,n35[2] ,n1492);
    nand g137(n793 ,n5[2] ,n557);
    nand g138(n665 ,n34[4] ,n426);
    nand g139(n1899 ,n32[0] ,n1489);
    nor g140(n1580 ,n952 ,n1411);
    nand g141(n1796 ,n25[0] ,n1477);
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2074), .Q(n20[9]));
    nor g143(n895 ,n59[3] ,n586);
    nand g144(n1605 ,n39[7] ,n1478);
    nand g145(n1424 ,n46[6] ,n1374);
    nand g146(n1481 ,n272 ,n1384);
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1186), .Q(n47[3]));
    buf g148(n14[4], 1'b0);
    nand g149(n1023 ,n47[7] ,n566);
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2010), .Q(n22[5]));
    not g151(n167 ,n166);
    nor g152(n466 ,n234 ,n379);
    not g153(n1314 ,n1269);
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1151), .Q(n51[5]));
    nand g155(n641 ,n28[0] ,n432);
    nand g156(n1751 ,n33[7] ,n1486);
    nand g157(n342 ,n18[1] ,n293);
    nand g158(n813 ,n5[2] ,n580);
    nand g159(n842 ,n17[1] ,n495);
    nand g160(n639 ,n35[0] ,n435);
    buf g161(n15[3], n13[1]);
    nor g162(n406 ,n2 ,n310);
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1296), .Q(n55[2]));
    nand g164(n1239 ,n2234 ,n889);
    not g165(n583 ,n584);
    nand g166(n649 ,n24[6] ,n428);
    nand g167(n757 ,n5[0] ,n555);
    nand g168(n1441 ,n52[2] ,n1368);
    nand g169(n381 ,n273 ,n326);
    nand g170(n2004 ,n1809 ,n1616);
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2069), .Q(n31[1]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1958), .Q(n20[0]));
    nand g173(n1772 ,n28[7] ,n1468);
    nand g174(n1016 ,n2195 ,n593);
    nor g175(n375 ,n198 ,n327);
    nand g176(n1879 ,n1545 ,n1531);
    nand g177(n1545 ,n47[1] ,n1371);
    nand g178(n767 ,n5[6] ,n583);
    nor g179(n871 ,n212 ,n595);
    nand g180(n874 ,n58[1] ,n589);
    nand g181(n1668 ,n39[2] ,n1467);
    not g182(n139 ,n138);
    nand g183(n1876 ,n1446 ,n1441);
    nand g184(n867 ,n58[0] ,n589);
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1295), .Q(n55[3]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2102), .Q(n21[2]));
    nand g187(n2018 ,n1823 ,n1628);
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n280), .Q(n15[7]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1301), .Q(n54[6]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1925), .Q(n62[0]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2101), .Q(n21[0]));
    nand g192(n779 ,n5[1] ,n567);
    nand g193(n399 ,n2230 ,n330);
    or g194(n248 ,n41[0] ,n41[2]);
    nand g195(n812 ,n5[3] ,n580);
    nor g196(n2153 ,n1949 ,n2143);
    nand g197(n558 ,n264 ,n480);
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1999), .Q(n24[0]));
    nor g199(n472 ,n362 ,n375);
    nand g200(n2038 ,n1859 ,n1635);
    or g201(n320 ,n222 ,n257);
    buf g202(n15[5], n13[5]);
    nand g203(n323 ,n37[1] ,n255);
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n292), .Q(n16[5]));
    nor g205(n1248 ,n193 ,n1084);
    dff g206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1510), .Q(n19[2]));
    nand g207(n1775 ,n28[4] ,n1468);
    or g208(n404 ,n60[0] ,n329);
    nor g209(n362 ,n196 ,n328);
    nor g210(n1507 ,n192 ,n1391);
    nand g211(n720 ,n5[1] ,n581);
    nand g212(n2175 ,n1559 ,n2169);
    not g213(n569 ,n570);
    nor g214(n2152 ,n1940 ,n2144);
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2104), .Q(n21[3]));
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1217), .Q(n44[2]));
    nand g217(n1698 ,n39[1] ,n1491);
    nand g218(n1414 ,n55[7] ,n1370);
    not g219(n1478 ,n1479);
    nand g220(n1642 ,n39[4] ,n1488);
    nand g221(n999 ,n633 ,n631);
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2081), .Q(n20[6]));
    nand g223(n2016 ,n1821 ,n1626);
    nand g224(n1557 ,n57[5] ,n1362);
    nor g225(n1483 ,n298 ,n1383);
    nor g226(n331 ,n192 ,n307);
    nand g227(n917 ,n620 ,n550);
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1974), .Q(n27[1]));
    nor g229(n317 ,n62[2] ,n274);
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1960), .Q(n59[1]));
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n287), .Q(n16[6]));
    nand g232(n1146 ,n905 ,n714);
    nand g233(n1897 ,n1460 ,n1459);
    nand g234(n1489 ,n272 ,n1382);
    nor g235(n2161 ,n1578 ,n2148);
    or g236(n370 ,n199 ,n319);
    nand g237(n1999 ,n1804 ,n1656);
    nand g238(n162 ,n37[2] ,n161);
    not g239(n1496 ,n1497);
    nand g240(n530 ,n30[3] ,n425);
    nor g241(n124 ,n20[7] ,n123);
    or g242(n1105 ,n1027 ,n1029);
    nand g243(n1964 ,n1724 ,n1713);
    nor g244(n108 ,n105 ,n103);
    nand g245(n94 ,n40[1] ,n40[0]);
    nand g246(n613 ,n27[1] ,n424);
    nor g247(n435 ,n258 ,n402);
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1140), .Q(n53[0]));
    nand g249(n173 ,n20[5] ,n171);
    nand g250(n689 ,n24[2] ,n428);
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2087), .Q(n20[7]));
    nand g252(n940 ,n46[7] ,n568);
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2063), .Q(n59[3]));
    not g254(n1470 ,n1471);
    nand g255(n1222 ,n971 ,n760);
    buf g256(n16[12], 1'b0);
    nand g257(n621 ,n2217 ,n421);
    nand g258(n715 ,n5[1] ,n571);
    nor g259(n1252 ,n192 ,n1088);
    nand g260(n1262 ,n19[2] ,n886);
    nand g261(n1957 ,n1110 ,n1589);
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2009), .Q(n22[7]));
    or g263(n1948 ,n1888 ,n1887);
    nand g264(n961 ,n44[7] ,n556);
    not g265(n586 ,n587);
    dff g266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1189), .Q(n47[0]));
    nand g267(n1826 ,n21[2] ,n1495);
    dff g268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1305), .Q(n54[2]));
    nand g269(n922 ,n50[2] ,n574);
    dff g270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1223), .Q(n43[4]));
    nand g271(n1172 ,n863 ,n815);
    not g272(n95 ,n94);
    nand g273(n1594 ,n39[3] ,n1474);
    nand g274(n808 ,n5[0] ,n554);
    nand g275(n1656 ,n39[0] ,n1478);
    nand g276(n1159 ,n1041 ,n725);
    nor g277(n1382 ,n204 ,n1202);
    nand g278(n1593 ,n39[4] ,n1474);
    nand g279(n1678 ,n39[1] ,n1483);
    not g280(n205 ,n60[0]);
    nand g281(n2006 ,n1811 ,n1618);
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1969), .Q(n27[5]));
    not g283(n221 ,n17[2]);
    nand g284(n1473 ,n260 ,n1382);
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2058), .Q(n32[1]));
    nor g286(n488 ,n473 ,n446);
    nand g287(n1230 ,n979 ,n768);
    not g288(n1492 ,n1493);
    nand g289(n2135 ,n1547 ,n2111);
    nand g290(n403 ,n37[2] ,n340);
    nand g291(n1452 ,n44[0] ,n1366);
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1164), .Q(n50[0]));
    nand g293(n726 ,n5[4] ,n573);
    nand g294(n925 ,n608 ,n626);
    or g295(n1098 ,n1011 ,n1010);
    nand g296(n1730 ,n27[2] ,n1482);
    nor g297(n395 ,n4 ,n332);
    nand g298(n690 ,n34[0] ,n426);
    not g299(n147 ,n146);
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1153), .Q(n51[3]));
    nor g301(n1720 ,n193 ,n1397);
    nand g302(n1625 ,n39[1] ,n1496);
    not g303(n226 ,n59[1]);
    nand g304(n1360 ,n333 ,n1195);
    nand g305(n1711 ,n39[3] ,n1469);
    nor g306(n1246 ,n192 ,n1083);
    dff g307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1272), .Q(n53[6]));
    nand g308(n712 ,n5[4] ,n571);
    nand g309(n189 ,n38[2] ,n188);
    nand g310(n1818 ,n22[2] ,n1497);
    nor g311(n2201 ,n172 ,n174);
    nand g312(n1079 ,n59[3] ,n587);
    nand g313(n988 ,n622 ,n509);
    xnor g314(n2234 ,n41[2] ,n158);
    nand g315(n631 ,n25[7] ,n476);
    nand g316(n1997 ,n1802 ,n1610);
    nand g317(n2043 ,n1871 ,n1653);
    dff g318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2020), .Q(n36[7]));
    nand g319(n384 ,n60[1] ,n331);
    nor g320(n93 ,n40[4] ,n40[3]);
    nor g321(n2167 ,n601 ,n2156);
    or g322(n1109 ,n1036 ,n1051);
    nand g323(n1219 ,n968 ,n757);
    or g324(n1941 ,n1870 ,n1869);
    nand g325(n1128 ,n2237 ,n885);
    nor g326(n369 ,n17[1] ,n336);
    dff g327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2096), .Q(n28[4]));
    dff g328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n291), .Q(n16[10]));
    dff g329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1250), .Q(n40[5]));
    nand g330(n322 ,n37[0] ,n255);
    nand g331(n1149 ,n910 ,n717);
    nand g332(n1208 ,n956 ,n775);
    not g333(n327 ,n328);
    nor g334(n889 ,n252 ,n493);
    nand g335(n949 ,n46[0] ,n568);
    nor g336(n127 ,n60[1] ,n60[0]);
    nand g337(n972 ,n43[4] ,n562);
    nand g338(n1120 ,n38[1] ,n888);
    nand g339(n81 ,n58[1] ,n58[0]);
    nand g340(n1635 ,n39[5] ,n1472);
    nand g341(n1291 ,n1071 ,n824);
    not g342(n1486 ,n1487);
    nand g343(n850 ,n49[2] ,n579);
    nand g344(n1731 ,n27[1] ,n1482);
    nand g345(n780 ,n5[7] ,n557);
    buf g346(n14[2], 1'b0);
    nand g347(n1053 ,n54[0] ,n582);
    nand g348(n1568 ,n50[1] ,n1364);
    nand g349(n2243 ,n115 ,n126);
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2085), .Q(n29[5]));
    nand g351(n1167 ,n848 ,n809);
    nand g352(n790 ,n5[5] ,n557);
    nand g353(n932 ,n47[6] ,n566);
    not g354(n1482 ,n1483);
    nand g355(n882 ,n57[6] ,n553);
    nand g356(n916 ,n51[1] ,n570);
    or g357(n313 ,n62[2] ,n308);
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1231), .Q(n42[4]));
    nor g359(n312 ,n62[2] ,n273);
    dff g360(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1978), .Q(n26[5]));
    nand g361(n2128 ,n518 ,n2116);
    xnor g362(n2216 ,n40[2] ,n143);
    nand g363(n1696 ,n39[2] ,n1491);
    nand g364(n879 ,n20[12] ,n585);
    nand g365(n1336 ,n18[1] ,n1312);
    xnor g366(n2218 ,n40[4] ,n146);
    nand g367(n804 ,n5[7] ,n554);
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1997), .Q(n24[2]));
    nand g369(n1154 ,n61[7] ,n887);
    dff g370(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2022), .Q(n36[5]));
    nand g371(n168 ,n20[2] ,n167);
    nand g372(n1916 ,n2213 ,n1498);
    nand g373(n1304 ,n1063 ,n796);
    nand g374(n2074 ,n837 ,n1910);
    nand g375(n1516 ,n57[7] ,n1362);
    nor g376(n376 ,n219 ,n327);
    nand g377(n1152 ,n913 ,n705);
    nand g378(n1995 ,n1800 ,n1608);
    nand g379(n1883 ,n1449 ,n1574);
    nor g380(n152 ,n40[7] ,n151);
    nand g381(n962 ,n44[6] ,n556);
    nand g382(n1269 ,n396 ,n874);
    nor g383(n137 ,n59[1] ,n59[0]);
    nor g384(n249 ,n19[2] ,n19[3]);
    nand g385(n1758 ,n2190 ,n1499);
    nand g386(n1551 ,n43[0] ,n1363);
    nand g387(n976 ,n43[0] ,n562);
    nand g388(n900 ,n53[0] ,n560);
    nand g389(n2014 ,n1819 ,n1625);
    nor g390(n2229 ,n133 ,n131);
    dff g391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2060), .Q(n31[7]));
    nand g392(n901 ,n52[7] ,n572);
    nand g393(n121 ,n116 ,n120);
    dff g394(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2016), .Q(n21[7]));
    nand g395(n539 ,n29[4] ,n433);
    nand g396(n762 ,n5[2] ,n561);
    nand g397(n1216 ,n1059 ,n755);
    nand g398(n1821 ,n21[7] ,n1495);
    nand g399(n733 ,n5[5] ,n565);
    nand g400(n386 ,n60[3] ,n331);
    nand g401(n185 ,n18[1] ,n18[0]);
    dff g402(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n484), .Q(n39[6]));
    nor g403(n2187 ,n129 ,n127);
    nand g404(n1403 ,n52[3] ,n1368);
    dff g405(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2088), .Q(n29[3]));
    nand g406(n1170 ,n850 ,n813);
    nand g407(n1130 ,n2239 ,n885);
    nand g408(n1530 ,n43[4] ,n1363);
    nor g409(n1352 ,n1099 ,n1098);
    nand g410(n634 ,n2219 ,n421);
    nand g411(n2034 ,n1746 ,n1682);
    nand g412(n1284 ,n1075 ,n808);
    not g413(n1476 ,n1477);
    nand g414(n960 ,n55[1] ,n558);
    nand g415(n1907 ,n30[4] ,n1485);
    dff g416(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1236), .Q(n42[0]));
    nor g417(n1510 ,n193 ,n1389);
    nand g418(n1303 ,n923 ,n795);
    nor g419(n1364 ,n262 ,n1196);
    nand g420(n1902 ,n2205 ,n1498);
    dff g421(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1981), .Q(n26[2]));
    dff g422(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n290), .Q(n16[2]));
    xnor g423(n1361 ,n885 ,n19[0]);
    nand g424(n1828 ,n21[0] ,n1495);
    nand g425(n968 ,n44[0] ,n556);
    nand g426(n1971 ,n1728 ,n1675);
    nand g427(n270 ,n37[0] ,n230);
    nand g428(n722 ,n5[0] ,n569);
    dff g429(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2043), .Q(n34[0]));
    dff g430(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1235), .Q(n42[1]));
    not g431(n1194 ,n1195);
    nand g432(n1856 ,n1412 ,n1442);
    nand g433(n747 ,n5[6] ,n577);
    dff g434(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n483), .Q(n39[4]));
    nand g435(n2114 ,n1119 ,n2099);
    dff g436(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1331), .Q(n58[3]));
    nand g437(n800 ,n339 ,n491);
    nand g438(n714 ,n5[2] ,n571);
    nand g439(n1903 ,n2204 ,n1498);
    nor g440(n436 ,n297 ,n380);
    not g441(n214 ,n40[1]);
    nand g442(n735 ,n5[3] ,n565);
    nand g443(n1963 ,n880 ,n1779);
    dff g444(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1989), .Q(n25[2]));
    nand g445(n855 ,n48[3] ,n563);
    nor g446(n2117 ,n698 ,n1954);
    nand g447(n1338 ,n481 ,n1132);
    nand g448(n680 ,n33[3] ,n434);
    nand g449(n933 ,n47[5] ,n566);
    nor g450(n1719 ,n193 ,n1396);
    nand g451(n1709 ,n39[5] ,n1469);
    or g452(n1099 ,n1014 ,n1012);
    nand g453(n778 ,n5[2] ,n559);
    nand g454(n1672 ,n39[7] ,n1483);
    or g455(n2146 ,n1881 ,n2135);
    not g456(n188 ,n187);
    nor g457(n424 ,n258 ,n403);
    dff g458(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2103), .Q(n21[1]));
    nand g459(n1786 ,n26[2] ,n1475);
    nor g460(n480 ,n205 ,n409);
    dff g461(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1212), .Q(n44[7]));
    nand g462(n1869 ,n1540 ,n1443);
    nor g463(n448 ,n17[1] ,n407);
    nand g464(n753 ,n5[5] ,n555);
    dff g465(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2001), .Q(n23[6]));
    or g466(n1933 ,n1843 ,n1842);
    nand g467(n1030 ,n683 ,n663);
    not g468(n272 ,n271);
    nand g469(n1040 ,n47[0] ,n566);
    nand g470(n2226 ,n84 ,n83);
    nand g471(n1268 ,n945 ,n781);
    nand g472(n301 ,n194 ,n2242);
    dff g473(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1156), .Q(n51[0]));
    nand g474(n918 ,n51[0] ,n570);
    dff g475(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2046), .Q(n33[5]));
    nor g476(n417 ,n17[1] ,n359);
    nand g477(n1647 ,n39[6] ,n1484);
    nand g478(n783 ,n5[5] ,n581);
    nor g479(n1469 ,n298 ,n1378);
    dff g480(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2128), .Q(n12[7]));
    nand g481(n675 ,n24[3] ,n428);
    nand g482(n1654 ,n39[0] ,n1474);
    nand g483(n324 ,n37[2] ,n255);
    nand g484(n1893 ,n32[4] ,n1489);
    nor g485(n290 ,n237 ,n193);
    nor g486(n87 ,n58[2] ,n58[0]);
    nand g487(n693 ,n35[1] ,n435);
    dff g488(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1159), .Q(n50[5]));
    or g489(n595 ,n444 ,n412);
    nand g490(n1258 ,n349 ,n1016);
    dff g491(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2125), .Q(n12[0]));
    not g492(n208 ,n37[3]);
    nand g493(n620 ,n27[2] ,n424);
    nand g494(n1867 ,n34[2] ,n1473);
    dff g495(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1279), .Q(n57[3]));
    nand g496(n1035 ,n53[4] ,n560);
    dff g497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1327), .Q(n60[3]));
    nor g498(n159 ,n37[1] ,n37[0]);
    nand g499(n512 ,n29[0] ,n433);
    nand g500(n2061 ,n1918 ,n1692);
    nand g501(n1881 ,n1448 ,n1569);
    nand g502(n810 ,n5[6] ,n580);
    nand g503(n1610 ,n39[2] ,n1478);
    nand g504(n515 ,n22[7] ,n423);
    buf g505(n16[11], 1'b0);
    nand g506(n519 ,n31[0] ,n427);
    nand g507(n1632 ,n39[1] ,n1494);
    dff g508(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1299), .Q(n55[0]));
    nor g509(n367 ,n316 ,n311);
    nand g510(n801 ,n5[6] ,n554);
    nand g511(n1743 ,n35[5] ,n1492);
    not g512(n441 ,n442);
    nand g513(n2071 ,n868 ,n1903);
    not g514(n114 ,n20[5]);
    not g515(n1484 ,n1485);
    dff g516(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1172), .Q(n49[0]));
    nand g517(n1572 ,n55[5] ,n1370);
    nand g518(n1840 ,n1561 ,n1265);
    nor g519(n334 ,n208 ,n301);
    nand g520(n1887 ,n1552 ,n1455);
    nand g521(n1676 ,n39[3] ,n1483);
    nand g522(n1910 ,n2203 ,n1498);
    nand g523(n2098 ,n2198 ,n1755);
    nand g524(n1564 ,n53[5] ,n1375);
    nor g525(n1385 ,n418 ,n1103);
    xnor g526(n2223 ,n40[9] ,n155);
    nand g527(n2033 ,n1747 ,n1681);
    nor g528(n1345 ,n275 ,n1309);
    dff g529(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2002), .Q(n23[5]));
    nand g530(n1526 ,n56[5] ,n1377);
    nand g531(n745 ,n5[7] ,n577);
    nand g532(n1270 ,n61[2] ,n887);
    nor g533(n293 ,n209 ,n213);
    nand g534(n1617 ,n39[2] ,n1480);
    not g535(n559 ,n560);
    not g536(n1088 ,n1002);
    nand g537(n122 ,n20[6] ,n121);
    nor g538(n412 ,n276 ,n393);
    nand g539(n1863 ,n34[3] ,n1473);
    nor g540(n256 ,n62[0] ,n62[1]);
    nand g541(n459 ,n40[6] ,n378);
    nand g542(n2052 ,n1886 ,n1639);
    nand g543(n826 ,n5[7] ,n576);
    nand g544(n1243 ,n41[1] ,n890);
    buf g545(n16[13], 1'b0);
    nor g546(n1341 ,n193 ,n1125);
    nand g547(n2127 ,n505 ,n2115);
    nor g548(n554 ,n300 ,n479);
    not g549(n1381 ,n1382);
    dff g550(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n285), .Q(n16[1]));
    nand g551(n730 ,n5[1] ,n583);
    nand g552(n1319 ,n1129 ,n1261);
    nand g553(n740 ,n5[5] ,n567);
    not g554(n244 ,n40[8]);
    nand g555(n1680 ,n39[4] ,n1493);
    nand g556(n1215 ,n964 ,n754);
    nand g557(n1289 ,n1072 ,n830);
    nor g558(n171 ,n163 ,n170);
    nand g559(n1238 ,n915 ,n776);
    nand g560(n819 ,n5[4] ,n564);
    not g561(n197 ,n39[1]);
    or g562(n1112 ,n221 ,n894);
    nand g563(n1576 ,n44[5] ,n1366);
    nand g564(n1033 ,n53[5] ,n560);
    xnor g565(n2237 ,n79 ,n19[4]);
    or g566(n1931 ,n1912 ,n1840);
    nand g567(n1917 ,n2201 ,n1498);
    nand g568(n1767 ,n29[4] ,n1470);
    nand g569(n184 ,n20[11] ,n183);
    dff g570(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n485), .Q(n39[5]));
    nand g571(n1694 ,n39[4] ,n1491);
    nand g572(n709 ,n5[5] ,n571);
    nand g573(n724 ,n5[7] ,n573);
    not g574(n697 ,n652);
    nand g575(n2183 ,n2243 ,n2182);
    nand g576(n2069 ,n1762 ,n1698);
    nand g577(n1333 ,n18[2] ,n1312);
    nand g578(n2178 ,n1549 ,n2170);
    nand g579(n1686 ,n39[3] ,n1493);
    dff g580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1221), .Q(n43[6]));
    dff g581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1171), .Q(n49[1]));
    nor g582(n178 ,n164 ,n177);
    nand g583(n1571 ,n54[5] ,n1373);
    nand g584(n522 ,n23[6] ,n429);
    nand g585(n521 ,n22[6] ,n423);
    dff g586(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2034), .Q(n35[2]));
    nand g587(n2210 ,n104 ,n113);
    nand g588(n744 ,n5[0] ,n567);
    nand g589(n997 ,n459 ,n632);
    nor g590(n1397 ,n1346 ,n1343);
    dff g591(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1252), .Q(n40[3]));
    nand g592(n955 ,n615 ,n544);
    or g593(n105 ,n20[3] ,n20[2]);
    nand g594(n1831 ,n1538 ,n1573);
    nand g595(n1022 ,n51[3] ,n570);
    nand g596(n1136 ,n1033 ,n703);
    nor g597(n2111 ,n1945 ,n1944);
    dff g598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2013), .Q(n22[2]));
    nand g599(n1427 ,n53[6] ,n1375);
    nand g600(n560 ,n269 ,n480);
    buf g601(n16[15], 1'b0);
    nand g602(n1077 ,n57[2] ,n553);
    nand g603(n1574 ,n52[1] ,n1368);
    dff g604(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1183), .Q(n47[6]));
    nand g605(n755 ,n5[3] ,n555);
    nand g606(n1503 ,n48[3] ,n1367);
    nand g607(n1207 ,n954 ,n748);
    dff g608(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1241), .Q(n57[6]));
    nand g609(n347 ,n17[0] ,n303);
    nand g610(n671 ,n25[2] ,n476);
    nand g611(n2125 ,n533 ,n2118);
    nand g612(n781 ,n5[3] ,n567);
    nand g613(n1181 ,n858 ,n823);
    nand g614(n1837 ,n1555 ,n1424);
    nor g615(n427 ,n258 ,n380);
    dff g616(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1177), .Q(n48[4]));
    nand g617(n2075 ,n1906 ,n1648);
    nand g618(n546 ,n22[1] ,n423);
    nand g619(n1192 ,n942 ,n740);
    nand g620(n821 ,n5[3] ,n564);
    nand g621(n1311 ,n194 ,n1080);
    nand g622(n1962 ,n1723 ,n1671);
    nand g623(n1895 ,n32[3] ,n1489);
    nand g624(n309 ,n2243 ,n221);
    nand g625(n2148 ,n1928 ,n2140);
    dff g626(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2176), .Q(n61[3]));
    not g627(n1085 ,n997);
    nor g628(n278 ,n193 ,n58[0]);
    nand g629(n759 ,n5[6] ,n561);
    nand g630(n1433 ,n44[6] ,n1366);
    nand g631(n1979 ,n1784 ,n1593);
    nand g632(n1909 ,n30[2] ,n1485);
    nor g633(n2241 ,n19[4] ,n191);
    nand g634(n1810 ,n23[2] ,n1481);
    nand g635(n685 ,n32[3] ,n436);
    dff g636(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1995), .Q(n24[4]));
    buf g637(n1499 ,n587);
    dff g638(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2172), .Q(n61[6]));
    nand g639(n2097 ,n1776 ,n1711);
    nand g640(n604 ,n32[4] ,n436);
    dff g641(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2055), .Q(n32[4]));
    nand g642(n527 ,n21[3] ,n430);
    nand g643(n1848 ,n1528 ,n1437);
    nand g644(n803 ,n5[2] ,n554);
    not g645(n1488 ,n1489);
    nor g646(n2116 ,n696 ,n1952);
    nor g647(n358 ,n257 ,n337);
    nand g648(n1645 ,n39[1] ,n1488);
    nand g649(n1789 ,n25[7] ,n1477);
    xnor g650(n2192 ,n59[3] ,n140);
    nand g651(n550 ,n29[2] ,n433);
    not g652(n156 ,n155);
    nand g653(n1292 ,n1024 ,n780);
    nand g654(n304 ,n14[1] ,n194);
    nand g655(n1959 ,n840 ,n1757);
    nand g656(n1032 ,n525 ,n552);
    nand g657(n1911 ,n30[1] ,n1485);
    dff g658(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1975), .Q(n27[0]));
    nand g659(n1058 ,n614 ,n664);
    nand g660(n1143 ,n1067 ,n709);
    nor g661(n2154 ,n1946 ,n2146);
    nor g662(n319 ,n17[0] ,n309);
    nand g663(n1624 ,n39[2] ,n1496);
    not g664(n195 ,n39[5]);
    nand g665(n1132 ,n353 ,n800);
    nand g666(n627 ,n33[1] ,n434);
    nand g667(n1621 ,n39[6] ,n1496);
    nand g668(n1861 ,n1503 ,n1439);
    nand g669(n306 ,n4 ,n233);
    not g670(n444 ,n443);
    nand g671(n1922 ,n33[2] ,n1486);
    nand g672(n993 ,n470 ,n682);
    nand g673(n1900 ,n2206 ,n1498);
    nand g674(n532 ,n29[3] ,n433);
    nand g675(n625 ,n27[0] ,n424);
    nand g676(n906 ,n52[1] ,n572);
    nand g677(n654 ,n34[6] ,n426);
    dff g678(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1259), .Q(n37[2]));
    nand g679(n1475 ,n260 ,n1379);
    nand g680(n545 ,n22[3] ,n423);
    nor g681(n2110 ,n1942 ,n1941);
    nand g682(n1998 ,n1803 ,n1611);
    nand g683(n1718 ,n39[0] ,n1471);
    nand g684(n1650 ,n39[3] ,n1484);
    nor g685(n282 ,n215 ,n192);
    not g686(n260 ,n259);
    nor g687(n289 ,n244 ,n193);
    not g688(n437 ,n438);
    nor g689(n251 ,n58[2] ,n58[3]);
    nand g690(n1993 ,n1798 ,n1606);
    nand g691(n676 ,n394 ,n474);
    nor g692(n2170 ,n600 ,n2163);
    nand g693(n1683 ,n39[7] ,n1487);
    not g694(n1089 ,n1003);
    nand g695(n782 ,n5[6] ,n557);
    nand g696(n1056 ,n55[4] ,n558);
    nand g697(n1822 ,n21[6] ,n1495);
    nand g698(n1570 ,n52[6] ,n1368);
    dff g699(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1307), .Q(n53[7]));
    or g700(n1943 ,n1876 ,n1875);
    nor g701(n454 ,n361 ,n372);
    nand g702(n1631 ,n39[2] ,n1494);
    nand g703(n2030 ,n1743 ,n1691);
    nor g704(n1374 ,n261 ,n1198);
    nand g705(n683 ,n26[4] ,n431);
    not g706(n63 ,n19[3]);
    nand g707(n1629 ,n39[4] ,n1494);
    nor g708(n2182 ,n18[0] ,n2179);
    nand g709(n1638 ,n39[1] ,n1472);
    dff g710(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1721), .Q(n62[1]));
    nand g711(n825 ,n5[2] ,n564);
    nand g712(n1921 ,n33[1] ,n1486);
    not g713(n1087 ,n1000);
    nor g714(n430 ,n268 ,n401);
    nand g715(n1793 ,n25[3] ,n1477);
    nand g716(n841 ,n58[4] ,n589);
    not g717(n135 ,n134);
    nand g718(n1832 ,n1536 ,n1422);
    nand g719(n1237 ,n834 ,n987);
    nand g720(n915 ,n51[2] ,n570);
    nand g721(n1068 ,n685 ,n680);
    nand g722(n2031 ,n1744 ,n1680);
    nand g723(n1690 ,n39[7] ,n1491);
    nand g724(n1844 ,n1572 ,n1571);
    nand g725(n930 ,n502 ,n510);
    not g726(n1468 ,n1469);
    nand g727(n568 ,n264 ,n442);
    nand g728(n506 ,n31[3] ,n427);
    not g729(n305 ,n304);
    not g730(n563 ,n564);
    nand g731(n1039 ,n46[6] ,n568);
    not g732(n181 ,n180);
    nand g733(n1183 ,n932 ,n732);
    nand g734(n835 ,n223 ,n595);
    nand g735(n725 ,n5[5] ,n573);
    nand g736(n746 ,n5[0] ,n557);
    nor g737(n1247 ,n192 ,n1081);
    not g738(n215 ,n40[7]);
    nand g739(n1841 ,n1560 ,n1429);
    nand g740(n721 ,n5[3] ,n569);
    nor g741(n489 ,n40[0] ,n420);
    nand g742(n2131 ,n536 ,n2120);
    nand g743(n1787 ,n26[1] ,n1475);
    nand g744(n705 ,n5[4] ,n569);
    nand g745(n1892 ,n1458 ,n1457);
    nand g746(n728 ,n5[1] ,n573);
    nand g747(n1875 ,n1543 ,n1270);
    or g748(n1092 ,n988 ,n983);
    nor g749(n1359 ,n313 ,n1194);
    nand g750(n964 ,n44[4] ,n556);
    nand g751(n1816 ,n22[4] ,n1497);
    dff g752(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1293), .Q(n55[6]));
    nand g753(n1693 ,n39[5] ,n1491);
    nor g754(n1398 ,n1344 ,n1359);
    nand g755(n180 ,n20[9] ,n178);
    nand g756(n951 ,n45[6] ,n578);
    dff g757(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1169), .Q(n49[3]));
    nand g758(n77 ,n74 ,n71);
    not g759(n222 ,n62[2]);
    dff g760(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1208), .Q(n45[3]));
    nand g761(n611 ,n24[1] ,n428);
    nand g762(n2160 ,n1434 ,n2155);
    not g763(n567 ,n568);
    dff g764(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2035), .Q(n35[0]));
    nand g765(n618 ,n35[4] ,n435);
    dff g766(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2049), .Q(n33[2]));
    nand g767(n1294 ,n1055 ,n790);
    nand g768(n1858 ,n1535 ,n1409);
    nand g769(n1072 ,n56[3] ,n575);
    nand g770(n622 ,n24[0] ,n428);
    dff g771(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1961), .Q(n28[2]));
    dff g772(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1188), .Q(n47[1]));
    nand g773(n1241 ,n882 ,n801);
    dff g774(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2045), .Q(n33[6]));
    nor g775(n1125 ,n836 ,n897);
    nand g776(n2102 ,n1826 ,n1631);
    nand g777(n1842 ,n1525 ,n1575);
    nand g778(n797 ,n5[2] ,n581);
    nand g779(n1595 ,n39[2] ,n1474);
    nand g780(n533 ,n30[0] ,n425);
    dff g781(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1342), .Q(n41[0]));
    buf g782(n893 ,n330);
    nand g783(n921 ,n50[3] ,n574);
    nand g784(n1612 ,n39[7] ,n1480);
    nand g785(n157 ,n40[9] ,n156);
    not g786(n577 ,n578);
    nand g787(n175 ,n20[6] ,n174);
    nand g788(n1459 ,n52[0] ,n1368);
    nor g789(n2109 ,n1939 ,n1938);
    nor g790(n273 ,n232 ,n62[0]);
    nand g791(n1461 ,n318 ,n1351);
    nand g792(n146 ,n40[3] ,n144);
    nand g793(n860 ,n59[3] ,n592);
    nand g794(n1681 ,n39[1] ,n1493);
    nand g795(n1599 ,n39[6] ,n1476);
    nor g796(n2199 ,n167 ,n165);
    dff g797(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2070), .Q(n31[0]));
    nand g798(n1843 ,n1558 ,n1419);
    nand g799(n1285 ,n1074 ,n826);
    nor g800(n1754 ,n192 ,n1393);
    nand g801(n792 ,n5[3] ,n557);
    nand g802(n1782 ,n26[6] ,n1475);
    nand g803(n710 ,n5[6] ,n571);
    nor g804(n111 ,n106 ,n110);
    nand g805(n786 ,n5[7] ,n559);
    or g806(n834 ,n222 ,n596);
    or g807(n2142 ,n1844 ,n2139);
    nand g808(n357 ,n223 ,n342);
    nand g809(n1546 ,n48[1] ,n1367);
    nand g810(n629 ,n24[7] ,n428);
    nand g811(n99 ,n40[6] ,n98);
    nand g812(n1559 ,n57[0] ,n1362);
    nand g813(n1436 ,n53[4] ,n1375);
    dff g814(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2121), .Q(n38[1]));
    dff g815(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1222), .Q(n43[5]));
    nand g816(n975 ,n43[1] ,n562);
    nand g817(n1797 ,n24[7] ,n1479);
    nand g818(n258 ,n37[1] ,n224);
    nand g819(n582 ,n264 ,n440);
    not g820(n68 ,n67);
    nand g821(n380 ,n229 ,n334);
    not g822(n439 ,n440);
    nand g823(n1974 ,n1731 ,n1678);
    or g824(n2244 ,n40[10] ,n102);
    nor g825(n126 ,n20[12] ,n125);
    nand g826(n902 ,n547 ,n497);
    dff g827(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1190), .Q(n46[7]));
    xnor g828(n2200 ,n20[3] ,n168);
    nor g829(n172 ,n20[5] ,n171);
    or g830(n103 ,n20[1] ,n20[0]);
    nand g831(n923 ,n54[4] ,n582);
    nor g832(n414 ,n19[4] ,n405);
    nand g833(n1323 ,n1112 ,n1244);
    dff g834(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1225), .Q(n43[2]));
    not g835(n174 ,n173);
    not g836(n1925 ,n1829);
    nand g837(n1573 ,n44[7] ,n1366);
    nand g838(n547 ,n22[2] ,n423);
    nand g839(n1458 ,n55[0] ,n1370);
    nand g840(n1835 ,n1517 ,n1462);
    nand g841(n1994 ,n1799 ,n1607);
    dff g842(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1251), .Q(n40[4]));
    nand g843(n1142 ,n909 ,n710);
    nand g844(n938 ,n611 ,n529);
    nand g845(n1805 ,n23[7] ,n1481);
    nand g846(n1232 ,n982 ,n770);
    dff g847(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1291), .Q(n56[1]));
    dff g848(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1971), .Q(n27[4]));
    nand g849(n1147 ,n906 ,n715);
    nand g850(n1692 ,n39[6] ,n1491);
    nand g851(n1860 ,n1504 ,n1407);
    nand g852(n566 ,n264 ,n438);
    not g853(n378 ,n379);
    nand g854(n138 ,n59[1] ,n59[0]);
    not g855(n1317 ,n1275);
    nand g856(n1443 ,n42[2] ,n1376);
    nand g857(n1328 ,n389 ,n1134);
    not g858(n1480 ,n1481);
    nand g859(n1829 ,n194 ,n1512);
    or g860(n400 ,n205 ,n329);
    buf g861(n14[6], 1'b0);
    nor g862(n2190 ,n139 ,n137);
    nand g863(n1162 ,n922 ,n772);
    dff g864(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1141), .Q(n52[7]));
    nor g865(n1396 ,n1348 ,n1345);
    nand g866(n1603 ,n39[2] ,n1476);
    or g867(n1127 ,n907 ,n902);
    nand g868(n827 ,n5[6] ,n576);
    dff g869(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2033), .Q(n35[1]));
    not g870(n1389 ,n1320);
    dff g871(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2097), .Q(n28[3]));
    nand g872(n513 ,n23[7] ,n429);
    or g873(n1944 ,n1878 ,n1877);
    nand g874(n2012 ,n1817 ,n1623);
    nand g875(n617 ,n36[1] ,n422);
    nand g876(n1463 ,n51[0] ,n1365);
    nand g877(n1422 ,n46[7] ,n1374);
    nand g878(n833 ,n278 ,n588);
    nand g879(n2089 ,n847 ,n1917);
    nor g880(n379 ,n345 ,n333);
    nand g881(n1437 ,n44[4] ,n1366);
    xnor g882(n2206 ,n184 ,n20[12]);
    nand g883(n1542 ,n56[2] ,n1377);
    xnor g884(n2230 ,n58[2] ,n132);
    dff g885(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2082), .Q(n29[7]));
    nand g886(n1025 ,n661 ,n679);
    dff g887(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2061), .Q(n31[6]));
    buf g888(n14[5], 1'b0);
    nand g889(n994 ,n625 ,n512);
    nand g890(n1282 ,n1076 ,n807);
    nand g891(n1536 ,n47[7] ,n1371);
    nand g892(n1400 ,n44[2] ,n1366);
    nand g893(n1532 ,n49[4] ,n1369);
    not g894(n2186 ,n1);
    nand g895(n845 ,n49[6] ,n579);
    or g896(n112 ,n20[12] ,n111);
    not g897(n573 ,n574);
    nand g898(n299 ,n59[1] ,n59[2]);
    nand g899(n1218 ,n967 ,n788);
    not g900(n1383 ,n1384);
    dff g901(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1139), .Q(n53[1]));
    nand g902(n1882 ,n1548 ,n1283);
    nor g903(n1251 ,n193 ,n1087);
    not g904(n161 ,n160);
    nor g905(n446 ,n222 ,n358);
    nand g906(n1210 ,n957 ,n750);
    nor g907(n296 ,n211 ,n192);
    not g908(n192 ,n194);
    nand g909(n1069 ,n2228 ,n587);
    nand g910(n1430 ,n50[4] ,n1364);
    nand g911(n681 ,n36[5] ,n422);
    nand g912(n752 ,n5[6] ,n555);
    nor g913(n2151 ,n1931 ,n2141);
    nand g914(n1050 ,n2225 ,n587);
    nand g915(n1435 ,n54[4] ,n1373);
    nand g916(n847 ,n20[5] ,n585);
    nand g917(n1630 ,n39[3] ,n1494);
    nand g918(n818 ,n5[5] ,n564);
    nand g919(n1833 ,n1414 ,n1423);
    nand g920(n552 ,n21[4] ,n430);
    nand g921(n630 ,n2222 ,n421);
    nand g922(n2029 ,n1742 ,n1697);
    xnor g923(n2232 ,n136 ,n58[4]);
    nand g924(n1981 ,n1786 ,n1595);
    nor g925(n452 ,n233 ,n408);
    nand g926(n1815 ,n22[5] ,n1497);
    nor g927(n487 ,n193 ,n451);
    nor g928(n245 ,n199 ,n221);
    nor g929(n1377 ,n299 ,n1196);
    nand g930(n832 ,n5[0] ,n576);
    nand g931(n1070 ,n53[6] ,n560);
    nand g932(n607 ,n28[3] ,n432);
    or g933(n1934 ,n1846 ,n1845);
    nor g934(n374 ,n217 ,n327);
    nand g935(n655 ,n35[6] ,n435);
    not g936(n183 ,n182);
    nand g937(n953 ,n45[5] ,n578);
    nand g938(n2156 ,n1428 ,n2151);
    dff g939(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n486), .Q(n39[3]));
    nand g940(n1990 ,n1795 ,n1604);
    nand g941(n1616 ,n39[3] ,n1480);
    nand g942(n708 ,n5[0] ,n559);
    nand g943(n492 ,n222 ,n455);
    nor g944(n836 ,n62[2] ,n594);
    or g945(n2143 ,n1892 ,n2136);
    nand g946(n382 ,n194 ,n317);
    nand g947(n1798 ,n24[6] ,n1479);
    nor g948(n428 ,n297 ,n401);
    nand g949(n946 ,n46[2] ,n568);
    nand g950(n1416 ,n354 ,n1353);
    nand g951(n637 ,n34[7] ,n426);
    nand g952(n1865 ,n1537 ,n1176);
    dff g953(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n419), .Q(n60[0]));
    nand g954(n398 ,n2232 ,n330);
    nand g955(n990 ,n653 ,n623);
    nor g956(n82 ,n58[2] ,n80);
    nand g957(n1259 ,n324 ,n1017);
    nor g958(n288 ,n216 ,n193);
    nand g959(n984 ,n42[2] ,n584);
    nor g960(n1349 ,n1105 ,n1109);
    nand g961(n1710 ,n39[4] ,n1469);
    nand g962(n551 ,n61[4] ,n475);
    nand g963(n1538 ,n45[7] ,n1372);
    nand g964(n534 ,n29[5] ,n433);
    nand g965(n1042 ,n667 ,n528);
    nand g966(n1453 ,n348 ,n1350);
    nand g967(n1556 ,n49[0] ,n1369);
    nor g968(n113 ,n20[9] ,n112);
    nand g969(n1455 ,n46[0] ,n1374);
    nand g970(n777 ,n5[7] ,n581);
    buf g971(n15[4], n13[2]);
    nand g972(n1462 ,n42[6] ,n1376);
    nand g973(n540 ,n61[2] ,n475);
    nand g974(n516 ,n31[7] ,n427);
    nand g975(n1060 ,n54[6] ,n582);
    nand g976(n252 ,n194 ,n2244);
    nand g977(n904 ,n52[3] ,n572);
    nor g978(n292 ,n210 ,n193);
    nand g979(n1627 ,n39[6] ,n1494);
    nand g980(n415 ,n222 ,n381);
    xor g981(n2233 ,n41[1] ,n41[0]);
    nand g982(n768 ,n5[5] ,n583);
    or g983(n1930 ,n1838 ,n1837);
    xnor g984(n2231 ,n58[3] ,n134);
    dff g985(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2029), .Q(n35[6]));
    nor g986(n343 ,n17[0] ,n276);
    nor g987(n91 ,n19[3] ,n89);
    nand g988(n1765 ,n29[6] ,n1470);
    nand g989(n1725 ,n27[7] ,n1482);
    nor g990(n475 ,n202 ,n382);
    nand g991(n820 ,n5[7] ,n580);
    nand g992(n526 ,n30[5] ,n425);
    nand g993(n1745 ,n35[3] ,n1492);
    nand g994(n1005 ,n640 ,n637);
    nand g995(n499 ,n31[2] ,n427);
    nand g996(n1504 ,n47[3] ,n1371);
    dff g997(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2064), .Q(n31[5]));
    nand g998(n1620 ,n39[5] ,n1496);
    nand g999(n857 ,n48[1] ,n563);
    nand g1000(n1059 ,n44[3] ,n556);
    nand g1001(n302 ,n2243 ,n223);
    xor g1002(n2227 ,n58[3] ,n82);
    or g1003(n1107 ,n1047 ,n1028);
    nand g1004(n2072 ,n1904 ,n1646);
    nor g1005(n1100 ,n1013 ,n1009);
    nand g1006(n791 ,n5[4] ,n557);
    nand g1007(n1590 ,n39[7] ,n1474);
    nand g1008(n1814 ,n22[6] ,n1497);
    nand g1009(n1885 ,n1550 ,n1452);
    nor g1010(n432 ,n297 ,n403);
    dff g1011(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1720), .Q(n17[0]));
    nand g1012(n543 ,n23[3] ,n429);
    nand g1013(n549 ,n61[5] ,n475);
    dff g1014(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2092), .Q(n29[0]));
    nand g1015(n1608 ,n39[4] ,n1478);
    nand g1016(n170 ,n20[3] ,n169);
    xnor g1017(n2224 ,n40[10] ,n157);
    nand g1018(n1622 ,n39[4] ,n1496);
    nand g1019(n1129 ,n2238 ,n885);
    nand g1020(n1062 ,n54[5] ,n582);
    nand g1021(n798 ,n5[0] ,n581);
    nand g1022(n1044 ,n609 ,n542);
    nand g1023(n396 ,n2229 ,n330);
    dff g1024(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1719), .Q(n17[2]));
    nand g1025(n1853 ,n1532 ,n1264);
    nor g1026(n2193 ,n161 ,n159);
    nand g1027(n2073 ,n1905 ,n1647);
    nand g1028(n1716 ,n39[0] ,n1487);
    nand g1029(n1794 ,n25[2] ,n1477);
    nand g1030(n1888 ,n1553 ,n1456);
    nand g1031(n497 ,n21[2] ,n430);
    nand g1032(n1144 ,n903 ,n712);
    nor g1033(n456 ,n364 ,n373);
    dff g1034(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2050), .Q(n33[1]));
    or g1035(n314 ,n37[0] ,n301);
    nand g1036(n1954 ,n1101 ,n1585);
    dff g1037(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2065), .Q(n31[4]));
    nand g1038(n1281 ,n1077 ,n803);
    not g1039(n897 ,n862);
    nand g1040(n1723 ,n28[1] ,n1468);
    nor g1041(n442 ,n60[3] ,n404);
    nand g1042(n1429 ,n42[5] ,n1376);
    nand g1043(n987 ,n8 ,n596);
    or g1044(n80 ,n58[1] ,n58[0]);
    nand g1045(n1968 ,n1726 ,n1673);
    nor g1046(n887 ,n475 ,n591);
    nor g1047(n345 ,n222 ,n256);
    dff g1048(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1209), .Q(n45[2]));
    not g1049(n141 ,n40[6]);
    nand g1050(n578 ,n269 ,n438);
    nand g1051(n1271 ,n61[0] ,n887);
    dff g1052(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2178), .Q(n61[1]));
    nor g1053(n1508 ,n192 ,n1387);
    dff g1054(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1230), .Q(n42[5]));
    nand g1055(n875 ,n56[6] ,n575);
    nor g1056(n1113 ,n192 ,n884);
    nand g1057(n1211 ,n959 ,n787);
    not g1058(n213 ,n18[2]);
    nand g1059(n1420 ,n52[4] ,n1368);
    nand g1060(n469 ,n40[10] ,n378);
    nand g1061(n1555 ,n47[6] ,n1371);
    nand g1062(n1771 ,n29[0] ,n1470);
    nand g1063(n2240 ,n70 ,n75);
    nor g1064(n1110 ,n1068 ,n1065);
    nand g1065(n2079 ,n1911 ,n1652);
    nand g1066(n899 ,n53[2] ,n560);
    nand g1067(n1744 ,n35[4] ,n1492);
    nand g1068(n741 ,n5[4] ,n567);
    nor g1069(n337 ,n41[1] ,n248);
    nand g1070(n839 ,n59[1] ,n592);
    not g1071(n1081 ,n989);
    nand g1072(n908 ,n52[0] ,n572);
    nand g1073(n1063 ,n54[3] ,n582);
    nand g1074(n155 ,n40[8] ,n154);
    nand g1075(n927 ,n606 ,n624);
    nand g1076(n2023 ,n1736 ,n1666);
    or g1077(n401 ,n37[2] ,n341);
    nand g1078(n1898 ,n32[1] ,n1489);
    dff g1079(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n487), .Q(n39[1]));
    nand g1080(n1729 ,n27[3] ,n1482);
    nor g1081(n1588 ,n1015 ,n1461);
    nor g1082(n109 ,n107 ,n108);
    nand g1083(n1038 ,n668 ,n539);
    nand g1084(n2048 ,n1923 ,n1707);
    nand g1085(n1784 ,n26[4] ,n1475);
    nand g1086(n2007 ,n1812 ,n1657);
    dff g1087(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1167), .Q(n49[5]));
    nand g1088(n911 ,n51[6] ,n570);
    nand g1089(n1852 ,n34[7] ,n1473);
    nand g1090(n717 ,n5[7] ,n569);
    nand g1091(n1450 ,n51[1] ,n1365);
    not g1092(n1312 ,n1311);
    nand g1093(n1206 ,n953 ,n743);
    nand g1094(n74 ,n19[2] ,n67);
    nand g1095(n1984 ,n1789 ,n1597);
    nand g1096(n2122 ,n1118 ,n2098);
    nor g1097(n64 ,n19[1] ,n19[0]);
    nand g1098(n1045 ,n53[7] ,n560);
    dff g1099(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2003), .Q(n23[4]));
    dff g1100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1192), .Q(n46[5]));
    or g1101(n2179 ,n18[2] ,n18[1]);
    nand g1102(n182 ,n20[10] ,n181);
    not g1103(n1083 ,n993);
    nand g1104(n275 ,n17[1] ,n221);
    nand g1105(n1918 ,n31[6] ,n1490);
    not g1106(n219 ,n39[2]);
    nand g1107(n2010 ,n1815 ,n1620);
    nand g1108(n1752 ,n33[6] ,n1486);
    nand g1109(n1234 ,n984 ,n771);
    nand g1110(n2172 ,n1523 ,n2167);
    nand g1111(n1577 ,n48[4] ,n1367);
    nand g1112(n1961 ,n1722 ,n1670);
    nand g1113(n658 ,n32[6] ,n436);
    nand g1114(n1254 ,n947 ,n779);
    nand g1115(n865 ,n57[7] ,n553);
    nand g1116(n769 ,n5[4] ,n583);
    dff g1117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2175), .Q(n61[0]));
    nand g1118(n1761 ,n31[2] ,n1490);
    dff g1119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1152), .Q(n51[4]));
    nand g1120(n562 ,n263 ,n438);
    nor g1121(n886 ,n2242 ,n590);
    nand g1122(n1539 ,n57[3] ,n1362);
    nor g1123(n1122 ,n1046 ,n1044);
    nand g1124(n1544 ,n45[1] ,n1372);
    nand g1125(n128 ,n60[1] ,n60[0]);
    nand g1126(n468 ,n2243 ,n357);
    nand g1127(n1412 ,n53[7] ,n1375);
    dff g1128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1321), .Q(n60[1]));
    nand g1129(n1332 ,n1069 ,n1315);
    nand g1130(n742 ,n5[2] ,n567);
    nand g1131(n1915 ,n2202 ,n1498);
    nand g1132(n2176 ,n1539 ,n2168);
    dff g1133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1329), .Q(n58[1]));
    nand g1134(n985 ,n42[1] ,n584);
    nand g1135(n1563 ,n43[1] ,n1363);
    dff g1136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1246), .Q(n40[9]));
    dff g1137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2072), .Q(n30[7]));
    nand g1138(n711 ,n5[7] ,n571);
    nand g1139(n584 ,n263 ,n442);
    nand g1140(n670 ,n36[3] ,n422);
    nand g1141(n1300 ,n936 ,n777);
    nand g1142(n1157 ,n1037 ,n724);
    nand g1143(n495 ,n221 ,n468);
    nand g1144(n410 ,n347 ,n356);
    nand g1145(n1989 ,n1794 ,n1603);
    nand g1146(n397 ,n2231 ,n330);
    not g1147(n555 ,n556);
    nor g1148(n2120 ,n702 ,n1956);
    nand g1149(n1992 ,n1797 ,n1605);
    nor g1150(n2118 ,n697 ,n1953);
    nand g1151(n1118 ,n38[3] ,n888);
    nor g1152(n440 ,n60[0] ,n409);
    nand g1153(n1175 ,n872 ,n818);
    nor g1154(n1721 ,n192 ,n1398);
    nand g1155(n959 ,n45[0] ,n578);
    nand g1156(n823 ,n5[0] ,n564);
    nand g1157(n523 ,n29[6] ,n433);
    nand g1158(n995 ,n629 ,n513);
    or g1159(n1937 ,n1854 ,n1853);
    nand g1160(n2040 ,n1863 ,n1637);
    nor g1161(n88 ,n58[3] ,n86);
    nor g1162(n1356 ,n1123 ,n1127);
    nand g1163(n420 ,n202 ,n379);
    nand g1164(n2035 ,n1749 ,n1715);
    nand g1165(n856 ,n48[2] ,n563);
    nand g1166(n1145 ,n904 ,n713);
    nor g1167(n2221 ,n152 ,n154);
    nand g1168(n941 ,n55[0] ,n558);
    nor g1169(n363 ,n217 ,n328);
    nor g1170(n1399 ,n192 ,n1340);
    nand g1171(n1666 ,n39[4] ,n1467);
    nand g1172(n1277 ,n865 ,n804);
    nand g1173(n1965 ,n873 ,n1777);
    not g1174(n235 ,n41[1]);
    nand g1175(n1121 ,n19[4] ,n886);
    nor g1176(n1354 ,n1095 ,n1092);
    nand g1177(n2096 ,n1775 ,n1710);
    nor g1178(n2168 ,n603 ,n2157);
    not g1179(n892 ,n891);
    nand g1180(n1080 ,n370 ,n666);
    nor g1181(n457 ,n377 ,n388);
    nand g1182(n308 ,n62[0] ,n232);
    not g1183(n210 ,n40[5]);
    or g1184(n1938 ,n1858 ,n1857);
    nand g1185(n1924 ,n1518 ,n1433);
    nor g1186(n590 ,n19[4] ,n443);
    not g1187(n581 ,n582);
    nand g1188(n612 ,n25[1] ,n476);
    nand g1189(n1065 ,n607 ,n506);
    nand g1190(n510 ,n21[5] ,n430);
    dff g1191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2075), .Q(n30[5]));
    nand g1192(n771 ,n5[2] ,n583);
    nand g1193(n2136 ,n1554 ,n2112);
    dff g1194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1213), .Q(n44[6]));
    dff g1195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1166), .Q(n49[6]));
    dff g1196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2089), .Q(n20[5]));
    nand g1197(n1244 ,n9 ,n894);
    nand g1198(n2158 ,n1413 ,n2149);
    nand g1199(n1640 ,n39[6] ,n1488);
    nand g1200(n1641 ,n39[5] ,n1488);
    dff g1201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1970), .Q(n20[3]));
    dff g1202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1249), .Q(n40[6]));
    nand g1203(n1031 ,n2226 ,n587);
    nand g1204(n1727 ,n27[5] ,n1482);
    nor g1205(n78 ,n63 ,n74);
    nand g1206(n1670 ,n39[2] ,n1469);
    or g1207(n1093 ,n948 ,n944);
    nand g1208(n1643 ,n39[3] ,n1488);
    nand g1209(n1442 ,n52[7] ,n1368);
    nand g1210(n776 ,n5[2] ,n569);
    dff g1211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1191), .Q(n46[6]));
    buf g1212(n15[0], 1'b0);
    nand g1213(n1567 ,n351 ,n1349);
    nand g1214(n1541 ,n47[2] ,n1371);
    nand g1215(n1428 ,n51[6] ,n1365);
    nand g1216(n1819 ,n22[1] ,n1497);
    not g1217(n885 ,n886);
    nand g1218(n751 ,n5[7] ,n555);
    nand g1219(n1657 ,n39[0] ,n1480);
    nand g1220(n2101 ,n1828 ,n1659);
    nand g1221(n351 ,n12[3] ,n255);
    nor g1222(n1200 ,n38[0] ,n891);
    nand g1223(n761 ,n5[3] ,n561);
    nand g1224(n1279 ,n1078 ,n806);
    dff g1225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1163), .Q(n50[1]));
    nor g1226(n2123 ,n701 ,n1950);
    nand g1227(n2139 ,n1526 ,n2107);
    not g1228(n154 ,n153);
    dff g1229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2114), .Q(n38[2]));
    nand g1230(n520 ,n21[6] ,n430);
    nand g1231(n548 ,n23[2] ,n429);
    nor g1232(n2171 ,n598 ,n2160);
    nand g1233(n500 ,n21[1] ,n430);
    not g1234(n240 ,n20[0]);
    nand g1235(n1712 ,n39[0] ,n1467);
    nand g1236(n684 ,n27[3] ,n424);
    xnor g1237(n2189 ,n60[3] ,n130);
    dff g1238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2027), .Q(n36[0]));
    nand g1239(n2011 ,n1816 ,n1622);
    or g1240(n86 ,n58[4] ,n58[1]);
    nor g1241(n411 ,n58[4] ,n408);
    nand g1242(n1687 ,n39[4] ,n1487);
    nand g1243(n1628 ,n39[5] ,n1494);
    dff g1244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1332), .Q(n58[4]));
    xnor g1245(n2188 ,n60[2] ,n128);
    nor g1246(n1367 ,n299 ,n1198);
    nand g1247(n402 ,n37[2] ,n334);
    buf g1248(n15[1], 1'b0);
    nor g1249(n423 ,n270 ,n401);
    nand g1250(n1830 ,n1502 ,n1451);
    nor g1251(n888 ,n193 ,n590);
    nand g1252(n1626 ,n39[7] ,n1494);
    nor g1253(n2115 ,n695 ,n1951);
    nand g1254(n2084 ,n1765 ,n1700);
    nand g1255(n1327 ,n386 ,n1133);
    nand g1256(n1274 ,n397 ,n877);
    dff g1257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1147), .Q(n52[1]));
    dff g1258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1399), .Q(n11));
    nand g1259(n177 ,n20[7] ,n176);
    nand g1260(n1004 ,n465 ,n638);
    dff g1261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1750), .Q(n18[1]));
    not g1262(n229 ,n37[2]);
    nand g1263(n1137 ,n1035 ,n704);
    nand g1264(n572 ,n269 ,n440);
    not g1265(n421 ,n420);
    not g1266(n206 ,n2);
    nand g1267(n840 ,n59[2] ,n592);
    not g1268(n600 ,n540);
    dff g1269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2023), .Q(n36[4]));
    dff g1270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1980), .Q(n26[3]));
    dff g1271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2077), .Q(n30[3]));
    nand g1272(n1652 ,n39[1] ,n1484);
    nand g1273(n1774 ,n28[5] ,n1468);
    nand g1274(n1263 ,n19[1] ,n886);
    dff g1275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2056), .Q(n32[3]));
    nand g1276(n1811 ,n23[1] ,n1481);
    nand g1277(n1334 ,n1257 ,n1201);
    nand g1278(n944 ,n692 ,n612);
    nand g1279(n1661 ,n39[0] ,n1484);
    nand g1280(n353 ,n17[1] ,n309);
    not g1281(n341 ,n340);
    nand g1282(n187 ,n38[1] ,n38[0]);
    nand g1283(n1133 ,n2189 ,n893);
    dff g1284(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1234), .Q(n42[2]));
    nand g1285(n1076 ,n57[1] ,n553);
    nand g1286(n796 ,n5[3] ,n581);
    nand g1287(n748 ,n5[4] ,n577);
    nand g1288(n891 ,n194 ,n590);
    not g1289(n447 ,n446);
    nand g1290(n1411 ,n355 ,n1355);
    nor g1291(n580 ,n300 ,n437);
    nand g1292(n862 ,n10 ,n594);
    nor g1293(n388 ,n206 ,n327);
    dff g1294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1158), .Q(n50[6]));
    nand g1295(n1679 ,n39[7] ,n1493);
    dff g1296(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1395), .Q(n19[0]));
    dff g1297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2122), .Q(n38[3]));
    nor g1298(n2166 ,n599 ,n2159);
    dff g1299(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1184), .Q(n47[5]));
    not g1300(n234 ,n40[0]);
    nand g1301(n1003 ,n471 ,n636);
    not g1302(n2235 ,n2182);
    nand g1303(n2036 ,n1852 ,n1633);
    nand g1304(n1777 ,n2212 ,n1498);
    nand g1305(n1741 ,n36[6] ,n1466);
    nand g1306(n1763 ,n31[0] ,n1490);
    nand g1307(n1184 ,n933 ,n733);
    not g1308(n601 ,n541);
    nand g1309(n764 ,n5[0] ,n561);
    nor g1310(n110 ,n20[6] ,n109);
    nand g1311(n455 ,n2244 ,n381);
    nand g1312(n1055 ,n55[5] ,n558);
    nand g1313(n1310 ,n842 ,n496);
    nor g1314(n485 ,n192 ,n449);
    nand g1315(n1446 ,n53[2] ,n1375);
    dff g1316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1298), .Q(n55[1]));
    nand g1317(n858 ,n48[0] ,n563);
    nand g1318(n2126 ,n535 ,n2123);
    nand g1319(n851 ,n49[1] ,n579);
    nand g1320(n1217 ,n966 ,n756);
    nand g1321(n1906 ,n30[5] ,n1485);
    nand g1322(n2067 ,n881 ,n1902);
    dff g1323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1155), .Q(n51[1]));
    or g1324(n1103 ,n448 ,n1080);
    not g1325(n696 ,n647);
    dff g1326(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1330), .Q(n58[2]));
    nand g1327(n980 ,n42[4] ,n584);
    or g1328(n2144 ,n1864 ,n2137);
    nand g1329(n1148 ,n908 ,n716);
    nand g1330(n1976 ,n1781 ,n1590);
    nand g1331(n98 ,n93 ,n97);
    not g1332(n239 ,n8);
    nor g1333(n486 ,n193 ,n472);
    not g1334(n65 ,n64);
    nand g1335(n462 ,n40[7] ,n378);
    nor g1336(n1384 ,n38[3] ,n1201);
    nand g1337(n525 ,n22[4] ,n423);
    dff g1338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2080), .Q(n30[0]));
    nand g1339(n1275 ,n399 ,n861);
    dff g1340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1218), .Q(n44[1]));
    not g1341(n265 ,n266);
    nand g1342(n1013 ,n650 ,n648);
    nand g1343(n645 ,n2221 ,n421);
    not g1344(n142 ,n40[2]);
    nand g1345(n2100 ,n2196 ,n1755);
    dff g1346(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1507), .Q(n9));
    nand g1347(n1750 ,n1336 ,n1534);
    nand g1348(n704 ,n5[4] ,n559);
    nand g1349(n1955 ,n1115 ,n1586);
    nor g1350(n481 ,n245 ,n367);
    nand g1351(n518 ,n30[7] ,n425);
    or g1352(n1946 ,n1883 ,n1882);
    nand g1353(n678 ,n27[5] ,n424);
    nand g1354(n1168 ,n878 ,n811);
    not g1355(n1755 ,n891);
    nand g1356(n2124 ,n530 ,n2113);
    nand g1357(n772 ,n5[2] ,n573);
    nand g1358(n1010 ,n521 ,n520);
    nand g1359(n1854 ,n1436 ,n1420);
    nand g1360(n2001 ,n1806 ,n1613);
    nand g1361(n992 ,n515 ,n511);
    or g1362(n2147 ,n1851 ,n2138);
    nand g1363(n632 ,n2220 ,n421);
    nand g1364(n859 ,n20[0] ,n585);
    nand g1365(n1637 ,n39[3] ,n1472);
    nand g1366(n738 ,n5[7] ,n567);
    buf g1367(n418 ,n2186);
    nand g1368(n817 ,n5[6] ,n564);
    nand g1369(n1054 ,n56[0] ,n575);
    nand g1370(n1697 ,n39[6] ,n1493);
    nand g1371(n1331 ,n1048 ,n1316);
    nand g1372(n1952 ,n1097 ,n1581);
    nand g1373(n1732 ,n27[0] ,n1482);
    nand g1374(n591 ,n194 ,n478);
    nor g1375(n476 ,n268 ,n403);
    nor g1376(n438 ,n60[3] ,n400);
    nand g1377(n1973 ,n1730 ,n1677);
    nand g1378(n1766 ,n29[5] ,n1470);
    nand g1379(n544 ,n31[1] ,n427);
    nand g1380(n2091 ,n1770 ,n1705);
    dff g1381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2059), .Q(n32[0]));
    dff g1382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n294), .Q(n13[6]));
    nand g1383(n463 ,n40[5] ,n378);
    nand g1384(n1850 ,n1577 ,n1430);
    nand g1385(n1778 ,n2200 ,n1498);
    nand g1386(n1330 ,n1031 ,n1317);
    nand g1387(n876 ,n56[4] ,n575);
    nand g1388(n977 ,n42[7] ,n584);
    nand g1389(n1537 ,n49[3] ,n1369);
    nand g1390(n732 ,n5[6] ,n565);
    nand g1391(n1205 ,n951 ,n747);
    nand g1392(n405 ,n249 ,n315);
    nand g1393(n656 ,n28[6] ,n432);
    nor g1394(n2108 ,n1936 ,n1935);
    dff g1395(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1248), .Q(n40[7]));
    not g1396(n695 ,n617);
    nor g1397(n85 ,n58[3] ,n83);
    nand g1398(n2039 ,n1862 ,n1636);
    nand g1399(n267 ,n59[1] ,n227);
    nand g1400(n501 ,n23[5] ,n429);
    not g1401(n209 ,n18[0]);
    nor g1402(n413 ,n17[1] ,n406);
    nor g1403(n1467 ,n298 ,n1381);
    nand g1404(n1177 ,n854 ,n819);
    nand g1405(n1280 ,n883 ,n802);
    nand g1406(n556 ,n269 ,n442);
    dff g1407(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1325), .Q(n41[2]));
    nand g1408(n1321 ,n384 ,n1135);
    nand g1409(n190 ,n19[3] ,n19[2]);
    nand g1410(n1029 ,n672 ,n669);
    nand g1411(n912 ,n51[5] ,n570);
    dff g1412(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1253), .Q(n40[2]));
    nand g1413(n1591 ,n39[6] ,n1474);
    not g1414(n257 ,n256);
    dff g1415(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1334), .Q(n38[0]));
    nand g1416(n1764 ,n29[7] ,n1470);
    dff g1417(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1168), .Q(n49[4]));
    nand g1418(n2059 ,n1899 ,n1660);
    dff g1419(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2032), .Q(n35[3]));
    nand g1420(n1896 ,n32[2] ,n1489);
    nand g1421(n148 ,n40[4] ,n147);
    nor g1422(n90 ,n19[2] ,n19[0]);
    nand g1423(n1756 ,n31[5] ,n1490);
    nand g1424(n657 ,n33[6] ,n434);
    nand g1425(n1991 ,n1796 ,n1655);
    nand g1426(n504 ,n26[2] ,n431);
    dff g1427(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2037), .Q(n34[6]));
    nor g1428(n264 ,n225 ,n60[1]);
    nand g1429(n1465 ,n350 ,n1352);
    nand g1430(n1497 ,n266 ,n1379);
    nor g1431(n2107 ,n1933 ,n1932);
    nand g1432(n2092 ,n1771 ,n1718);
    dff g1433(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1587), .Q(n18[0]));
    dff g1434(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2174), .Q(n61[5]));
    nand g1435(n2053 ,n1889 ,n1640);
    not g1436(n236 ,n40[4]);
    nand g1437(n1046 ,n604 ,n674);
    xor g1438(n2215 ,n40[1] ,n40[0]);
    nor g1439(n361 ,n219 ,n328);
    dff g1440(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2084), .Q(n29[6]));
    nand g1441(n1847 ,n1530 ,n1438);
    nand g1442(n1790 ,n25[6] ,n1477);
    nand g1443(n1407 ,n46[3] ,n1374);
    nand g1444(n392 ,n308 ,n312);
    nand g1445(n1877 ,n1563 ,n1447);
    nand g1446(n1724 ,n28[0] ,n1468);
    nand g1447(n1747 ,n35[1] ,n1492);
    nand g1448(n1322 ,n1131 ,n1263);
    xnor g1449(n2191 ,n59[2] ,n138);
    dff g1450(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n385), .Q(n37[0]));
    nand g1451(n952 ,n693 ,n646);
    nand g1452(n1970 ,n843 ,n1778);
    not g1453(n383 ,n382);
    nand g1454(n837 ,n20[9] ,n585);
    nand g1455(n785 ,n5[6] ,n559);
    nor g1456(n1370 ,n261 ,n1197);
    nand g1457(n926 ,n50[0] ,n574);
    nor g1458(n291 ,n243 ,n193);
    nand g1459(n1512 ,n1339 ,n1360);
    nand g1460(n298 ,n38[1] ,n38[2]);
    nand g1461(n682 ,n2223 ,n421);
    nor g1462(n2106 ,n1930 ,n1929);
    nor g1463(n1347 ,n199 ,n1310);
    dff g1464(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1754), .Q(n62[2]));
    not g1465(n228 ,n38[2]);
    dff g1466(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1966), .Q(n20[1]));
    nand g1467(n1739 ,n36[0] ,n1466);
    nand g1468(n2060 ,n1919 ,n1690);
    nand g1469(n1845 ,n1527 ,n1233);
    dff g1470(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2130), .Q(n12[5]));
    not g1471(n1390 ,n1322);
    or g1472(n1102 ,n938 ,n931);
    nand g1473(n1836 ,n2192 ,n1499);
    not g1474(n589 ,n588);
    dff g1475(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1304), .Q(n54[3]));
    or g1476(n1108 ,n1042 ,n1032);
    nand g1477(n1880 ,n1546 ,n1568);
    nand g1478(n1987 ,n1791 ,n1601);
    nand g1479(n1769 ,n29[2] ,n1470);
    nand g1480(n1851 ,n1421 ,n1435);
    nand g1481(n261 ,n59[2] ,n226);
    dff g1482(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n288), .Q(n16[9]));
    or g1483(n1932 ,n1901 ,n1841);
    nand g1484(n1781 ,n26[7] ,n1475);
    xor g1485(n2208 ,n18[1] ,n18[0]);
    nand g1486(n1417 ,n50[6] ,n1364);
    nand g1487(n854 ,n48[4] ,n563);
    nand g1488(n765 ,n5[7] ,n583);
    nand g1489(n648 ,n33[0] ,n434);
    nand g1490(n749 ,n5[2] ,n577);
    dff g1491(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1277), .Q(n57[7]));
    nand g1492(n1402 ,n352 ,n1356);
    nand g1493(n1799 ,n24[5] ,n1479);
    nand g1494(n981 ,n55[3] ,n558);
    nor g1495(n1355 ,n1093 ,n1102);
    nand g1496(n2064 ,n1756 ,n1693);
    nand g1497(n1180 ,n857 ,n822);
    not g1498(n193 ,n194);
    not g1499(n561 ,n562);
    nand g1500(n958 ,n616 ,n498);
    dff g1501(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n452), .Q(n13[3]));
    nand g1502(n1534 ,n2208 ,n1385);
    nand g1503(n355 ,n12[1] ,n255);
    nand g1504(n1695 ,n39[3] ,n1491);
    nand g1505(n1006 ,n639 ,n690);
    nand g1506(n1078 ,n57[3] ,n553);
    nor g1507(n104 ,n20[11] ,n20[10]);
    nand g1508(n1547 ,n56[1] ,n1377);
    nand g1509(n1734 ,n36[7] ,n1466);
    nand g1510(n2132 ,n1521 ,n2105);
    nand g1511(n2057 ,n1896 ,n1644);
    nand g1512(n1514 ,n49[7] ,n1369);
    not g1513(n224 ,n37[0]);
    not g1514(n163 ,n20[4]);
    nand g1515(n1958 ,n859 ,n1662);
    dff g1516(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1157), .Q(n50[7]));
    nor g1517(n433 ,n268 ,n380);
    nand g1518(n1305 ,n1064 ,n797);
    nand g1519(n496 ,n417 ,n467);
    nand g1520(n1533 ,n57[4] ,n1362);
    dff g1521(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1300), .Q(n54[7]));
    nand g1522(n1434 ,n51[2] ,n1365);
    nand g1523(n1874 ,n1418 ,n1445);
    nand g1524(n390 ,n2244 ,n337);
    nand g1525(n830 ,n5[3] ,n576);
    nand g1526(n1432 ,n46[4] ,n1374);
    not g1527(n1466 ,n1467);
    dff g1528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1220), .Q(n43[7]));
    nand g1529(n408 ,n251 ,n321);
    nor g1530(n1392 ,n18[0] ,n1386);
    dff g1531(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1215), .Q(n44[4]));
    nand g1532(n723 ,n5[1] ,n569);
    nand g1533(n1231 ,n980 ,n769);
    nand g1534(n1735 ,n36[5] ,n1466);
    nor g1535(n1101 ,n1021 ,n1020);
    nand g1536(n844 ,n20[1] ,n585);
    nor g1537(n1583 ,n1006 ,n1415);
    nand g1538(n503 ,n22[0] ,n423);
    nand g1539(n1558 ,n48[5] ,n1367);
    dff g1540(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1977), .Q(n26[6]));
    dff g1541(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1255), .Q(n46[2]));
    nor g1542(n1585 ,n1018 ,n1465);
    nor g1543(n340 ,n37[3] ,n301);
    dff g1544(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1302), .Q(n54[5]));
    nand g1545(n814 ,n5[1] ,n580);
    not g1546(n227 ,n59[2]);
    not g1547(n207 ,n19[4]);
    dff g1548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2025), .Q(n36[2]));
    dff g1549(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1508), .Q(n19[4]));
    nand g1550(n692 ,n26[1] ,n431);
    nand g1551(n2129 ,n538 ,n2117);
    not g1552(n339 ,n338);
    nand g1553(n1298 ,n960 ,n774);
    nand g1554(n1051 ,n545 ,n527);
    nand g1555(n96 ,n40[9] ,n40[8]);
    dff g1556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n295), .Q(n13[7]));
    dff g1557(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1138), .Q(n46[4]));
    nand g1558(n1618 ,n39[1] ,n1480);
    nand g1559(n1908 ,n30[3] ,n1485);
    nor g1560(n1581 ,n1005 ,n1416);
    nand g1561(n1713 ,n39[0] ,n1469);
    nand g1562(n1445 ,n54[2] ,n1373);
    or g1563(n1196 ,n59[0] ,n1079);
    dff g1564(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1509), .Q(n19[3]));
    nand g1565(n1806 ,n23[6] ,n1481);
    nand g1566(n1199 ,n59[0] ,n895);
    nor g1567(n294 ,n212 ,n192);
    nand g1568(n1553 ,n48[0] ,n1367);
    dff g1569(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1238), .Q(n51[2]));
    dff g1570(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1214), .Q(n44[5]));
    dff g1571(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1185), .Q(n47[4]));
    nand g1572(n727 ,n5[3] ,n573);
    nor g1573(n2119 ,n700 ,n1955);
    nor g1574(n426 ,n270 ,n402);
    not g1575(n92 ,n40[5]);
    dff g1576(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1148), .Q(n52[0]));
    nand g1577(n616 ,n28[5] ,n432);
    nand g1578(n1664 ,n39[6] ,n1467);
    nand g1579(n1007 ,n642 ,n516);
    not g1580(n220 ,n39[0]);
    nand g1581(n2225 ,n81 ,n80);
    dff g1582(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1226), .Q(n43[1]));
    nand g1583(n2076 ,n1907 ,n1649);
    nand g1584(n2086 ,n1767 ,n1702);
    nand g1585(n498 ,n31[5] ,n427);
    nor g1586(n2140 ,n1833 ,n2132);
    nand g1587(n1413 ,n51[4] ,n1365);
    nand g1588(n1505 ,n43[3] ,n1363);
    nor g1589(n1369 ,n299 ,n1199);
    nand g1590(n1479 ,n272 ,n1379);
    not g1591(n1490 ,n1491);
    nand g1592(n1283 ,n61[1] ,n887);
    nand g1593(n873 ,n20[4] ,n585);
    nand g1594(n628 ,n2224 ,n421);
    nor g1595(n1358 ,n254 ,n1194);
    not g1596(n565 ,n566);
    nand g1597(n1726 ,n27[6] ,n1482);
    nor g1598(n186 ,n38[1] ,n38[0]);
    nand g1599(n72 ,n68 ,n70);
    or g1600(n1939 ,n1861 ,n1860);
    or g1601(n1096 ,n1001 ,n999);
    buf g1602(n14[3], 1'b0);
    nor g1603(n482 ,n192 ,n454);
    nand g1604(n1502 ,n43[7] ,n1363);
    nand g1605(n919 ,n50[6] ,n574);
    nand g1606(n1067 ,n52[5] ,n572);
    nand g1607(n443 ,n17[2] ,n369);
    nor g1608(n101 ,n40[7] ,n100);
    nand g1609(n770 ,n5[3] ,n583);
    nand g1610(n1140 ,n900 ,n708);
    dff g1611(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2052), .Q(n32[7]));
    nand g1612(n1174 ,n853 ,n817);
    nand g1613(n1138 ,n943 ,n741);
    buf g1614(n14[0], 1'b0);
    nand g1615(n1951 ,n1091 ,n1580);
    nand g1616(n1665 ,n39[5] ,n1467);
    nand g1617(n311 ,n199 ,n277);
    nand g1618(n2099 ,n2197 ,n1755);
    nand g1619(n1808 ,n23[4] ,n1481);
    nand g1620(n461 ,n40[8] ,n378);
    xor g1621(n2238 ,n77 ,n19[3]);
    nand g1622(n166 ,n20[1] ,n20[0]);
    not g1623(n593 ,n301);
    nor g1624(n458 ,n363 ,n365);
    nand g1625(n588 ,n331 ,n478);
    nand g1626(n2085 ,n1766 ,n1701);
    nand g1627(n815 ,n5[0] ,n580);
    nand g1628(n535 ,n30[2] ,n425);
    nand g1629(n1655 ,n39[0] ,n1476);
    nand g1630(n1021 ,n658 ,n657);
    nand g1631(n1673 ,n39[6] ,n1483);
    dff g1632(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n494), .Q(n39[7]));
    nand g1633(n2024 ,n1737 ,n1667);
    nand g1634(n409 ,n60[3] ,n330);
    not g1635(n1388 ,n1319);
    nand g1636(n716 ,n5[0] ,n571);
    dff g1637(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n482), .Q(n39[2]));
    nand g1638(n465 ,n40[1] ,n378);
    nand g1639(n1017 ,n2194 ,n593);
    nand g1640(n1028 ,n677 ,n673);
    nand g1641(n1596 ,n39[1] ,n1474);
    nand g1642(n1792 ,n25[5] ,n1477);
    not g1643(n1084 ,n996);
    dff g1644(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2031), .Q(n35[4]));
    dff g1645(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1113), .Q(n59[0]));
    nand g1646(n969 ,n43[7] ,n562);
    nand g1647(n1161 ,n921 ,n727);
    nand g1648(n1760 ,n31[3] ,n1490);
    nand g1649(n1426 ,n54[6] ,n1373);
    nor g1650(n365 ,n218 ,n327);
    nand g1651(n1501 ,n48[2] ,n1367);
    dff g1652(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1988), .Q(n25[3]));
    nand g1653(n1134 ,n2188 ,n893);
    nand g1654(n69 ,n2207 ,n66);
    nand g1655(n1684 ,n39[6] ,n1487);
    nand g1656(n460 ,n40[3] ,n378);
    nand g1657(n878 ,n49[4] ,n579);
    not g1658(n603 ,n551);
    not g1659(n1082 ,n991);
    nand g1660(n1264 ,n61[4] ,n887);
    dff g1661(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1289), .Q(n56[3]));
    nand g1662(n2133 ,n1520 ,n2106);
    nand g1663(n471 ,n40[2] ,n378);
    dff g1664(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1206), .Q(n45[5]));
    nand g1665(n134 ,n58[2] ,n133);
    not g1666(n274 ,n273);
    nand g1667(n1456 ,n50[0] ,n1364);
    nand g1668(n638 ,n2215 ,n421);
    nand g1669(n667 ,n24[4] ,n428);
    nand g1670(n1506 ,n56[3] ,n1377);
    nand g1671(n84 ,n58[2] ,n80);
    nand g1672(n1169 ,n849 ,n812);
    not g1673(n575 ,n576);
    nand g1674(n387 ,n2235 ,n338);
    nor g1675(n1491 ,n271 ,n1380);
    nor g1676(n1366 ,n267 ,n1198);
    nand g1677(n1809 ,n23[3] ,n1481);
    nand g1678(n942 ,n46[5] ,n568);
    nor g1679(n144 ,n142 ,n143);
    nand g1680(n1188 ,n1043 ,n736);
    nor g1681(n1373 ,n261 ,n1196);
    not g1682(n243 ,n40[10]);
    nand g1683(n1295 ,n981 ,n792);
    nand g1684(n1531 ,n46[1] ,n1374);
    nand g1685(n635 ,n2218 ,n421);
    dff g1686(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1165), .Q(n49[7]));
    nor g1687(n1362 ,n299 ,n1197);
    dff g1688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1964), .Q(n28[0]));
    dff g1689(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1324), .Q(n41[1]));
    nand g1690(n1975 ,n1732 ,n1714);
    nand g1691(n2046 ,n1753 ,n1685);
    dff g1692(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2095), .Q(n28[5]));
    nand g1693(n650 ,n32[0] ,n436);
    nand g1694(n1607 ,n39[5] ,n1478);
    nand g1695(n966 ,n44[2] ,n556);
    nand g1696(n1540 ,n43[2] ,n1363);
    nand g1697(n1983 ,n1788 ,n1654);
    nand g1698(n470 ,n40[9] ,n378);
    nand g1699(n624 ,n34[2] ,n426);
    nand g1700(n822 ,n5[1] ,n564);
    nor g1701(n1928 ,n1856 ,n1834);
    nand g1702(n2173 ,n1533 ,n2165);
    nand g1703(n1037 ,n50[7] ,n574);
    nand g1704(n140 ,n59[2] ,n139);
    nor g1705(n371 ,n197 ,n327);
    nand g1706(n754 ,n5[4] ,n555);
    not g1707(n329 ,n330);
    nand g1708(n2015 ,n1820 ,n1658);
    nand g1709(n647 ,n36[7] ,n422);
    nand g1710(n1615 ,n39[4] ,n1480);
    nor g1711(n576 ,n300 ,n439);
    not g1712(n2185 ,n17[2]);
    dff g1713(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2079), .Q(n30[1]));
    nand g1714(n677 ,n26[5] ,n431);
    nor g1715(n585 ,n192 ,n481);
    nand g1716(n1839 ,n1566 ,n1426);
    nand g1717(n473 ,n2244 ,n392);
    dff g1718(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1288), .Q(n56[4]));
    nor g1719(n1582 ,n192 ,n1394);
    nand g1720(n1193 ,n1026 ,n706);
    nand g1721(n529 ,n23[1] ,n429);
    nand g1722(n615 ,n28[1] ,n432);
    nand g1723(n1800 ,n24[4] ,n1479);
    buf g1724(n14[7], 1'b0);
    nand g1725(n2163 ,n1450 ,n2154);
    nand g1726(n541 ,n61[7] ,n475);
    nor g1727(n431 ,n270 ,n403);
    nand g1728(n1189 ,n1040 ,n737);
    dff g1729(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2026), .Q(n36[1]));
    dff g1730(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1990), .Q(n25[1]));
    nand g1731(n1980 ,n1785 ,n1594);
    dff g1732(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n284), .Q(n16[0]));
    nand g1733(n2027 ,n1739 ,n1712);
    nor g1734(n864 ,n466 ,n489);
    nand g1735(n1803 ,n24[1] ,n1479);
    nand g1736(n686 ,n33[5] ,n434);
    nand g1737(n1401 ,n50[2] ,n1364);
    nor g1738(n2150 ,n1934 ,n2142);
    nor g1739(n1117 ,n925 ,n928);
    nor g1740(n315 ,n193 ,n250);
    not g1741(n479 ,n480);
    nand g1742(n872 ,n48[5] ,n563);
    nand g1743(n644 ,n32[7] ,n436);
    nand g1744(n706 ,n5[3] ,n559);
    nand g1745(n2134 ,n1542 ,n2110);
    nor g1746(n1365 ,n262 ,n1197);
    nor g1747(n1126 ,n192 ,n864);
    nand g1748(n1012 ,n694 ,n619);
    nand g1749(n2164 ,n1425 ,n2161);
    nand g1750(n756 ,n5[2] ,n555);
    nand g1751(n1163 ,n924 ,n728);
    dff g1752(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1748), .Q(n18[2]));
    nand g1753(n1619 ,n39[7] ,n1496);
    or g1754(n247 ,n193 ,n2241);
    nor g1755(n1487 ,n259 ,n1380);
    nand g1756(n2159 ,n1431 ,n2150);
    nor g1757(n596 ,n333 ,n445);
    dff g1758(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1303), .Q(n54[4]));
    nand g1759(n2049 ,n1922 ,n1688);
    nand g1760(n967 ,n44[1] ,n556);
    dff g1761(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1959), .Q(n59[2]));
    nand g1762(n1677 ,n39[2] ,n1483);
    dff g1763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1181), .Q(n48[0]));
    nand g1764(n1639 ,n39[7] ,n1488);
    nor g1765(n359 ,n277 ,n335);
    nand g1766(n659 ,n36[6] ,n422);
    nand g1767(n805 ,n5[5] ,n554);
    nand g1768(n1706 ,n39[7] ,n1469);
    nand g1769(n1733 ,n36[2] ,n1466);
    nor g1770(n151 ,n141 ,n150);
    nand g1771(n619 ,n25[6] ,n476);
    nand g1772(n119 ,n20[9] ,n20[8]);
    nand g1773(n354 ,n12[7] ,n255);
    nand g1774(n1187 ,n937 ,n789);
    nand g1775(n1804 ,n24[0] ,n1479);
    nand g1776(n160 ,n37[1] ,n37[0]);
    nor g1777(n1350 ,n1107 ,n1106);
    nor g1778(n263 ,n60[1] ,n60[2]);
    dff g1779(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2038), .Q(n34[5]));
    nor g1780(n360 ,n197 ,n328);
    nand g1781(n2068 ,n1761 ,n1696);
    nand g1782(n774 ,n5[1] ,n557);
    nand g1783(n903 ,n52[4] ,n572);
    nand g1784(n352 ,n12[2] ,n255);
    nand g1785(n843 ,n20[3] ,n585);
    nand g1786(n1703 ,n39[3] ,n1471);
    nand g1787(n1972 ,n1729 ,n1676);
    nand g1788(n758 ,n5[7] ,n561);
    nand g1789(n679 ,n34[5] ,n426);
    nand g1790(n1186 ,n935 ,n735);
    nand g1791(n2083 ,n869 ,n1913);
    dff g1792(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2164), .Q(n61[7]));
    nand g1793(n1226 ,n975 ,n763);
    or g1794(n75 ,n67 ,n73);
    nor g1795(n587 ,n193 ,n478);
    nor g1796(n2165 ,n602 ,n2158);
    not g1797(n198 ,n39[4]);
    dff g1798(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1245), .Q(n40[10]));
    nand g1799(n1604 ,n39[1] ,n1476);
    nand g1800(n1740 ,n35[7] ,n1492);
    nand g1801(n794 ,n5[6] ,n581);
    nand g1802(n1736 ,n36[4] ,n1466);
    dff g1803(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2019), .Q(n21[4]));
    not g1804(n598 ,n517);
    nand g1805(n2070 ,n1763 ,n1717);
    nand g1806(n787 ,n5[0] ,n577);
    nand g1807(n1158 ,n919 ,n784);
    dff g1808(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1276), .Q(n58[0]));
    not g1809(n1309 ,n1310);
    nand g1810(n1649 ,n39[4] ,n1484);
    or g1811(n1106 ,n929 ,n930);
    dff g1812(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2018), .Q(n21[5]));
    nand g1813(n1636 ,n39[4] ,n1472);
    or g1814(n1104 ,n1038 ,n1030);
    nand g1815(n1131 ,n2240 ,n885);
    nand g1816(n719 ,n5[5] ,n569);
    dff g1817(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2086), .Q(n29[4]));
    nor g1818(n333 ,n62[2] ,n257);
    nand g1819(n1431 ,n51[5] ,n1365);
    nand g1820(n1560 ,n43[5] ,n1363);
    not g1821(n1315 ,n1273);
    nand g1822(n1552 ,n47[0] ,n1371);
    nor g1823(n1376 ,n262 ,n1198);
    xnor g1824(n2219 ,n40[5] ,n148);
    nand g1825(n1700 ,n39[6] ,n1471);
    nand g1826(n1171 ,n851 ,n814);
    nand g1827(n1609 ,n39[3] ,n1478);
    dff g1828(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2066), .Q(n31[3]));
    nor g1829(n1249 ,n192 ,n1085);
    nor g1830(n1308 ,n192 ,n1090);
    nand g1831(n2054 ,n1890 ,n1641);
    nand g1832(n640 ,n35[7] ,n435);
    dff g1833(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1328), .Q(n60[2]));
    nand g1834(n939 ,n660 ,n686);
    nor g1835(n338 ,n221 ,n302);
    dff g1836(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1145), .Q(n52[3]));
    nand g1837(n1717 ,n39[0] ,n1491);
    dff g1838(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2028), .Q(n35[7]));
    dff g1839(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2040), .Q(n34[3]));
    dff g1840(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n296), .Q(n15[6]));
    nand g1841(n1524 ,n45[5] ,n1372);
    nand g1842(n1408 ,n50[7] ,n1364);
    nor g1843(n286 ,n242 ,n193);
    not g1844(n1378 ,n1379);
    nand g1845(n1019 ,n2193 ,n593);
    nand g1846(n509 ,n23[0] ,n429);
    nand g1847(n1688 ,n39[2] ,n1487);
    dff g1848(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n289), .Q(n16[8]));
    nand g1849(n1195 ,n838 ,n594);
    nor g1850(n100 ,n92 ,n99);
    dff g1851(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2017), .Q(n21[6]));
    nand g1852(n2037 ,n1855 ,n1634);
    dff g1853(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n283), .Q(n16[4]));
    nand g1854(n1015 ,n618 ,n665);
    nand g1855(n1824 ,n21[4] ,n1495);
    nor g1856(n1343 ,n344 ,n1309);
    not g1857(n571 ,n572);
    nand g1858(n1601 ,n39[4] ,n1476);
    nand g1859(n1202 ,n38[0] ,n892);
    nor g1860(n494 ,n192 ,n457);
    nand g1861(n957 ,n45[1] ,n578);
    nand g1862(n1527 ,n49[5] ,n1369);
    nand g1863(n947 ,n46[1] ,n568);
    dff g1864(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1996), .Q(n24[3]));
    or g1865(n1197 ,n200 ,n1079);
    nand g1866(n1296 ,n1057 ,n793);
    nor g1867(n1498 ,n192 ,n1338);
    nand g1868(n1052 ,n53[1] ,n560);
    dff g1869(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1278), .Q(n57[5]));
    nand g1870(n1849 ,n1522 ,n1432);
    nand g1871(n1255 ,n946 ,n742);
    nand g1872(n1691 ,n39[5] ,n1493);
    nand g1873(n1276 ,n867 ,n833);
    nor g1874(n372 ,n196 ,n327);
    nand g1875(n1500 ,n45[2] ,n1372);
    dff g1876(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n414), .Q(n13[4]));
    or g1877(n1094 ,n995 ,n992);
    nor g1878(n449 ,n366 ,n374);
    nand g1879(n1671 ,n39[1] ,n1469);
    dff g1880(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1962), .Q(n28[1]));
    nand g1881(n1419 ,n50[5] ,n1364);
    nor g1882(n1375 ,n267 ,n1197);
    not g1883(n237 ,n40[2]);
    nand g1884(n246 ,n17[0] ,n206);
    not g1885(n211 ,n9);
    nand g1886(n849 ,n49[3] ,n579);
    nand g1887(n1742 ,n35[6] ,n1492);
    nand g1888(n1267 ,n1054 ,n832);
    dff g1889(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1983), .Q(n26[0]));
    xnor g1890(n2209 ,n185 ,n18[2]);
    dff g1891(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2126), .Q(n12[2]));
    nand g1892(n1405 ,n53[3] ,n1375);
    nand g1893(n1287 ,n1073 ,n828);
    nand g1894(n2174 ,n1557 ,n2166);
    nand g1895(n300 ,n60[1] ,n60[2]);
    nand g1896(n707 ,n5[1] ,n559);
    nand g1897(n1318 ,n1128 ,n1121);
    dff g1898(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n411), .Q(n13[5]));
    nand g1899(n517 ,n61[3] ,n475);
    nor g1900(n2113 ,n699 ,n1957);
    dff g1901(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1292), .Q(n55[7]));
    nor g1902(n284 ,n234 ,n193);
    nand g1903(n2050 ,n1921 ,n1689);
    nand g1904(n1862 ,n34[4] ,n1473);
    dff g1905(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2057), .Q(n32[2]));
    nand g1906(n1956 ,n1122 ,n1588);
    nand g1907(n773 ,n5[0] ,n583);
    nand g1908(n1674 ,n39[5] ,n1483);
    xor g1909(n2239 ,n72 ,n19[2]);
    nand g1910(n795 ,n5[4] ,n581);
    not g1911(n1090 ,n1004);
    nand g1912(n1606 ,n39[6] ,n1478);
    nand g1913(n737 ,n5[0] ,n565);
    nand g1914(n1795 ,n25[1] ,n1477);
    not g1915(n701 ,n687);
    nand g1916(n2088 ,n1768 ,n1703);
    nand g1917(n1440 ,n55[3] ,n1370);
    xnor g1918(n2213 ,n20[6] ,n173);
    nor g1919(n564 ,n300 ,n441);
    nor g1920(n1346 ,n223 ,n1310);
    nand g1921(n1737 ,n36[3] ,n1466);
    dff g1922(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1178), .Q(n48[3]));
    nand g1923(n2242 ,n90 ,n91);
    nand g1924(n909 ,n52[6] ,n572);
    nand g1925(n1708 ,n39[6] ,n1469);
    nand g1926(n511 ,n21[7] ,n430);
    nand g1927(n536 ,n30[4] ,n425);
    dff g1928(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2005), .Q(n23[2]));
    dff g1929(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1162), .Q(n50[2]));
    dff g1930(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n799), .Q(n6));
    nand g1931(n1914 ,n30[0] ,n1485);
    dff g1932(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1973), .Q(n27[2]));
    dff g1933(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1287), .Q(n56[5]));
    nand g1934(n1485 ,n266 ,n1382);
    or g1935(n268 ,n37[0] ,n37[1]);
    nand g1936(n1066 ,n54[1] ,n582);
    nand g1937(n931 ,n546 ,n500);
    nand g1938(n277 ,n17[2] ,n223);
    nand g1939(n1212 ,n961 ,n751);
    nand g1940(n73 ,n65 ,n69);
    nor g1941(n429 ,n258 ,n401);
    dff g1942(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1137), .Q(n53[4]));
    nand g1943(n2042 ,n1868 ,n1638);
    dff g1944(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1180), .Q(n48[1]));
    or g1945(n1929 ,n1924 ,n1835);
    nand g1946(n389 ,n60[2] ,n331);
    or g1947(n1123 ,n917 ,n914);
    dff g1948(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1173), .Q(n48[7]));
    nand g1949(n2162 ,n1463 ,n2153);
    nand g1950(n1969 ,n1727 ,n1674);
    nand g1951(n130 ,n60[2] ,n129);
    or g1952(n1198 ,n59[0] ,n896);
    nand g1953(n2236 ,n87 ,n88);
    nand g1954(n643 ,n33[7] ,n434);
    nand g1955(n1477 ,n260 ,n1384);
    nor g1956(n1372 ,n267 ,n1199);
    nand g1957(n1872 ,n1541 ,n1444);
    nor g1958(n1586 ,n1025 ,n1453);
    nor g1959(n1253 ,n193 ,n1089);
    nand g1960(n1884 ,n1551 ,n1464);
    nand g1961(n1179 ,n856 ,n825);
    nand g1962(n1008 ,n644 ,n643);
    nand g1963(n542 ,n31[4] ,n427);
    nand g1964(n1857 ,n1505 ,n1410);
    dff g1965(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1258), .Q(n37[3]));
    nand g1966(n1521 ,n56[7] ,n1377);
    not g1967(n702 ,n691);
    nand g1968(n788 ,n5[1] ,n555);
    nor g1969(n1250 ,n193 ,n1086);
    not g1970(n194 ,n2186);
    nand g1971(n2025 ,n1733 ,n1668);
    nand g1972(n1757 ,n2191 ,n1499);
    xor g1973(n2228 ,n58[4] ,n85);
    dff g1974(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1179), .Q(n48[2]));
    not g1975(n407 ,n406);
    nand g1976(n914 ,n504 ,n671);
    nand g1977(n1160 ,n920 ,n726);
    not g1978(n1386 ,n1385);
    dff g1979(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1986), .Q(n25[5]));
    nand g1980(n1868 ,n34[1] ,n1473);
    nand g1981(n1518 ,n45[6] ,n1372);
    nand g1982(n718 ,n5[6] ,n569);
    nand g1983(n2013 ,n1818 ,n1624);
    nor g1984(n1344 ,n232 ,n1195);
    nor g1985(n1097 ,n1008 ,n1007);
    nand g1986(n1448 ,n55[1] ,n1370);
    dff g1987(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1256), .Q(n55[4]));
    nand g1988(n1213 ,n962 ,n752);
    nand g1989(n1513 ,n48[7] ,n1367);
    nand g1990(n1011 ,n649 ,n522);
    not g1991(n698 ,n659);
    nand g1992(n691 ,n36[4] ,n422);
    nand g1993(n1185 ,n934 ,n734);
    nor g1994(n125 ,n119 ,n124);
    dff g1995(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1160), .Q(n50[4]));
    xnor g1996(n884 ,n478 ,n200);
    nand g1997(n1454 ,n52[5] ,n1368);
    nand g1998(n1651 ,n39[2] ,n1484);
    nand g1999(n1048 ,n2227 ,n587);
    nand g2000(n136 ,n58[3] ,n135);
    nand g2001(n2207 ,n2181 ,n2184);
    nand g2002(n1562 ,n56[4] ,n1377);
    nand g2003(n848 ,n49[5] ,n579);
    nand g2004(n1151 ,n912 ,n719);
    nand g2005(n254 ,n62[1] ,n222);
    nand g2006(n2003 ,n1808 ,n1615);
    nand g2007(n1996 ,n1801 ,n1609);
    dff g2008(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1993), .Q(n24[6]));
    nor g2009(n266 ,n38[1] ,n38[2]);
    nand g2010(n419 ,n391 ,n404);
    nand g2011(n1905 ,n30[6] ,n1485);
    nand g2012(n1812 ,n23[0] ,n1481);
    dff g2013(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1965), .Q(n20[4]));
    nand g2014(n1977 ,n1782 ,n1591);
    nand g2015(n1776 ,n28[3] ,n1468);
    nand g2016(n1236 ,n986 ,n773);
    nand g2017(n982 ,n42[3] ,n584);
    nand g2018(n883 ,n57[4] ,n553);
    xnor g2019(n2202 ,n20[7] ,n175);
    nand g2020(n1873 ,n1501 ,n1401);
    nand g2021(n2026 ,n1738 ,n1669);
    dff g2022(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1161), .Q(n50[3]));
    nand g2023(n1064 ,n54[2] ,n582);
    nand g2024(n1565 ,n44[1] ,n1366);
    or g2025(n1926 ,n1831 ,n1830);
    nor g2026(n1111 ,n17[2] ,n835);
    nand g2027(n775 ,n5[3] ,n577);
    nand g2028(n760 ,n5[5] ,n561);
    not g2029(n279 ,n278);
    nand g2030(n963 ,n44[5] ,n556);
    dff g2031(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1143), .Q(n52[5]));
    nand g2032(n2056 ,n1895 ,n1643);
    nand g2033(n1920 ,n33[0] ,n1486);
    not g2034(n83 ,n82);
    not g2035(n238 ,n40[6]);
    buf g2036(n16[14], 1'b0);
    nand g2037(n672 ,n26[3] ,n431);
    or g2038(n1942 ,n1873 ,n1872);
    nand g2039(n493 ,n415 ,n447);
    dff g2040(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2073), .Q(n30[6]));
    nand g2041(n1913 ,n2214 ,n1498);
    not g2042(n1313 ,n1237);
    not g2043(n241 ,n10);
    dff g2044(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1144), .Q(n52[4]));
    nor g2045(n366 ,n195 ,n328);
    nor g2046(n483 ,n192 ,n456);
    nand g2047(n1598 ,n39[2] ,n1472);
    dff g2048(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1280), .Q(n57[4]));
    nand g2049(n1953 ,n1100 ,n1583);
    nand g2050(n1749 ,n35[0] ,n1492);
    nand g2051(n1817 ,n22[3] ,n1497);
    nor g2052(n328 ,n302 ,n275);
    dff g2053(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2008), .Q(n22[6]));
    dff g2054(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1210), .Q(n45[1]));
    nand g2055(n1682 ,n39[2] ,n1493);
    nand g2056(n1225 ,n974 ,n762);
    xnor g2057(n2212 ,n20[4] ,n170);
    nand g2058(n934 ,n47[4] ,n566);
    nor g2059(n330 ,n192 ,n306);
    dff g2060(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2048), .Q(n33[3]));
    or g2061(n262 ,n59[1] ,n59[2]);
    not g2062(n1316 ,n1274);
    dff g2063(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1341), .Q(n10));
    nand g2064(n1260 ,n323 ,n1019);
    nand g2065(n1675 ,n39[4] ,n1483);
    dff g2066(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1203), .Q(n46[0]));
    nand g2067(n538 ,n30[6] ,n425);
    or g2068(n1945 ,n1880 ,n1879);
    dff g2069(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1260), .Q(n37[1]));
    nand g2070(n1233 ,n61[5] ,n887);
    dff g2071(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1174), .Q(n48[6]));
    nor g2072(n484 ,n193 ,n458);
    nand g2073(n1460 ,n53[0] ,n1375);
    nand g2074(n1214 ,n963 ,n753);
    not g2075(n202 ,n2244);
    nor g2076(n490 ,n193 ,n450);
    nor g2077(n2155 ,n1943 ,n2145);
    nand g2078(n2130 ,n526 ,n2119);
    nand g2079(n626 ,n33[2] ,n434);
    not g2080(n599 ,n531);
    nand g2081(n66 ,n19[1] ,n19[0]);
    not g2082(n1201 ,n1200);
    nand g2083(n1738 ,n36[1] ,n1466);
    not g2084(n133 ,n132);
    nand g2085(n1410 ,n42[3] ,n1376);
    nand g2086(n913 ,n51[4] ,n570);
    nand g2087(n811 ,n5[4] ,n580);
    nand g2088(n1519 ,n48[6] ,n1367);
    nand g2089(n2044 ,n1751 ,n1683);
    nand g2090(n1141 ,n901 ,n711);
    nor g2091(n422 ,n297 ,n402);
    dff g2092(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2042), .Q(n34[1]));
    nand g2093(n663 ,n25[4] ,n476);
    dff g2094(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1991), .Q(n25[0]));
    dff g2095(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1284), .Q(n57[0]));
    nand g2096(n1825 ,n21[3] ,n1495);
    nand g2097(n2032 ,n1745 ,n1686);
    nor g2098(n2217 ,n145 ,n147);
    dff g2099(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2011), .Q(n22[4]));
    not g2100(n344 ,n343);
    nor g2101(n1394 ,n448 ,n1347);
    or g2102(n2145 ,n1874 ,n2134);
    dff g2103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1982), .Q(n26[1]));
    nand g2104(n2045 ,n1752 ,n1684);
    nand g2105(n1293 ,n1061 ,n782);
    dff g2106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2131), .Q(n12[4]));
    nand g2107(n1780 ,n2199 ,n1498);
    nor g2108(n1368 ,n267 ,n1196);
    nand g2109(n614 ,n35[3] ,n435);
    nand g2110(n898 ,n20[6] ,n585);
    xnor g2111(n2205 ,n20[11] ,n182);
    nand g2112(n1266 ,n899 ,n778);
    nand g2113(n928 ,n605 ,n499);
    dff g2114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2094), .Q(n28[6]));
    nor g2115(n115 ,n20[11] ,n20[10]);
    nand g2116(n2008 ,n1814 ,n1621);
    nand g2117(n1985 ,n1790 ,n1599);
    nand g2118(n1982 ,n1787 ,n1596);
    nand g2119(n318 ,n12[4] ,n255);
    nand g2120(n2081 ,n898 ,n1916);
    nand g2121(n1139 ,n1052 ,n707);
    nand g2122(n2078 ,n1909 ,n1651);
    dff g2123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1182), .Q(n47[7]));
    nand g2124(n1722 ,n28[2] ,n1468);
    dff g2125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1219), .Q(n44[0]));
    nand g2126(n1036 ,n675 ,n543);
    nand g2127(n979 ,n42[5] ,n584);
    nand g2128(n1592 ,n39[5] ,n1474);
    nand g2129(n570 ,n263 ,n480);
    xnor g2130(n2197 ,n38[2] ,n187);
    nand g2131(n2093 ,n1772 ,n1706);
    not g2132(n201 ,n60[1]);
    dff g2133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1337), .Q(n14[1]));
    nand g2134(n1423 ,n54[7] ,n1373);
    nand g2135(n2063 ,n860 ,n1836);
    nand g2136(n1444 ,n46[2] ,n1374);
    nor g2137(n1363 ,n262 ,n1199);
    nand g2138(n674 ,n33[4] ,n434);
    nand g2139(n750 ,n5[1] ,n577);
    nand g2140(n971 ,n43[5] ,n562);
    not g2141(n199 ,n17[1]);
    nand g2142(n713 ,n5[3] ,n571);
    nand g2143(n986 ,n42[0] ,n584);
    nand g2144(n1813 ,n22[7] ,n1497);
    nand g2145(n668 ,n27[4] ,n424);
    not g2146(n699 ,n670);
    nand g2147(n1846 ,n1564 ,n1454);
    nand g2148(n2022 ,n1735 ,n1665);
    nand g2149(n1768 ,n29[3] ,n1470);
    not g2150(n307 ,n306);
    nand g2151(n1421 ,n55[4] ,n1370);
    or g2152(n250 ,n19[0] ,n19[1]);
    dff g2153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1984), .Q(n25[7]));
    dff g2154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1126), .Q(n40[0]));
    nand g2155(n1699 ,n39[7] ,n1471);
    nand g2156(n1707 ,n39[3] ,n1487);
    not g2157(n602 ,n549);
    nand g2158(n1178 ,n855 ,n821);
    nor g2159(n1371 ,n261 ,n1199);
    nand g2160(n1520 ,n56[6] ,n1377);
    nand g2161(n1164 ,n926 ,n729);
    nand g2162(n1114 ,n444 ,n888);
    not g2163(n223 ,n17[0]);
    nand g2164(n143 ,n40[1] ,n40[0]);
    dff g2165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1326), .Q(n8));
    nand g2166(n2051 ,n1920 ,n1716);
    nand g2167(n1715 ,n39[0] ,n1493);
    nand g2168(n1644 ,n39[2] ,n1488);
    dff g2169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2173), .Q(n61[4]));
    not g2170(n233 ,n58[4]);
    not g2171(n129 ,n128);
    nand g2172(n1153 ,n1022 ,n721);
    or g2173(n1940 ,n1866 ,n1865);
    nand g2174(n1265 ,n61[6] ,n887);
    nor g2175(n434 ,n268 ,n402);
    nand g2176(n609 ,n28[4] ,n432);
    nor g2177(n335 ,n2235 ,n302);
    dff g2178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n247), .Q(n7));
    nand g2179(n1425 ,n51[7] ,n1365);
    nand g2180(n1779 ,n2211 ,n1498);
    nand g2181(n1223 ,n972 ,n766);
    dff g2182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1232), .Q(n42[3]));
    nand g2183(n605 ,n28[2] ,n432);
    nand g2184(n651 ,n27[6] ,n424);
    nand g2185(n1535 ,n45[3] ,n1372);
    dff g2186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2015), .Q(n22[0]));
    dff g2187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n490), .Q(n39[0]));
    or g2188(n310 ,n17[2] ,n303);
    nand g2189(n1890 ,n32[5] ,n1489);
    nand g2190(n1204 ,n950 ,n745);
    nor g2191(n1471 ,n265 ,n1380);
    nor g2192(n364 ,n198 ,n328);
    dff g2193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2054), .Q(n32[5]));
    nand g2194(n1704 ,n39[2] ,n1471);
    nand g2195(n2094 ,n1773 ,n1708);
    nand g2196(n1669 ,n39[1] ,n1467);
    nand g2197(n1662 ,n240 ,n1498);
    nand g2198(n1116 ,n231 ,n889);
    dff g2199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1228), .Q(n42[7]));
    nand g2200(n606 ,n35[2] ,n435);
    nand g2201(n991 ,n469 ,n628);
    nand g2202(n1165 ,n846 ,n820);
    dff g2203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2004), .Q(n23[3]));
    nor g2204(n79 ,n78 ,n76);
    dff g2205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1136), .Q(n53[5]));
    nand g2206(n1820 ,n22[0] ,n1497);
    nand g2207(n1569 ,n54[1] ,n1373);
    nand g2208(n608 ,n32[2] ,n436);
    nand g2209(n2019 ,n1824 ,n1629);
    nand g2210(n1002 ,n460 ,n621);
    nand g2211(n1273 ,n398 ,n841);
    nand g2212(n1904 ,n30[7] ,n1485);
    nand g2213(n1337 ,n304 ,n1114);
    nand g2214(n920 ,n50[4] ,n574);
    nor g2215(n1348 ,n221 ,n1310);
    dff g2216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2071), .Q(n20[10]));
    dff g2217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1985), .Q(n25[6]));
    nand g2218(n824 ,n5[1] ,n576);
    nand g2219(n2055 ,n1893 ,n1642);
    nand g2220(n652 ,n36[0] ,n422);
    not g2221(n204 ,n38[3]);
    dff g2222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1976), .Q(n26[7]));
    dff g2223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2076), .Q(n30[4]));
    nand g2224(n467 ,n221 ,n410);
    nand g2225(n853 ,n48[6] ,n563);
    nand g2226(n1024 ,n55[7] ,n558);
    nand g2227(n936 ,n54[7] ,n582);
    nand g2228(n2021 ,n1741 ,n1664);
    dff g2229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1229), .Q(n42[6]));
    nand g2230(n349 ,n37[3] ,n255);
    nand g2231(n2065 ,n1759 ,n1694);
    nand g2232(n1229 ,n978 ,n767);
    nor g2233(n97 ,n40[2] ,n95);
    nand g2234(n983 ,n503 ,n508);
    nor g2235(n287 ,n238 ,n192);
    nor g2236(n2169 ,n597 ,n2162);
    nand g2237(n1220 ,n969 ,n758);
    nand g2238(n1891 ,n1513 ,n1408);
    nand g2239(n1871 ,n34[0] ,n1473);
    dff g2240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2068), .Q(n31[2]));
    nand g2241(n943 ,n46[4] ,n568);
    nand g2242(n1600 ,n39[5] ,n1476);
    nand g2243(n507 ,n61[1] ,n475);
    dff g2244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2024), .Q(n36[3]));
    dff g2245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2093), .Q(n28[7]));
    not g2246(n1494 ,n1495);
    nand g2247(n802 ,n5[4] ,n554);
    dff g2248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1511), .Q(n19[1]));
    dff g2249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1286), .Q(n56[6]));
    nand g2250(n734 ,n5[4] ,n565);
    not g2251(n216 ,n40[9]);
    nor g2252(n368 ,n220 ,n328);
    not g2253(n1086 ,n998);
    nor g2254(n491 ,n17[1] ,n416);
    nand g2255(n1307 ,n1045 ,n786);
    nand g2256(n1864 ,n1440 ,n1406);
    nand g2257(n1119 ,n38[2] ,n888);
    or g2258(n1587 ,n1335 ,n1392);
    nand g2259(n660 ,n32[5] ,n436);
    nand g2260(n1464 ,n42[0] ,n1376);
    nand g2261(n528 ,n23[4] ,n429);
    nand g2262(n763 ,n5[1] ,n561);
    dff g2263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1193), .Q(n53[3]));
    nand g2264(n1306 ,n1053 ,n798);
    nand g2265(n1623 ,n39[3] ,n1496);
    nand g2266(n646 ,n34[1] ,n426);
    nand g2267(n1190 ,n940 ,n738);
    nor g2268(n1509 ,n193 ,n1388);
    nand g2269(n1978 ,n1783 ,n1592);
    nand g2270(n831 ,n5[2] ,n576);
    nand g2271(n117 ,n20[1] ,n20[0]);
    nand g2272(n1001 ,n610 ,n514);
    dff g2273(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1149), .Q(n51[7]));
    nand g2274(n464 ,n40[4] ,n378);
    nor g2275(n1115 ,n939 ,n958);
    nand g2276(n2157 ,n1404 ,n2152);
    nand g2277(n1646 ,n39[7] ,n1484);
    nand g2278(n2080 ,n1914 ,n1661);
    not g2279(n242 ,n40[3]);
    nand g2280(n1203 ,n949 ,n744);
    nor g2281(n281 ,n231 ,n235);
    nand g2282(n107 ,n20[5] ,n20[4]);
    nand g2283(n1041 ,n50[5] ,n574);
    not g2284(n218 ,n39[7]);
    nor g2285(n894 ,n343 ,n590);
    or g2286(n1935 ,n1848 ,n1847);
    nand g2287(n1135 ,n2187 ,n893);
    nand g2288(n391 ,n60[0] ,n331);
    nand g2289(n1827 ,n21[1] ,n1495);
    nand g2290(n1960 ,n839 ,n1758);
    nor g2291(n285 ,n214 ,n193);
    nand g2292(n1320 ,n1130 ,n1262);
    nand g2293(n537 ,n29[1] ,n433);
    nand g2294(n866 ,n56[2] ,n575);
    nand g2295(n1528 ,n45[4] ,n1372);
    nand g2296(n1728 ,n27[4] ,n1482);
    nand g2297(n1406 ,n54[3] ,n1373);
    not g2298(n212 ,n11);
    or g2299(n1949 ,n1897 ,n1894);
    nand g2300(n393 ,n246 ,n356);
    nand g2301(n70 ,n2207 ,n64);
    nand g2302(n276 ,n199 ,n221);
    nand g2303(n929 ,n662 ,n501);
    or g2304(n2141 ,n1839 ,n2133);
    nor g2305(n67 ,n2207 ,n66);
    nand g2306(n1667 ,n39[3] ,n1467);
    nand g2307(n1967 ,n1725 ,n1672);
    dff g2308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1254), .Q(n46[1]));
    nand g2309(n1342 ,n1124 ,n1116);
    nand g2310(n948 ,n613 ,n537);
    nand g2311(n2082 ,n1764 ,n1699);
    nand g2312(n1714 ,n39[0] ,n1483);
    nand g2313(n729 ,n5[0] ,n573);
    nand g2314(n1823 ,n21[5] ,n1495);
    nand g2315(n2137 ,n1506 ,n2109);
    nor g2316(n450 ,n368 ,n371);
    nor g2317(n280 ,n239 ,n192);
    nand g2318(n1415 ,n346 ,n1354);
    nor g2319(n116 ,n20[4] ,n20[3]);
    nand g2320(n954 ,n45[4] ,n578);
    nand g2321(n1788 ,n26[0] ,n1475);
    nand g2322(n1807 ,n23[5] ,n1481);
    nand g2323(n1702 ,n39[4] ,n1471);
    dff g2324(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1285), .Q(n56[7]));
    nor g2325(n253 ,n206 ,n17[0]);
    dff g2326(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n282), .Q(n16[7]));
    dff g2327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1170), .Q(n49[2]));
    nand g2328(n1018 ,n655 ,n654);
    nand g2329(n1288 ,n876 ,n829);
    nand g2330(n2009 ,n1813 ,n1619);
    nand g2331(n1451 ,n42[7] ,n1376);
    nand g2332(n1889 ,n32[6] ,n1489);
    nand g2333(n1659 ,n39[0] ,n1494);
    nand g2334(n2090 ,n1769 ,n1704);
    nor g2335(n2181 ,n2185 ,n17[1]);
    nand g2336(n998 ,n463 ,n634);
    dff g2337(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2091), .Q(n29[1]));
    nor g2338(n283 ,n236 ,n192);
    dff g2339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n453), .Q(n13[2]));
    nand g2340(n1759 ,n31[4] ,n1490);
    nand g2341(n1404 ,n51[3] ,n1365);
    nand g2342(n385 ,n314 ,n322);
    nand g2343(n524 ,n31[6] ,n427);
    nor g2344(n453 ,n207 ,n405);
    not g2345(n579 ,n580);
    nand g2346(n1548 ,n49[1] ,n1369);
    nand g2347(n2104 ,n1825 ,n1630);
    nand g2348(n1075 ,n57[0] ,n553);
    dff g2349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2006), .Q(n23[1]));
    nand g2350(n2177 ,n1515 ,n2171);
    not g2351(n225 ,n60[2]);
    nor g2352(n1340 ,n871 ,n1111);
    buf g2353(n13[0], 1'b0);
    dff g2354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2044), .Q(n33[7]));
    dff g2355(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2000), .Q(n23[7]));
    nand g2356(n2000 ,n1805 ,n1612);
    not g2357(n592 ,n591);
    nand g2358(n1457 ,n54[0] ,n1373);
    nand g2359(n828 ,n5[5] ,n576);
    nand g2360(n978 ,n42[6] ,n584);
    not g2361(n232 ,n62[1]);
    nand g2362(n956 ,n45[3] ,n578);
    dff g2363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1247), .Q(n40[8]));
    nand g2364(n394 ,n6 ,n345);
    or g2365(n1095 ,n994 ,n990);
    dff g2366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2177), .Q(n61[2]));
    nand g2367(n2087 ,n1034 ,n1915);
    nand g2368(n863 ,n49[0] ,n579);
    nand g2369(n703 ,n5[5] ,n559);
    not g2370(n553 ,n554);
    nor g2371(n102 ,n96 ,n101);
    nand g2372(n1209 ,n1049 ,n749);
    dff g2373(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1294), .Q(n55[5]));
    nand g2374(n1770 ,n29[1] ,n1470);
    nand g2375(n1049 ,n45[2] ,n578);
    nor g2376(n316 ,n17[2] ,n253);
    or g2377(n1927 ,n1891 ,n1832);
    nand g2378(n1150 ,n911 ,n718);
    nand g2379(n1447 ,n42[1] ,n1376);
    nor g2380(n255 ,n193 ,n2242);
    nand g2381(n1543 ,n49[2] ,n1369);
    dff g2382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1308), .Q(n40[1]));
    dff g2383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2062), .Q(n20[12]));
    nand g2384(n502 ,n22[5] ,n423);
    dff g2385(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2090), .Q(n29[2]));
    nand g2386(n1923 ,n33[3] ,n1486);
    nand g2387(n2005 ,n1810 ,n1617);
    nand g2388(n743 ,n5[5] ,n577);
    not g2389(n336 ,n335);
    nand g2390(n303 ,n17[0] ,n2210);
    nand g2391(n1685 ,n39[5] ,n1487);
    nand g2392(n870 ,n57[5] ,n553);
    nand g2393(n514 ,n29[7] ,n433);
    nand g2394(n2017 ,n1822 ,n1627);
    nand g2395(n1748 ,n1333 ,n1529);
    nand g2396(n508 ,n21[0] ,n430);
    nor g2397(n1353 ,n1096 ,n1094);
    not g2398(n557 ,n558);
    nand g2399(n1783 ,n26[5] ,n1475);
    nand g2400(n1439 ,n50[3] ,n1364);
    nand g2401(n1227 ,n976 ,n764);
    nand g2402(n348 ,n12[5] ,n255);
    nand g2403(n297 ,n37[0] ,n37[1]);
    dff g2404(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n305), .Q(n13[1]));
    nand g2405(n1550 ,n45[0] ,n1372);
    nor g2406(n1379 ,n38[3] ,n1202);
    dff g2407(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1297), .Q(n54[1]));
    nor g2408(n1357 ,n222 ,n1195);
    or g2409(n799 ,n325 ,n676);
    dff g2410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1267), .Q(n56[0]));
    nor g2411(n2196 ,n188 ,n186);
    nor g2412(n1579 ,n927 ,n1402);
    nand g2413(n1027 ,n684 ,n532);
    nand g2414(n2103 ,n1827 ,n1632);
    nand g2415(n1554 ,n56[0] ,n1377);
    nand g2416(n271 ,n38[1] ,n228);
    dff g2417(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1207), .Q(n45[4]));
    nand g2418(n1525 ,n47[5] ,n1371);
    nor g2419(n451 ,n360 ,n376);
    nand g2420(n1176 ,n61[3] ,n887);
    nand g2421(n736 ,n5[1] ,n565);
    nand g2422(n1950 ,n1117 ,n1579);
    dff g2423(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2014), .Q(n22[1]));
    dff g2424(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1992), .Q(n24[7]));
    nand g2425(n1074 ,n56[7] ,n575);
    nand g2426(n1791 ,n25[4] ,n1477);
    nor g2427(n295 ,n241 ,n192);
    nand g2428(n531 ,n61[6] ,n475);
    nand g2429(n610 ,n27[7] ,n424);
    nand g2430(n974 ,n43[2] ,n562);
    nand g2431(n1660 ,n39[0] ,n1488);
    nand g2432(n1886 ,n32[7] ,n1489);
    nand g2433(n666 ,n387 ,n413);
    nand g2434(n1324 ,n1243 ,n1242);
    dff g2435(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1204), .Q(n45[7]));
    nand g2436(n1043 ,n47[1] ,n566);
    nand g2437(n687 ,n36[2] ,n422);
    nor g2438(n1395 ,n193 ,n1361);
    nor g2439(n2112 ,n1948 ,n1947);
    dff g2440(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1150), .Q(n51[6]));
    nand g2441(n1228 ,n977 ,n765);
    nand g2442(n838 ,n257 ,n492);
    nand g2443(n1689 ,n39[1] ,n1487);
    nand g2444(n1901 ,n1524 ,n1576);
    nand g2445(n2077 ,n1908 ,n1650);
    nand g2446(n350 ,n12[6] ,n255);
    nand g2447(n1866 ,n1405 ,n1403);
    nand g2448(n1235 ,n985 ,n730);
    not g2449(n1472 ,n1473);
    nand g2450(n1753 ,n33[5] ,n1486);
    nor g2451(n321 ,n58[1] ,n279);
    dff g2452(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2047), .Q(n33[4]));
    nand g2453(n861 ,n58[2] ,n589);
    nor g2454(n594 ,n477 ,n445);
    xnor g2455(n2220 ,n40[6] ,n150);
    not g2456(n191 ,n190);
    nor g2457(n1393 ,n1357 ,n1358);
    dff g2458(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2036), .Q(n34[7]));
    nor g2459(n120 ,n20[2] ,n118);
    nand g2460(n877 ,n58[3] ,n589);
    nand g2461(n1057 ,n55[2] ,n558);
    nand g2462(n2041 ,n1867 ,n1598);
    nand g2463(n1380 ,n38[3] ,n1200);
    nand g2464(n1894 ,n1556 ,n1271);
    not g2465(n896 ,n895);
    nand g2466(n2062 ,n879 ,n1900);
    nor g2467(n123 ,n114 ,n122);
    dff g2468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1211), .Q(n45[0]));
    nand g2469(n1191 ,n1039 ,n739);
    dff g2470(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1187), .Q(n47[2]));
    nand g2471(n739 ,n5[6] ,n567);
    nand g2472(n1000 ,n464 ,n635);
    dff g2473(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1987), .Q(n25[4]));
    not g2474(n230 ,n37[1]);
    nor g2475(n179 ,n20[9] ,n178);
    nand g2476(n970 ,n43[6] ,n562);
    dff g2477(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1281), .Q(n57[2]));
    nand g2478(n937 ,n47[2] ,n566);
    nand g2479(n1611 ,n39[1] ,n1478);
    nand g2480(n1762 ,n31[1] ,n1490);
    nor g2481(n445 ,n320 ,n390);
    nand g2482(n661 ,n35[5] ,n435);
    nand g2483(n907 ,n689 ,n548);
    dff g2484(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2078), .Q(n30[2]));
    not g2485(n217 ,n39[6]);
    nand g2486(n688 ,n32[1] ,n436);
    not g2487(n176 ,n175);
    dff g2488(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1175), .Q(n48[5]));
    dff g2489(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1306), .Q(n54[0]));
    nor g2490(n425 ,n270 ,n380);
    nand g2491(n642 ,n28[7] ,n432);
    nor g2492(n2203 ,n179 ,n181);
    nand g2493(n1278 ,n870 ,n805);
    nand g2494(n950 ,n45[7] ,n578);
    nand g2495(n1257 ,n38[0] ,n888);
    nand g2496(n2138 ,n1562 ,n2108);
    nand g2497(n2095 ,n1774 ,n1709);
    not g2498(n200 ,n59[0]);
    nand g2499(n868 ,n20[10] ,n585);
    nand g2500(n1912 ,n1427 ,n1570);
    nand g2501(n989 ,n461 ,n630);
    nand g2502(n1256 ,n1056 ,n791);
    not g2503(n149 ,n148);
    nand g2504(n1802 ,n24[2] ,n1479);
    nand g2505(n784 ,n5[6] ,n573);
    nand g2506(n1240 ,n41[2] ,n890);
    nand g2507(n1549 ,n57[1] ,n1362);
    nand g2508(n1648 ,n39[5] ,n1484);
    not g2509(n196 ,n39[3]);
    nand g2510(n1449 ,n53[1] ,n1375);
    dff g2511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2124), .Q(n12[3]));
    nand g2512(n1409 ,n44[3] ,n1366);
    nor g2513(n416 ,n17[2] ,n410);
    nor g2514(n131 ,n58[1] ,n58[0]);
    nand g2515(n1047 ,n678 ,n534);
    nand g2516(n1071 ,n56[1] ,n575);
    nand g2517(n731 ,n5[7] ,n565);
    nand g2518(n694 ,n26[6] ,n431);
    not g2519(n203 ,n38[1]);
    nand g2520(n1329 ,n1050 ,n1314);
    nand g2521(n2047 ,n1584 ,n1687);
    dff g2522(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1290), .Q(n56[2]));
    nand g2523(n1061 ,n55[6] ,n558);
    nand g2524(n1597 ,n39[7] ,n1476);
    nor g2525(n1493 ,n298 ,n1380);
    dff g2526(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1142), .Q(n52[6]));
    nand g2527(n1286 ,n875 ,n827);
    nand g2528(n1034 ,n20[7] ,n585);
    nand g2529(n259 ,n38[2] ,n203);
    dff g2530(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2067), .Q(n20[11]));
    nand g2531(n636 ,n2216 ,n421);
    nand g2532(n1009 ,n641 ,n519);
    not g2533(n164 ,n20[8]);
    not g2534(n169 ,n168);
    not g2535(n332 ,n333);
    dff g2536(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2041), .Q(n34[2]));
    nand g2537(n846 ,n49[7] ,n579);
    dff g2538(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2021), .Q(n36[6]));
    nand g2539(n1773 ,n28[6] ,n1468);
    nand g2540(n1242 ,n2233 ,n889);
    nand g2541(n623 ,n25[0] ,n476);
    nor g2542(n1091 ,n965 ,n955);
    dff g2543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2129), .Q(n12[6]));
    nand g2544(n1224 ,n973 ,n761);
    or g2545(n71 ,n19[2] ,n70);
    xnor g2546(n2198 ,n38[3] ,n189);
    nand g2547(n2028 ,n1740 ,n1679);
    dff g2548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1967), .Q(n27[7]));
    dff g2549(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1227), .Q(n43[0]));
    dff g2550(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2030), .Q(n35[5]));
    nand g2551(n809 ,n5[5] ,n580);
    nand g2552(n1658 ,n39[0] ,n1496);
    nand g2553(n574 ,n263 ,n440);
    nand g2554(n766 ,n5[4] ,n561);
    nand g2555(n1302 ,n1062 ,n783);
    nand g2556(n1561 ,n49[6] ,n1369);
    or g2557(n89 ,n19[4] ,n19[1]);
    nor g2558(n269 ,n201 ,n60[2]);
    dff g2559(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1282), .Q(n57[1]));
    nand g2560(n662 ,n24[5] ,n428);
    nand g2561(n1602 ,n39[3] ,n1476);
    nand g2562(n807 ,n5[1] ,n554);
    dff g2563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1979), .Q(n26[4]));
    dff g2564(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2039), .Q(n34[4]));
    xnor g2565(n2194 ,n37[2] ,n160);
    xnor g2566(n2222 ,n40[8] ,n153);
    nand g2567(n346 ,n12[0] ,n255);
    nand g2568(n673 ,n25[5] ,n476);
    nand g2569(n1701 ,n39[5] ,n1471);
endmodule
