module top (n0, n1, n5, n6, n2, n3, n9, n14, n15, n7, n8, n4, n16, n17, n10, n11, n12, n13);
    input n0, n1, n2, n3, n4;
    input [31:0] n5, n6;
    input [3:0] n7;
    input [1:0] n8;
    output [31:0] n9, n10, n11, n12, n13;
    output n14, n15, n16;
    output [7:0] n17;
    wire n0, n1, n2, n3, n4;
    wire [31:0] n5, n6;
    wire [3:0] n7;
    wire [1:0] n8;
    wire [31:0] n9, n10, n11, n12, n13;
    wire n14, n15, n16;
    wire [7:0] n17;
    wire [2:0] n18;
    wire [7:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [7:0] n23;
    wire [7:0] n24;
    wire [7:0] n25;
    wire [15:0] n26;
    wire [1:0] n27;
    wire [15:0] n28;
    wire [15:0] n29;
    wire [7:0] n30;
    wire [15:0] n31;
    wire [15:0] n32;
    wire n33, n34, n35, n36, n37, n38, n39, n40;
    wire n41, n42, n43, n44, n45, n46, n47, n48;
    wire n49, n50, n51, n52, n53, n54, n55, n56;
    wire n57, n58, n59, n60, n61, n62, n63, n64;
    wire n65, n66, n67, n68, n69, n70, n71, n72;
    wire n73, n74, n75, n76, n77, n78, n79, n80;
    wire n81, n82, n83, n84, n85, n86, n87, n88;
    wire n89, n90, n91, n92, n93, n94, n95, n96;
    wire n97, n98, n99, n100, n101, n102, n103, n104;
    wire n105, n106, n107, n108, n109, n110, n111, n112;
    wire n113, n114, n115, n116, n117, n118, n119, n120;
    wire n121, n122, n123, n124, n125, n126, n127, n128;
    wire n129, n130, n131, n132, n133, n134, n135, n136;
    wire n137, n138, n139, n140, n141, n142, n143, n144;
    wire n145, n146, n147, n148, n149, n150, n151, n152;
    wire n153, n154, n155, n156, n157, n158, n159, n160;
    wire n161, n162, n163, n164, n165, n166, n167, n168;
    wire n169, n170, n171, n172, n173, n174, n175, n176;
    wire n177, n178, n179, n180, n181, n182, n183, n184;
    wire n185, n186, n187, n188, n189, n190, n191, n192;
    wire n193, n194, n195, n196, n197, n198, n199, n200;
    wire n201, n202, n203, n204, n205, n206, n207, n208;
    wire n209, n210, n211, n212, n213, n214, n215, n216;
    wire n217, n218, n219, n220, n221, n222, n223, n224;
    wire n225, n226, n227, n228, n229, n230, n231, n232;
    wire n233, n234, n235, n236, n237, n238, n239, n240;
    wire n241, n242, n243, n244, n245, n246, n247, n248;
    wire n249, n250, n251, n252, n253, n254, n255, n256;
    wire n257, n258, n259, n260, n261, n262, n263, n264;
    wire n265, n266, n267, n268, n269, n270, n271, n272;
    wire n273, n274, n275, n276, n277, n278, n279, n280;
    wire n281, n282, n283, n284, n285, n286, n287, n288;
    wire n289, n290, n291, n292, n293, n294, n295, n296;
    wire n297, n298, n299, n300, n301, n302, n303, n304;
    wire n305, n306, n307, n308, n309, n310, n311, n312;
    wire n313, n314, n315, n316, n317, n318, n319, n320;
    wire n321, n322, n323, n324, n325, n326, n327, n328;
    wire n329, n330, n331, n332, n333, n334, n335, n336;
    wire n337, n338, n339, n340, n341, n342, n343, n344;
    wire n345, n346, n347, n348, n349, n350, n351, n352;
    wire n353, n354, n355, n356, n357, n358, n359, n360;
    wire n361, n362, n363, n364, n365, n366, n367, n368;
    wire n369, n370, n371, n372, n373, n374, n375, n376;
    wire n377, n378, n379, n380, n381, n382, n383, n384;
    wire n385, n386, n387, n388, n389, n390, n391, n392;
    wire n393, n394, n395, n396, n397, n398, n399, n400;
    wire n401, n402, n403, n404, n405, n406, n407, n408;
    wire n409, n410, n411, n412, n413, n414, n415, n416;
    wire n417, n418, n419, n420, n421, n422, n423, n424;
    wire n425, n426, n427, n428, n429, n430, n431, n432;
    wire n433, n434, n435, n436, n437, n438, n439, n440;
    wire n441, n442, n443, n444, n445, n446, n447, n448;
    wire n449, n450, n451, n452, n453, n454, n455, n456;
    wire n457, n458, n459, n460, n461, n462, n463, n464;
    wire n465, n466, n467, n468, n469, n470, n471, n472;
    wire n473, n474, n475, n476, n477, n478, n479, n480;
    wire n481, n482, n483, n484, n485, n486, n487, n488;
    wire n489, n490, n491, n492, n493, n494, n495, n496;
    wire n497, n498, n499, n500, n501, n502, n503, n504;
    wire n505, n506, n507, n508, n509, n510, n511, n512;
    wire n513, n514, n515, n516, n517, n518, n519, n520;
    wire n521, n522, n523, n524, n525, n526, n527, n528;
    wire n529, n530, n531, n532, n533, n534, n535, n536;
    wire n537, n538, n539, n540, n541, n542, n543, n544;
    wire n545, n546, n547, n548, n549, n550, n551, n552;
    wire n553, n554, n555, n556, n557, n558, n559, n560;
    wire n561, n562, n563, n564, n565, n566, n567, n568;
    wire n569, n570, n571, n572, n573, n574, n575, n576;
    wire n577, n578, n579, n580, n581, n582, n583, n584;
    wire n585, n586, n587, n588, n589, n590, n591, n592;
    wire n593, n594, n595, n596, n597, n598, n599, n600;
    wire n601, n602, n603, n604, n605, n606, n607, n608;
    wire n609, n610, n611, n612, n613, n614, n615, n616;
    wire n617, n618, n619, n620, n621, n622, n623, n624;
    wire n625, n626, n627, n628, n629, n630, n631, n632;
    wire n633, n634, n635, n636, n637, n638, n639, n640;
    wire n641, n642, n643, n644, n645, n646, n647, n648;
    wire n649, n650, n651, n652, n653, n654, n655, n656;
    wire n657, n658, n659, n660, n661, n662, n663, n664;
    wire n665, n666, n667, n668, n669, n670, n671, n672;
    wire n673, n674, n675, n676, n677, n678, n679, n680;
    wire n681, n682, n683, n684, n685, n686, n687, n688;
    wire n689, n690, n691, n692, n693, n694, n695, n696;
    wire n697, n698, n699, n700, n701, n702, n703, n704;
    wire n705, n706, n707, n708, n709, n710, n711, n712;
    wire n713, n714, n715, n716, n717, n718, n719, n720;
    wire n721, n722, n723, n724, n725, n726, n727, n728;
    wire n729, n730, n731, n732, n733, n734, n735, n736;
    wire n737, n738, n739, n740, n741, n742, n743, n744;
    wire n745, n746, n747, n748, n749, n750, n751, n752;
    wire n753, n754, n755, n756, n757, n758, n759, n760;
    wire n761, n762, n763, n764, n765, n766, n767, n768;
    wire n769, n770, n771, n772, n773, n774, n775, n776;
    wire n777, n778, n779, n780, n781, n782, n783, n784;
    wire n785, n786, n787, n788, n789, n790, n791, n792;
    wire n793, n794, n795, n796, n797, n798, n799, n800;
    wire n801, n802, n803, n804, n805, n806, n807, n808;
    wire n809, n810, n811, n812, n813, n814, n815, n816;
    wire n817, n818, n819, n820, n821, n822, n823, n824;
    wire n825, n826, n827, n828, n829, n830, n831, n832;
    wire n833, n834, n835, n836, n837, n838, n839, n840;
    wire n841, n842, n843, n844, n845, n846, n847, n848;
    wire n849, n850, n851, n852, n853, n854, n855, n856;
    wire n857, n858, n859, n860, n861, n862, n863, n864;
    wire n865, n866, n867, n868, n869, n870, n871, n872;
    wire n873, n874, n875, n876, n877, n878, n879, n880;
    wire n881, n882, n883, n884, n885, n886, n887, n888;
    wire n889, n890, n891, n892, n893, n894, n895, n896;
    wire n897, n898, n899, n900, n901, n902, n903, n904;
    wire n905, n906, n907, n908, n909, n910, n911, n912;
    wire n913, n914, n915, n916, n917, n918, n919, n920;
    wire n921, n922, n923, n924, n925, n926, n927, n928;
    wire n929, n930, n931, n932, n933, n934, n935, n936;
    wire n937, n938, n939, n940, n941, n942, n943, n944;
    wire n945, n946, n947, n948, n949, n950, n951, n952;
    wire n953, n954, n955, n956, n957, n958, n959, n960;
    wire n961, n962, n963, n964, n965, n966, n967, n968;
    wire n969, n970, n971, n972, n973, n974, n975, n976;
    wire n977, n978, n979, n980, n981, n982, n983, n984;
    wire n985, n986, n987, n988, n989, n990, n991, n992;
    wire n993, n994, n995, n996, n997, n998, n999, n1000;
    wire n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008;
    wire n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016;
    wire n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
    wire n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
    wire n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040;
    wire n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
    wire n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056;
    wire n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064;
    wire n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072;
    wire n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080;
    wire n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088;
    wire n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096;
    wire n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104;
    wire n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112;
    wire n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120;
    wire n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128;
    wire n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136;
    wire n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144;
    wire n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152;
    wire n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160;
    wire n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168;
    wire n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176;
    wire n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184;
    wire n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192;
    wire n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200;
    wire n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208;
    wire n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216;
    wire n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224;
    wire n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232;
    wire n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240;
    wire n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248;
    wire n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256;
    wire n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264;
    wire n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272;
    wire n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;
    wire n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288;
    wire n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296;
    wire n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304;
    wire n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312;
    wire n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320;
    wire n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;
    wire n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336;
    wire n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344;
    wire n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352;
    wire n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360;
    wire n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368;
    wire n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376;
    wire n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384;
    wire n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392;
    wire n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400;
    wire n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408;
    wire n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416;
    wire n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424;
    wire n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432;
    wire n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440;
    wire n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448;
    wire n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456;
    wire n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464;
    wire n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472;
    wire n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480;
    wire n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488;
    wire n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496;
    wire n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504;
    wire n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512;
    wire n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520;
    wire n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528;
    wire n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536;
    wire n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544;
    wire n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552;
    wire n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560;
    wire n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568;
    wire n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576;
    wire n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584;
    wire n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592;
    wire n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600;
    wire n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608;
    wire n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616;
    wire n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624;
    wire n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632;
    wire n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640;
    wire n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648;
    wire n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656;
    wire n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664;
    wire n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672;
    wire n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680;
    wire n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688;
    wire n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696;
    wire n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704;
    wire n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712;
    wire n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720;
    wire n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728;
    wire n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736;
    wire n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744;
    wire n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752;
    wire n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760;
    wire n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768;
    wire n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776;
    wire n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784;
    wire n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792;
    wire n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800;
    wire n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808;
    wire n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816;
    wire n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824;
    wire n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832;
    wire n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840;
    wire n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848;
    wire n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856;
    wire n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864;
    wire n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872;
    wire n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880;
    wire n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888;
    wire n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896;
    wire n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904;
    wire n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912;
    wire n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920;
    wire n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928;
    wire n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936;
    wire n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944;
    wire n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952;
    wire n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960;
    wire n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968;
    wire n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976;
    wire n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984;
    wire n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992;
    wire n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000;
    wire n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008;
    wire n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016;
    wire n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024;
    wire n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032;
    wire n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040;
    wire n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048;
    wire n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056;
    wire n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064;
    wire n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072;
    wire n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080;
    wire n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088;
    wire n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096;
    wire n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104;
    wire n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112;
    wire n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120;
    wire n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128;
    wire n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136;
    wire n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144;
    wire n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152;
    wire n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160;
    wire n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168;
    wire n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176;
    wire n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184;
    wire n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192;
    wire n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200;
    wire n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208;
    wire n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216;
    wire n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224;
    wire n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232;
    wire n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240;
    wire n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248;
    wire n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256;
    wire n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264;
    wire n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272;
    wire n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280;
    wire n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288;
    wire n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296;
    wire n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304;
    wire n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312;
    wire n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320;
    wire n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328;
    wire n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336;
    wire n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344;
    wire n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352;
    wire n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360;
    wire n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368;
    wire n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376;
    wire n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384;
    wire n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392;
    wire n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400;
    wire n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408;
    wire n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416;
    wire n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424;
    wire n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432;
    wire n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440;
    wire n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448;
    wire n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456;
    wire n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464;
    wire n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472;
    wire n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480;
    wire n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488;
    wire n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496;
    wire n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504;
    wire n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512;
    wire n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520;
    wire n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528;
    wire n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536;
    wire n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544;
    wire n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552;
    wire n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560;
    wire n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568;
    wire n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576;
    wire n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584;
    wire n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592;
    wire n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600;
    wire n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608;
    wire n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616;
    wire n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624;
    wire n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632;
    wire n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640;
    wire n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648;
    wire n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656;
    wire n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664;
    wire n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672;
    wire n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680;
    wire n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688;
    wire n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696;
    wire n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704;
    wire n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712;
    wire n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720;
    wire n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728;
    wire n2729, n2730, n2731;
    nand g0(n1660 ,n20[0] ,n22[4]);
    nor g1(n974 ,n929 ,n928);
    buf g2(n9[24], 1'b0);
    xnor g3(n1968 ,n1818 ,n1593);
    nand g4(n2389 ,n2336 ,n2370);
    xnor g5(n1068 ,n958 ,n1012);
    dff g6(.RN(n1), .SN(1'b1), .CK(n0), .D(n662), .Q(n19[2]));
    nand g7(n2048 ,n1912 ,n1996);
    xnor g8(n1864 ,n1619 ,n1616);
    nand g9(n1701 ,n20[5] ,n22[1]);
    xnor g10(n779 ,n21[2] ,n21[1]);
    xnor g11(n2377 ,n2352 ,n2280);
    nand g12(n520 ,n6[5] ,n475);
    nor g13(n1153 ,n1099 ,n1122);
    or g14(n2071 ,n1872 ,n1989);
    nor g15(n1229 ,n1212 ,n1188);
    xnor g16(n1829 ,n1685 ,n1573);
    dff g17(.RN(n1), .SN(1'b1), .CK(n0), .D(n362), .Q(n29[11]));
    nor g18(n1323 ,n1268 ,n1280);
    dff g19(.RN(n1), .SN(1'b1), .CK(n0), .D(n732), .Q(n9[4]));
    nand g20(n560 ,n24[4] ,n461);
    nand g21(n274 ,n31[13] ,n141);
    nand g22(n221 ,n26[7] ,n140);
    xnor g23(n2129 ,n2025 ,n1987);
    nand g24(n856 ,n2717 ,n825);
    buf g25(n11[15], 1'b0);
    xnor g26(n2181 ,n2091 ,n1978);
    or g27(n1256 ,n1236 ,n1255);
    xnor g28(n2692 ,n2410 ,n2430);
    nor g29(n2544 ,n2721 ,n32[12]);
    nor g30(n1955 ,n1726 ,n1903);
    not g31(n1631 ,n1630);
    nand g32(n835 ,n2717 ,n820);
    nand g33(n1574 ,n20[6] ,n22[6]);
    nand g34(n2226 ,n2145 ,n2184);
    nand g35(n558 ,n24[7] ,n461);
    not g36(n2498 ,n2497);
    nand g37(n1086 ,n757 ,n1029);
    nand g38(n1805 ,n1685 ,n1573);
    buf g39(n9[19], 1'b0);
    dff g40(.RN(n1), .SN(1'b1), .CK(n0), .D(n660), .Q(n19[3]));
    nand g41(n2119 ,n2005 ,n2073);
    nand g42(n2009 ,n1656 ,n1946);
    nand g43(n2308 ,n2153 ,n2287);
    buf g44(n12[8], n10[0]);
    nand g45(n262 ,n25[1] ,n142);
    nand g46(n2350 ,n2309 ,n2331);
    nor g47(n466 ,n344 ,n459);
    nor g48(n760 ,n20[5] ,n21[5]);
    xnor g49(n2708 ,n1243 ,n1255);
    nand g50(n515 ,n6[4] ,n462);
    or g51(n2405 ,n2388 ,n2395);
    nor g52(n169 ,n150 ,n148);
    buf g53(n12[26], 1'b0);
    xnor g54(n1223 ,n1191 ,n1202);
    nand g55(n1257 ,n1256 ,n1235);
    xnor g56(n1076 ,n1019 ,n980);
    not g57(n463 ,n464);
    nor g58(n1169 ,n1148 ,n1116);
    xnor g59(n1435 ,n1374 ,n1390);
    nand g60(n2435 ,n2367 ,n2434);
    nand g61(n1509 ,n1501 ,n1499);
    nand g62(n428 ,n327 ,n246);
    nand g63(n116 ,n5[3] ,n5[2]);
    nand g64(n160 ,n18[0] ,n108);
    nand g65(n1912 ,n1806 ,n1855);
    nor g66(n1322 ,n1268 ,n1279);
    nor g67(n2542 ,n2727 ,n32[6]);
    nand g68(n1541 ,n1523 ,n1530);
    not g69(n2190 ,n2189);
    nand g70(n618 ,n22[2] ,n469);
    nor g71(n1314 ,n1266 ,n1280);
    nand g72(n1649 ,n21[0] ,n23[0]);
    xnor g73(n1010 ,n951 ,n817);
    xnor g74(n2023 ,n1927 ,n1937);
    nand g75(n195 ,n29[1] ,n87);
    xnor g76(n1072 ,n998 ,n962);
    xnor g77(n2701 ,n1164 ,n1204);
    xnor g78(n1835 ,n1584 ,n1677);
    or g79(n1419 ,n1370 ,n1388);
    nand g80(n1610 ,n21[5] ,n23[4]);
    xnor g81(n1021 ,n816 ,n937);
    nand g82(n883 ,n2712 ,n846);
    buf g83(n12[10], n10[2]);
    xnor g84(n1526 ,n1481 ,n1508);
    nand g85(n234 ,n29[7] ,n87);
    not g86(n1393 ,n1392);
    xnor g87(n1142 ,n1096 ,n1101);
    or g88(n1272 ,n2679 ,n23[7]);
    nand g89(n1361 ,n24[0] ,n1299);
    nand g90(n531 ,n6[1] ,n470);
    nand g91(n121 ,n18[0] ,n18[1]);
    nand g92(n2246 ,n2156 ,n2208);
    nand g93(n398 ,n224 ,n343);
    xnor g94(n1434 ,n1372 ,n1395);
    nor g95(n1329 ,n1267 ,n1283);
    nand g96(n792 ,n2713 ,n783);
    nor g97(n1155 ,n1135 ,n1125);
    nor g98(n1321 ,n1268 ,n1281);
    not g99(n2533 ,n27[0]);
    not g100(n59 ,n58);
    dff g101(.RN(n1), .SN(1'b1), .CK(n0), .D(n361), .Q(n29[9]));
    nand g102(n1583 ,n20[5] ,n22[7]);
    nand g103(n2202 ,n2121 ,n2143);
    nand g104(n1603 ,n20[0] ,n22[7]);
    nand g105(n1778 ,n1589 ,n1652);
    not g106(n1011 ,n1010);
    nor g107(n716 ,n673 ,n672);
    nand g108(n704 ,n630 ,n631);
    nand g109(n1886 ,n1614 ,n1774);
    nor g110(n74 ,n25[5] ,n73);
    nand g111(n351 ,n234 ,n176);
    nand g112(n1708 ,n21[3] ,n23[2]);
    nand g113(n253 ,n126 ,n133);
    nand g114(n486 ,n6[0] ,n466);
    nand g115(n865 ,n2713 ,n824);
    nand g116(n2358 ,n2285 ,n2343);
    nor g117(n1353 ,n1266 ,n1304);
    nand g118(n2652 ,n2587 ,n2586);
    nand g119(n2336 ,n2268 ,n2301);
    dff g120(.RN(n1), .SN(1'b1), .CK(n0), .D(n658), .Q(n19[5]));
    nand g121(n891 ,n2715 ,n846);
    xor g122(n2030 ,n1949 ,n1935);
    nand g123(n1910 ,n1807 ,n1857);
    not g124(n1114 ,n1113);
    xnor g125(n747 ,n25[2] ,n68);
    nand g126(n1235 ,n1220 ,n1231);
    nand g127(n298 ,n29[4] ,n141);
    nand g128(n31[14] ,n2607 ,n2653);
    nand g129(n644 ,n538 ,n483);
    xnor g130(n2193 ,n2092 ,n2020);
    nand g131(n2560 ,n27[1] ,n27[0]);
    not g132(n54 ,n30[4]);
    not g133(n142 ,n143);
    buf g134(n13[1], 1'b0);
    xnor g135(n32[6] ,n1539 ,n1551);
    nand g136(n528 ,n6[3] ,n479);
    dff g137(.RN(n1), .SN(1'b1), .CK(n0), .D(n447), .Q(n14));
    not g138(n1039 ,n1032);
    nand g139(n423 ,n321 ,n240);
    nand g140(n1381 ,n1333 ,n1346);
    nand g141(n2477 ,n2707 ,n2691);
    dff g142(.RN(n1), .SN(1'b1), .CK(n0), .D(n379), .Q(n28[2]));
    nand g143(n218 ,n26[11] ,n140);
    xnor g144(n2092 ,n2017 ,n2013);
    nand g145(n191 ,n29[6] ,n87);
    nand g146(n333 ,n28[15] ,n141);
    or g147(n1738 ,n1685 ,n1573);
    or g148(n172 ,n87 ,n134);
    xnor g149(n2709 ,n1233 ,n1257);
    nand g150(n440 ,n258 ,n337);
    nand g151(n456 ,n84 ,n79);
    nand g152(n254 ,n25[3] ,n142);
    xor g153(n812 ,n798 ,n784);
    nand g154(n503 ,n6[4] ,n466);
    not g155(n1645 ,n1644);
    nand g156(n1887 ,n1621 ,n1798);
    nand g157(n389 ,n218 ,n292);
    not g158(n474 ,n475);
    not g159(n1567 ,n21[3]);
    nand g160(n653 ,n546 ,n485);
    nor g161(n53 ,n25[7] ,n52);
    nand g162(n1917 ,n1750 ,n1880);
    nand g163(n2237 ,n2080 ,n2207);
    xor g164(n1265 ,n1263 ,n1427);
    xnor g165(n2016 ,n1843 ,n1694);
    nor g166(n1340 ,n1266 ,n1307);
    or g167(n763 ,n20[2] ,n20[1]);
    nor g168(n2565 ,n2560 ,n2538);
    nand g169(n2317 ,n2259 ,n2282);
    nand g170(n545 ,n20[2] ,n465);
    nor g171(n1399 ,n1312 ,n1349);
    nand g172(n1482 ,n1411 ,n1464);
    dff g173(.RN(n1), .SN(1'b1), .CK(n0), .D(n382), .Q(n17[4]));
    xor g174(n2714 ,n2453 ,n2457);
    nand g175(n1934 ,n1788 ,n1862);
    nand g176(n1617 ,n21[2] ,n23[7]);
    nand g177(n1126 ,n1094 ,n1097);
    xnor g178(n139 ,n19[6] ,n28[6]);
    nand g179(n539 ,n21[0] ,n463);
    xnor g180(n967 ,n806 ,n898);
    buf g181(n12[12], n10[4]);
    nor g182(n1921 ,n1757 ,n1902);
    nand g183(n220 ,n26[8] ,n87);
    nand g184(n1533 ,n1515 ,n1517);
    nor g185(n1767 ,n1701 ,n1615);
    xnor g186(n1907 ,n1658 ,n1809);
    nand g187(n549 ,n19[6] ,n476);
    nand g188(n371 ,n200 ,n273);
    xnor g189(n1837 ,n1599 ,n1590);
    or g190(n2222 ,n2148 ,n2197);
    not g191(n1225 ,n1224);
    nand g192(n334 ,n28[14] ,n141);
    or g193(n1735 ,n1695 ,n1686);
    not g194(n1077 ,n1076);
    nand g195(n400 ,n260 ,n299);
    nor g196(n2584 ,n2534 ,n2560);
    nand g197(n708 ,n575 ,n526);
    nor g198(n1290 ,n1266 ,n1285);
    not g199(n2083 ,n2070);
    xnor g200(n1548 ,n1529 ,n1522);
    nor g201(n1494 ,n1476 ,n1477);
    xnor g202(n1472 ,n1435 ,n1449);
    nor g203(n1345 ,n1269 ,n1304);
    nand g204(n892 ,n2713 ,n846);
    nand g205(n2635 ,n2582 ,n2581);
    buf g206(n11[27], n10[11]);
    dff g207(.RN(n1), .SN(1'b1), .CK(n0), .D(n381), .Q(n28[0]));
    not g208(n1563 ,n1564);
    nand g209(n2337 ,n2311 ,n2321);
    xor g210(n2673 ,n20[1] ,n21[1]);
    buf g211(n9[10], 1'b0);
    nor g212(n1160 ,n1093 ,n1134);
    nand g213(n2115 ,n1927 ,n2043);
    nand g214(n859 ,n2712 ,n825);
    not g215(n1641 ,n1640);
    nand g216(n2427 ,n2426 ,n2412);
    xnor g217(n1438 ,n1391 ,n1394);
    nor g218(n1400 ,n1323 ,n1360);
    nor g219(n115 ,n5[27] ,n5[26]);
    nand g220(n2227 ,n2144 ,n2185);
    xor g221(n2697 ,n969 ,n851);
    nand g222(n2294 ,n2244 ,n2267);
    nand g223(n1594 ,n20[0] ,n22[1]);
    nor g224(n1377 ,n1286 ,n1356);
    dff g225(.RN(n1), .SN(1'b1), .CK(n0), .D(n712), .Q(n21[7]));
    nand g226(n377 ,n205 ,n331);
    nand g227(n194 ,n29[2] ,n87);
    nand g228(n899 ,n799 ,n871);
    nand g229(n1599 ,n20[6] ,n22[5]);
    or g230(n2300 ,n2259 ,n2282);
    nand g231(n45 ,n30[5] ,n44);
    nor g232(n101 ,n5[21] ,n5[20]);
    nand g233(n1490 ,n1452 ,n1468);
    xnor g234(n2099 ,n1993 ,n1928);
    xnor g235(n2717 ,n2463 ,n2451);
    nor g236(n118 ,n26[4] ,n26[5]);
    xnor g237(n2728 ,n2499 ,n2507);
    nor g238(n720 ,n699 ,n696);
    xnor g239(n1858 ,n1707 ,n1719);
    xnor g240(n2305 ,n2250 ,n2192);
    xnor g241(n982 ,n930 ,n932);
    nand g242(n158 ,n102 ,n95);
    nand g243(n2042 ,n1952 ,n1997);
    nand g244(n568 ,n23[4] ,n474);
    or g245(n1463 ,n1429 ,n1448);
    nor g246(n1352 ,n1266 ,n1296);
    buf g247(n13[3], 1'b0);
    buf g248(n11[31], n10[15]);
    nand g249(n1369 ,n1329 ,n1362);
    xnor g250(n2298 ,n2276 ,n2231);
    nand g251(n2359 ,n2305 ,n2344);
    nand g252(n225 ,n26[4] ,n87);
    dff g253(.RN(n1), .SN(1'b1), .CK(n0), .D(n648), .Q(n20[5]));
    nand g254(n2589 ,n2667 ,n2559);
    nand g255(n1686 ,n21[2] ,n23[6]);
    dff g256(.RN(n1), .SN(1'b1), .CK(n0), .D(n665), .Q(n27[1]));
    nor g257(n1100 ,n1043 ,n1081);
    nand g258(n1576 ,n20[5] ,n22[2]);
    xnor g259(n2497 ,n2709 ,n2693);
    nor g260(n1359 ,n1267 ,n1300);
    nand g261(n2637 ,n2579 ,n2608);
    xor g262(n1847 ,n1625 ,n1591);
    buf g263(n11[30], n10[14]);
    nand g264(n564 ,n24[0] ,n461);
    not g265(n2491 ,n2490);
    nand g266(n2611 ,n2703 ,n2547);
    nor g267(n2482 ,n2704 ,n2688);
    buf g268(n12[7], 1'b0);
    nor g269(n1935 ,n1743 ,n1881);
    xnor g270(n2230 ,n2126 ,n2132);
    nand g271(n898 ,n794 ,n855);
    nor g272(n1416 ,n1386 ,n1380);
    nor g273(n1326 ,n1267 ,n1278);
    xnor g274(n1221 ,n1198 ,n1190);
    nand g275(n1557 ,n1542 ,n1556);
    xnor g276(n2485 ,n2704 ,n2688);
    dff g277(.RN(n1), .SN(1'b1), .CK(n0), .D(n423), .Q(n10[7]));
    nand g278(n2662 ,n2599 ,n2648);
    nand g279(n2094 ,n1972 ,n2049);
    nor g280(n2438 ,n22[7] ,n23[7]);
    not g281(n1984 ,n1983);
    nand g282(n358 ,n285 ,n178);
    buf g283(n13[6], 1'b0);
    xnor g284(n1001 ,n930 ,n928);
    nand g285(n1281 ,n2674 ,n23[2]);
    xnor g286(n2144 ,n2029 ,n1952);
    not g287(n1855 ,n1854);
    nor g288(n1176 ,n1121 ,n1145);
    nand g289(n2097 ,n1971 ,n2050);
    nand g290(n911 ,n2715 ,n876);
    nor g291(n1177 ,n1101 ,n1159);
    nand g292(n881 ,n2713 ,n848);
    nand g293(n2007 ,n1929 ,n1908);
    nand g294(n2152 ,n1979 ,n1565);
    nor g295(n1253 ,n1237 ,n1252);
    nand g296(n1676 ,n20[2] ,n22[5]);
    nand g297(n213 ,n26[15] ,n140);
    nand g298(n1496 ,n1428 ,n1470);
    or g299(n765 ,n20[6] ,n20[5]);
    nand g300(n335 ,n29[9] ,n141);
    xnor g301(n2131 ,n2028 ,n1965);
    xnor g302(n1987 ,n1837 ,n1713);
    nand g303(n1300 ,n1285 ,n1272);
    nand g304(n689 ,n562 ,n517);
    xnor g305(n1974 ,n1839 ,n1655);
    nand g306(n1784 ,n1684 ,n1606);
    nor g307(n718 ,n680 ,n679);
    nand g308(n591 ,n19[7] ,n481);
    nand g309(n905 ,n789 ,n860);
    nor g310(n1105 ,n1045 ,n1082);
    xnor g311(n1485 ,n1458 ,n1459);
    nand g312(n2153 ,n2119 ,n2052);
    nor g313(n1394 ,n1313 ,n1343);
    nand g314(n418 ,n317 ,n237);
    nand g315(n1127 ,n1089 ,n1094);
    nor g316(n1195 ,n1103 ,n1172);
    nor g317(n1240 ,n1210 ,n1226);
    nand g318(n401 ,n226 ,n300);
    not g319(n461 ,n462);
    buf g320(n9[31], 1'b0);
    nor g321(n446 ,n185 ,n383);
    dff g322(.RN(n1), .SN(1'b1), .CK(n0), .D(n352), .Q(n29[5]));
    nand g323(n871 ,n2719 ,n825);
    dff g324(.RN(n1), .SN(1'b1), .CK(n0), .D(n735), .Q(n9[3]));
    nor g325(n1479 ,n1453 ,n1456);
    nand g326(n872 ,n2719 ,n824);
    nand g327(n1874 ,n1646 ,n1776);
    nor g328(n475 ,n344 ,n460);
    nand g329(n1908 ,n1763 ,n1858);
    nor g330(n1051 ,n987 ,n985);
    or g331(n2356 ,n2318 ,n2345);
    nand g332(n1588 ,n20[4] ,n22[4]);
    nand g333(n946 ,n862 ,n895);
    nand g334(n151 ,n113 ,n106);
    xnor g335(n1224 ,n1183 ,n1136);
    nand g336(n1697 ,n20[3] ,n22[5]);
    xnor g337(n1440 ,n1396 ,n1326);
    dff g338(.RN(n1), .SN(1'b1), .CK(n0), .D(n705), .Q(n22[7]));
    buf g339(n12[2], 1'b0);
    nand g340(n1597 ,n20[1] ,n22[2]);
    nand g341(n1794 ,n1697 ,n1575);
    buf g342(n13[25], n10[1]);
    nand g343(n2416 ,n2396 ,n1566);
    dff g344(.RN(n1), .SN(1'b1), .CK(n0), .D(n652), .Q(n20[2]));
    nand g345(n1483 ,n1406 ,n1463);
    nand g346(n1423 ,n1390 ,n1374);
    nand g347(n2400 ,n2361 ,n2390);
    not g348(n1614 ,n1613);
    nand g349(n2658 ,n2614 ,n2636);
    nor g350(n1442 ,n1427 ,n1263);
    nand g351(n639 ,n533 ,n495);
    nand g352(n2479 ,n2710 ,n2694);
    nor g353(n1335 ,n1266 ,n1303);
    dff g354(.RN(n1), .SN(1'b1), .CK(n0), .D(n708), .Q(n22[5]));
    or g355(n2041 ,n1969 ,n1967);
    nand g356(n629 ,n20[1] ,n468);
    xnor g357(n32[5] ,n1538 ,n1546);
    dff g358(.RN(n1), .SN(1'b1), .CK(n0), .D(n435), .Q(n29[14]));
    xor g359(n1026 ,n931 ,n970);
    nand g360(n2597 ,n2668 ,n2559);
    xor g361(n813 ,n797 ,n775);
    nand g362(n1952 ,n1747 ,n1876);
    dff g363(.RN(n1), .SN(1'b1), .CK(n0), .D(n656), .Q(n19[7]));
    nand g364(n1791 ,n1580 ,n1680);
    nand g365(n659 ,n551 ,n509);
    dff g366(.RN(n1), .SN(1'b1), .CK(n0), .D(n731), .Q(n9[7]));
    xnor g367(n2689 ,n2420 ,n2424);
    xnor g368(n773 ,n20[1] ,n21[1]);
    nor g369(n123 ,n89 ,n5[3]);
    nand g370(n699 ,n626 ,n625);
    nand g371(n882 ,n2716 ,n848);
    nand g372(n419 ,n318 ,n238);
    nand g373(n505 ,n6[2] ,n466);
    or g374(n1543 ,n1523 ,n1530);
    nand g375(n2349 ,n2291 ,n2332);
    buf g376(n12[21], n10[13]);
    xor g377(n757 ,n981 ,n971);
    dff g378(.RN(n1), .SN(1'b1), .CK(n0), .D(n406), .Q(n25[7]));
    nand g379(n1867 ,n1659 ,n1809);
    nand g380(n138 ,n90 ,n108);
    nand g381(n2264 ,n2192 ,n2226);
    nand g382(n1500 ,n1409 ,n1480);
    xnor g383(n2492 ,n2697 ,n2681);
    nand g384(n1575 ,n21[5] ,n23[3]);
    nand g385(n442 ,n221 ,n295);
    dff g386(.RN(n1), .SN(1'b1), .CK(n0), .D(n349), .Q(n26[8]));
    nand g387(n2643 ,n2622 ,n2591);
    nor g388(n1005 ,n849 ,n963);
    nand g389(n1793 ,n1655 ,n1604);
    nand g390(n2361 ,n2318 ,n2345);
    nor g391(n1102 ,n1090 ,n1062);
    xnor g392(n1064 ,n985 ,n987);
    nand g393(n604 ,n19[5] ,n481);
    nand g394(n887 ,n2717 ,n846);
    dff g395(.RN(n1), .SN(1'b1), .CK(n0), .D(n736), .Q(n9[0]));
    nand g396(n1656 ,n21[7] ,n23[6]);
    nand g397(n530 ,n6[7] ,n464);
    nand g398(n2293 ,n2227 ,n2264);
    nand g399(n514 ,n6[5] ,n462);
    nand g400(n1705 ,n21[3] ,n23[5]);
    nand g401(n63 ,n30[5] ,n61);
    nor g402(n851 ,n807 ,n823);
    nand g403(n544 ,n20[3] ,n465);
    xnor g404(n1191 ,n1095 ,n1140);
    nand g405(n2608 ,n2709 ,n2547);
    xnor g406(n778 ,n20[6] ,n21[6]);
    nand g407(n1692 ,n20[3] ,n22[3]);
    nand g408(n2575 ,n32[10] ,n2561);
    nand g409(n245 ,n31[3] ,n155);
    xnor g410(n1439 ,n1392 ,n1308);
    nand g411(n1999 ,n1852 ,n1948);
    nand g412(n1608 ,n21[1] ,n23[7]);
    nand g413(n2548 ,n2725 ,n32[8]);
    nand g414(n2460 ,n2455 ,n2459);
    not g415(n2081 ,n2065);
    or g416(n2413 ,n2393 ,n2404);
    nand g417(n1552 ,n1533 ,n1551);
    nor g418(n2471 ,n2699 ,n2683);
    nor g419(n2522 ,n2501 ,n2521);
    nand g420(n2255 ,n2149 ,n2236);
    nand g421(n518 ,n6[7] ,n475);
    buf g422(n13[19], 1'b0);
    buf g423(n13[4], 1'b0);
    xnor g424(n2249 ,n2212 ,n2188);
    xnor g425(n2706 ,n1242 ,n1251);
    nand g426(n605 ,n22[4] ,n469);
    xnor g427(n1827 ,n1588 ,n1601);
    xnor g428(n2411 ,n2398 ,n2381);
    nor g429(n2536 ,n2724 ,n32[9]);
    nand g430(n546 ,n20[1] ,n465);
    nand g431(n1883 ,n1618 ,n1781);
    buf g432(n11[11], 1'b0);
    dff g433(.RN(n1), .SN(1'b1), .CK(n0), .D(n692), .Q(n24[0]));
    not g434(n1311 ,n1310);
    nand g435(n2630 ,n2557 ,n2566);
    buf g436(n9[25], 1'b0);
    nand g437(n390 ,n219 ,n293);
    nand g438(n525 ,n6[6] ,n479);
    nor g439(n1291 ,n1269 ,n1281);
    xnor g440(n32[2] ,n1467 ,n1426);
    or g441(n31[0] ,n2634 ,n2654);
    nor g442(n42 ,n30[2] ,n30[0]);
    nand g443(n146 ,n122 ,n86);
    dff g444(.RN(n1), .SN(1'b1), .CK(n0), .D(n738), .Q(n9[2]));
    or g445(n2257 ,n2157 ,n2230);
    nand g446(n880 ,n2715 ,n847);
    nor g447(n1396 ,n1290 ,n1359);
    or g448(n1747 ,n1687 ,n1591);
    nand g449(n2386 ,n2292 ,n2357);
    not g450(n787 ,n21[0]);
    dff g451(.RN(n1), .SN(1'b1), .CK(n0), .D(n682), .Q(n24[7]));
    xnor g452(n811 ,n787 ,n773);
    not g453(n128 ,n127);
    nor g454(n1870 ,n1586 ,n1765);
    xnor g455(n1830 ,n1682 ,n1579);
    nand g456(n1605 ,n20[1] ,n22[5]);
    nand g457(n1571 ,n21[5] ,n23[2]);
    xor g458(n2679 ,n20[7] ,n21[7]);
    buf g459(n12[9], n10[1]);
    nand g460(n357 ,n194 ,n175);
    nand g461(n1879 ,n1624 ,n1771);
    or g462(n31[6] ,n2628 ,n2655);
    nor g463(n1902 ,n1648 ,n1812);
    nand g464(n290 ,n29[13] ,n141);
    not g465(n478 ,n479);
    dff g466(.RN(n1), .SN(1'b1), .CK(n0), .D(n711), .Q(n22[2]));
    dff g467(.RN(n1), .SN(1'b1), .CK(n0), .D(n433), .Q(n29[15]));
    xnor g468(n2090 ,n1970 ,n1973);
    nand g469(n1367 ,n24[0] ,n1306);
    nor g470(n97 ,n26[1] ,n26[2]);
    or g471(n1245 ,n1208 ,n1244);
    xnor g472(n1969 ,n1820 ,n1702);
    nand g473(n733 ,n725 ,n716);
    buf g474(n13[31], n10[7]);
    nand g475(n2177 ,n2141 ,n2130);
    not g476(n1609 ,n1608);
    or g477(n2328 ,n2260 ,n2303);
    xnor g478(n2143 ,n2024 ,n1926);
    nand g479(n833 ,n2714 ,n819);
    nand g480(n1296 ,n1282 ,n1273);
    nand g481(n1906 ,n1627 ,n1793);
    xnor g482(n968 ,n817 ,n908);
    not g483(n934 ,n933);
    nand g484(n2507 ,n2481 ,n2506);
    nand g485(n666 ,n587 ,n586);
    nand g486(n2390 ,n2329 ,n2373);
    nand g487(n2287 ,n2128 ,n2274);
    nand g488(n651 ,n585 ,n584);
    xnor g489(n131 ,n19[5] ,n28[5]);
    dff g490(.RN(n1), .SN(1'b1), .CK(n0), .D(n384), .Q(n17[3]));
    nand g491(n1542 ,n1522 ,n1529);
    nor g492(n1390 ,n1324 ,n1358);
    nand g493(n224 ,n26[5] ,n87);
    dff g494(.RN(n1), .SN(1'b1), .CK(n0), .D(n663), .Q(n19[0]));
    not g495(n2532 ,n27[1]);
    dff g496(.RN(n1), .SN(1'b1), .CK(n0), .D(n430), .Q(n10[1]));
    xnor g497(n1015 ,n817 ,n954);
    or g498(n1736 ,n1660 ,n1592);
    xnor g499(n2344 ,n2299 ,n2283);
    nor g500(n1766 ,n1707 ,n1719);
    nand g501(n1632 ,n21[6] ,n23[1]);
    nor g502(n1382 ,n1319 ,n1354);
    xnor g503(n2684 ,n2326 ,n2294);
    nand g504(n943 ,n836 ,n896);
    dff g505(.RN(n1), .SN(1'b1), .CK(n0), .D(n365), .Q(n28[10]));
    nand g506(n941 ,n831 ,n879);
    nand g507(n2620 ,n2711 ,n2547);
    nor g508(n2515 ,n2472 ,n2514);
    nand g509(n623 ,n24[1] ,n482);
    nand g510(n1408 ,n1348 ,n1383);
    nand g511(n2236 ,n2163 ,n2181);
    or g512(n764 ,n20[4] ,n20[3]);
    nand g513(n1876 ,n1625 ,n1799);
    nand g514(n1639 ,n21[3] ,n23[6]);
    or g515(n2506 ,n2496 ,n2505);
    nand g516(n928 ,n837 ,n910);
    xnor g517(n2499 ,n2699 ,n2683);
    nand g518(n953 ,n865 ,n883);
    not g519(n2495 ,n2494);
    xnor g520(n1964 ,n1846 ,n1676);
    nor g521(n1356 ,n1267 ,n1296);
    not g522(n1714 ,n1713);
    nor g523(n1877 ,n1639 ,n1811);
    nor g524(n1342 ,n1267 ,n1305);
    not g525(n2653 ,n2644);
    nand g526(n2646 ,n2554 ,n2569);
    nor g527(n1405 ,n1395 ,n1372);
    not g528(n57 ,n56);
    xnor g529(n2722 ,n2487 ,n2519);
    nand g530(n2554 ,n2722 ,n32[11]);
    not g531(n1199 ,n1198);
    nor g532(n1726 ,n1602 ,n1653);
    nand g533(n590 ,n20[7] ,n468);
    nand g534(n2068 ,n2014 ,n2016);
    or g535(n175 ,n87 ,n137);
    nand g536(n2008 ,n1871 ,n1923);
    xnor g537(n817 ,n800 ,n785);
    nor g538(n114 ,n5[13] ,n5[12]);
    dff g539(.RN(n1), .SN(1'b1), .CK(n0), .D(n646), .Q(n20[7]));
    nand g540(n2010 ,n1784 ,n1957);
    nand g541(n2621 ,n2700 ,n2547);
    nand g542(n569 ,n23[3] ,n474);
    nand g543(n77 ,n25[6] ,n76);
    nor g544(n2541 ,n2729 ,n32[4]);
    xnor g545(n2724 ,n2486 ,n2515);
    nand g546(n1939 ,n1735 ,n1899);
    xnor g547(n1013 ,n955 ,n817);
    not g548(n1094 ,n1095);
    nor g549(n1320 ,n1269 ,n1283);
    nand g550(n2650 ,n2603 ,n2601);
    nand g551(n1950 ,n1758 ,n1900);
    nand g552(n2632 ,n2549 ,n2564);
    nand g553(n838 ,n2717 ,n819);
    nand g554(n264 ,n30[4] ,n87);
    nand g555(n207 ,n28[2] ,n87);
    nand g556(n1604 ,n21[7] ,n23[4]);
    nor g557(n1343 ,n1269 ,n1300);
    nor g558(n1213 ,n1199 ,n1190);
    nand g559(n2366 ,n2304 ,n2350);
    buf g560(n12[28], 1'b0);
    xnor g561(n1517 ,n1485 ,n1472);
    not g562(n1430 ,n1422);
    nand g563(n522 ,n6[3] ,n475);
    not g564(n1709 ,n1708);
    nand g565(n1209 ,n1181 ,n1187);
    xnor g566(n1228 ,n1180 ,n1187);
    nand g567(n2263 ,n2157 ,n2230);
    not g568(n2082 ,n2067);
    xnor g569(n2015 ,n1835 ,n1767);
    nand g570(n380 ,n210 ,n283);
    nand g571(n1535 ,n1520 ,n1524);
    xnor g572(n1966 ,n1842 ,n1711);
    nand g573(n1629 ,n21[0] ,n23[5]);
    nand g574(n2275 ,n2202 ,n2222);
    buf g575(n13[12], 1'b0);
    nand g576(n263 ,n30[3] ,n87);
    nor g577(n1426 ,n1348 ,n1383);
    nand g578(n1215 ,n1179 ,n1193);
    nand g579(n1200 ,n1143 ,n1167);
    nand g580(n1725 ,n20[0] ,n22[0]);
    or g581(n1754 ,n1675 ,n1668);
    dff g582(.RN(n1), .SN(1'b1), .CK(n0), .D(n368), .Q(n28[15]));
    nor g583(n2569 ,n2560 ,n2545);
    nor g584(n1078 ,n998 ,n1028);
    nor g585(n1627 ,n1569 ,n1568);
    xnor g586(n2017 ,n1833 ,n1720);
    nand g587(n136 ,n124 ,n85);
    not g588(n2136 ,n2135);
    nand g589(n2002 ,n1915 ,n1916);
    xnor g590(n1121 ,n1073 ,n989);
    xor g591(n756 ,n979 ,n967);
    not g592(n1700 ,n1699);
    nand g593(n392 ,n256 ,n335);
    nor g594(n1058 ,n980 ,n1019);
    nand g595(n241 ,n31[6] ,n155);
    not g596(n90 ,n2);
    not g597(n1364 ,n1363);
    xnor g598(n2715 ,n2454 ,n2459);
    not g599(n1190 ,n1189);
    nand g600(n1280 ,n2673 ,n23[1]);
    nand g601(n1869 ,n1667 ,n1766);
    nor g602(n2439 ,n22[6] ,n23[6]);
    buf g603(n12[20], n10[12]);
    nand g604(n1109 ,n1048 ,n1085);
    nor g605(n2468 ,n2448 ,n2467);
    nand g606(n1279 ,n2676 ,n23[4]);
    nand g607(n1803 ,n1602 ,n1653);
    nor g608(n1313 ,n1268 ,n1285);
    nand g609(n196 ,n31[5] ,n155);
    nand g610(n799 ,n2720 ,n783);
    nand g611(n2383 ,n2363 ,n2368);
    buf g612(n9[14], 1'b0);
    xnor g613(n1222 ,n1193 ,n1179);
    nand g614(n1704 ,n20[7] ,n22[0]);
    dff g615(.RN(n1), .SN(1'b1), .CK(n0), .D(n357), .Q(n29[2]));
    nor g616(n1378 ,n1316 ,n1339);
    nand g617(n555 ,n27[1] ,n471);
    xnor g618(n1826 ,n1695 ,n1686);
    nand g619(n2244 ,n2078 ,n2191);
    nand g620(n648 ,n542 ,n502);
    buf g621(n12[6], 1'b0);
    or g622(n2367 ,n2302 ,n2351);
    xnor g623(n2125 ,n2015 ,n2047);
    nor g624(n1088 ,n1017 ,n1027);
    nand g625(n2201 ,n2048 ,n2134);
    dff g626(.RN(n1), .SN(1'b1), .CK(n0), .D(n375), .Q(n28[6]));
    nand g627(n1949 ,n1756 ,n1898);
    nand g628(n2001 ,n1853 ,n1947);
    nand g629(n1154 ,n1096 ,n1117);
    nor g630(n1218 ,n1198 ,n1189);
    nand g631(n559 ,n24[5] ,n461);
    nand g632(n921 ,n832 ,n878);
    xnor g633(n1402 ,n1365 ,n1310);
    not g634(n1812 ,n1782);
    nand g635(n2037 ,n1922 ,n1998);
    dff g636(.RN(n1), .SN(1'b1), .CK(n0), .D(n431), .Q(n10[0]));
    nand g637(n2586 ,n2666 ,n2561);
    not g638(n2450 ,n2449);
    nand g639(n1658 ,n21[6] ,n23[4]);
    nor g640(n445 ,n26[3] ,n348);
    nand g641(n1555 ,n1545 ,n1554);
    nand g642(n707 ,n574 ,n525);
    nand g643(n1927 ,n1741 ,n1888);
    nand g644(n2617 ,n2698 ,n2547);
    nand g645(n609 ,n20[4] ,n468);
    not g646(n1182 ,n1178);
    nand g647(n372 ,n222 ,n267);
    nand g648(n2070 ,n2013 ,n2017);
    dff g649(.RN(n1), .SN(1'b1), .CK(n0), .D(n694), .Q(n23[6]));
    xnor g650(n1865 ,n1660 ,n1623);
    nand g651(n1936 ,n1751 ,n1885);
    or g652(n1406 ,n1373 ,n1375);
    nand g653(n2067 ,n1973 ,n1970);
    not g654(n1414 ,n1408);
    or g655(n2415 ,n2397 ,n2403);
    nand g656(n233 ,n31[15] ,n155);
    not g657(n92 ,n18[2]);
    dff g658(.RN(n1), .SN(1'b1), .CK(n0), .D(n698), .Q(n23[3]));
    or g659(n31[1] ,n2652 ,n2658);
    nand g660(n2292 ,n2243 ,n2255);
    dff g661(.RN(n1), .SN(1'b1), .CK(n0), .D(n650), .Q(n20[3]));
    xnor g662(n2173 ,n2021 ,n2099);
    nand g663(n626 ,n19[1] ,n481);
    nand g664(n297 ,n753 ,n141);
    xnor g665(n1958 ,n1863 ,n1666);
    buf g666(n12[16], n10[8]);
    dff g667(.RN(n1), .SN(1'b1), .CK(n0), .D(n392), .Q(n26[9]));
    nand g668(n1084 ,n970 ,n1054);
    xnor g669(n1959 ,n1860 ,n1691);
    or g670(n1480 ,n1417 ,n1460);
    not g671(n2130 ,n2129);
    dff g672(.RN(n1), .SN(1'b1), .CK(n0), .D(n709), .Q(n22[4]));
    dff g673(.RN(n1), .SN(1'b1), .CK(n0), .D(n707), .Q(n22[6]));
    xnor g674(n2325 ,n2258 ,n2282);
    nand g675(n1484 ,n1425 ,n1466);
    nand g676(n630 ,n23[0] ,n480);
    nand g677(n2116 ,n2019 ,n2068);
    nand g678(n211 ,n31[9] ,n155);
    not g679(n1299 ,n1300);
    nor g680(n1053 ,n933 ,n1014);
    nand g681(n884 ,n2714 ,n848);
    nand g682(n2392 ,n2349 ,n2382);
    nand g683(n1202 ,n1128 ,n1175);
    nand g684(n1590 ,n20[7] ,n22[4]);
    xnor g685(n2696 ,n806 ,n823);
    nor g686(n2469 ,n2703 ,n2687);
    xnor g687(n1993 ,n1856 ,n1807);
    nor g688(n1338 ,n1269 ,n1307);
    nand g689(n1699 ,n21[5] ,n23[7]);
    buf g690(n10[22], 1'b0);
    or g691(n2176 ,n1962 ,n2146);
    nand g692(n2178 ,n2142 ,n2129);
    nand g693(n2313 ,n2269 ,n2283);
    nand g694(n2588 ,n2695 ,n2546);
    or g695(n1410 ,n1384 ,n1382);
    dff g696(.RN(n1), .SN(1'b1), .CK(n0), .D(n639), .Q(n21[6]));
    nor g697(n1216 ,n1202 ,n1192);
    buf g698(n10[31], 1'b0);
    or g699(n1749 ,n1607 ,n1578);
    buf g700(n11[24], n10[8]);
    nand g701(n581 ,n21[7] ,n463);
    or g702(n1728 ,n1672 ,n1577);
    nand g703(n1130 ,n977 ,n1111);
    nand g704(n2273 ,n2200 ,n2228);
    or g705(n2309 ,n2269 ,n2283);
    dff g706(.RN(n1), .SN(1'b1), .CK(n0), .D(n415), .Q(n10[14]));
    or g707(n1499 ,n1428 ,n1470);
    nand g708(n223 ,n26[6] ,n87);
    nand g709(n425 ,n324 ,n196);
    xor g710(n1263 ,n1346 ,n1333);
    or g711(n1143 ,n1075 ,n1120);
    xnor g712(n984 ,n942 ,n816);
    nand g713(n1522 ,n1491 ,n1506);
    not g714(n806 ,n807);
    nand g715(n1087 ,n968 ,n1046);
    not g716(n1862 ,n1861);
    dff g717(.RN(n1), .SN(1'b1), .CK(n0), .D(n380), .Q(n28[1]));
    nand g718(n449 ,n97 ,n445);
    nand g719(n2399 ,n2362 ,n2389);
    nor g720(n1134 ,n1107 ,n1092);
    xnor g721(n2681 ,n1761 ,n2086);
    not g722(n1473 ,n1472);
    nand g723(n2574 ,n2685 ,n2546);
    or g724(n2209 ,n2099 ,n2133);
    nand g725(n192 ,n28[10] ,n87);
    xnor g726(n2304 ,n2249 ,n2273);
    xnor g727(n935 ,n852 ,n807);
    nand g728(n2372 ,n2319 ,n2347);
    nand g729(n1771 ,n1660 ,n1592);
    nand g730(n1592 ,n20[2] ,n22[2]);
    nand g731(n554 ,n19[1] ,n476);
    nand g732(n664 ,n557 ,n532);
    not g733(n1657 ,n1656);
    buf g734(n9[29], 1'b0);
    nand g735(n193 ,n29[14] ,n140);
    nand g736(n1786 ,n1588 ,n1601);
    nand g737(n556 ,n19[0] ,n476);
    nand g738(n1593 ,n21[3] ,n23[0]);
    nor g739(n2195 ,n2120 ,n2158);
    or g740(n179 ,n158 ,n159);
    or g741(n1734 ,n1670 ,n1674);
    nor g742(n1012 ,n971 ,n981);
    nand g743(n582 ,n27[0] ,n472);
    nand g744(n2644 ,n2598 ,n2594);
    nand g745(n940 ,n833 ,n886);
    xnor g746(n32[9] ,n1549 ,n1557);
    dff g747(.RN(n1), .SN(1'b1), .CK(n0), .D(n400), .Q(n26[3]));
    nor g748(n1308 ,n1267 ,n1284);
    xnor g749(n2084 ,n1961 ,n1968);
    nand g750(n1801 ,n1689 ,n1654);
    nand g751(n1885 ,n1796 ,n1767);
    nand g752(n2053 ,n1753 ,n2000);
    buf g753(n12[4], 1'b0);
    nand g754(n875 ,n21[7] ,n822);
    nand g755(n519 ,n6[6] ,n475);
    nand g756(n2353 ,n2317 ,n2338);
    nand g757(n1889 ,n1723 ,n1786);
    nor g758(n1194 ,n1104 ,n1171);
    xnor g759(n2364 ,n2325 ,n2293);
    nand g760(n78 ,n161 ,n81);
    nand g761(n640 ,n534 ,n496);
    nand g762(n535 ,n21[4] ,n463);
    or g763(n2062 ,n2013 ,n2017);
    nor g764(n2278 ,n2270 ,n2261);
    or g765(n1347 ,n1268 ,n1301);
    nor g766(n83 ,n146 ,n158);
    nand g767(n683 ,n595 ,n513);
    xnor g768(n803 ,n762 ,n776);
    nand g769(n1544 ,n1519 ,n1528);
    nand g770(n2524 ,n2495 ,n2523);
    nand g771(n2580 ,n2680 ,n2546);
    nand g772(n489 ,n6[1] ,n462);
    xnor g773(n957 ,n818 ,n904);
    nand g774(n768 ,n20[2] ,n20[1]);
    not g775(n1022 ,n1021);
    nor g776(n482 ,n252 ,n458);
    nand g777(n301 ,n29[3] ,n87);
    nand g778(n349 ,n220 ,n294);
    buf g779(n10[26], 1'b0);
    or g780(n2210 ,n1966 ,n2132);
    nor g781(n2665 ,n1268 ,n1296);
    nor g782(n2393 ,n2375 ,n2385);
    or g783(n1746 ,n1597 ,n1669);
    nand g784(n2612 ,n2707 ,n2547);
    nand g785(n1711 ,n21[7] ,n23[5]);
    nand g786(n1675 ,n20[2] ,n22[3]);
    buf g787(n9[18], 1'b0);
    xnor g788(n1468 ,n1433 ,n1448);
    not g789(n1332 ,n1331);
    nand g790(n1298 ,n1278 ,n1275);
    nand g791(n1892 ,n1709 ,n1790);
    xor g792(n2297 ,n2260 ,n2275);
    or g793(n1732 ,n1598 ,n1593);
    xnor g794(n2685 ,n2340 ,n2355);
    nor g795(n1350 ,n1269 ,n1301);
    nor g796(n2066 ,n1936 ,n1986);
    nand g797(n1802 ,n1676 ,n1576);
    nand g798(n374 ,n265 ,n279);
    nand g799(n156 ,n18[2] ,n119);
    nor g800(n1368 ,n1328 ,n1363);
    nand g801(n863 ,n2718 ,n824);
    not g802(n1040 ,n1034);
    nand g803(n2149 ,n2040 ,n2098);
    nor g804(n1287 ,n1268 ,n1278);
    nand g805(n867 ,n2715 ,n824);
    xnor g806(n1549 ,n1530 ,n1523);
    not g807(n2145 ,n2144);
    xnor g808(n1538 ,n1514 ,n1516);
    nand g809(n70 ,n25[2] ,n69);
    not g810(n758 ,n2717);
    buf g811(n10[21], 1'b0);
    nand g812(n680 ,n614 ,n613);
    xor g813(n819 ,n805 ,n809);
    nand g814(n916 ,n2719 ,n848);
    nor g815(n481 ,n252 ,n457);
    dff g816(.RN(n1), .SN(1'b1), .CK(n0), .D(n425), .Q(n10[5]));
    xnor g817(n991 ,n816 ,n922);
    nand g818(n1655 ,n20[5] ,n22[6]);
    xnor g819(n2028 ,n1924 ,n1917);
    nand g820(n1642 ,n21[0] ,n23[2]);
    dff g821(.RN(n1), .SN(1'b1), .CK(n0), .D(n701), .Q(n23[1]));
    xnor g822(n1184 ,n1113 ,n1146);
    nand g823(n904 ,n2720 ,n848);
    xnor g824(n1071 ,n1008 ,n966);
    nand g825(n2147 ,n2036 ,n2114);
    dff g826(.RN(n1), .SN(1'b1), .CK(n0), .D(n683), .Q(n24[6]));
    nor g827(n725 ,n635 ,n674);
    xnor g828(n2013 ,n1865 ,n1592);
    nor g829(n1740 ,n1580 ,n1680);
    nor g830(n1349 ,n1266 ,n1300);
    nand g831(n2613 ,n2696 ,n2547);
    nand g832(n361 ,n257 ,n269);
    not g833(n2101 ,n2100);
    nand g834(n1925 ,n1734 ,n1883);
    nand g835(n2354 ,n2310 ,n2335);
    nand g836(n2398 ,n2358 ,n2386);
    nand g837(n50 ,n48 ,n47);
    nand g838(n1582 ,n20[6] ,n22[7]);
    nand g839(n2664 ,n2615 ,n2630);
    nor g840(n1427 ,n1367 ,n1377);
    nand g841(n1796 ,n1584 ,n1677);
    dff g842(.RN(n1), .SN(1'b1), .CK(n0), .D(n399), .Q(n26[4]));
    nand g843(n260 ,n26[3] ,n87);
    nand g844(n1478 ,n1426 ,n1462);
    not g845(n1059 ,n1058);
    nand g846(n1651 ,n20[7] ,n22[6]);
    nand g847(n186 ,n126 ,n142);
    nand g848(n1578 ,n20[7] ,n22[3]);
    nand g849(n2603 ,n2689 ,n2546);
    buf g850(n13[18], 1'b0);
    nand g851(n2321 ,n2263 ,n2289);
    nand g852(n533 ,n21[6] ,n463);
    dff g853(.RN(n1), .SN(1'b1), .CK(n0), .D(n386), .Q(n26[14]));
    nand g854(n204 ,n28[6] ,n87);
    nand g855(n972 ,n815 ,n937);
    dff g856(.RN(n1), .SN(1'b1), .CK(n0), .D(n647), .Q(n20[6]));
    or g857(n98 ,n5[1] ,n5[0]);
    nand g858(n281 ,n31[5] ,n141);
    nand g859(n2615 ,n2704 ,n2547);
    nor g860(n144 ,n18[2] ,n117);
    nand g861(n2064 ,n1988 ,n1976);
    nand g862(n577 ,n22[3] ,n478);
    nand g863(n606 ,n21[4] ,n467);
    nand g864(n243 ,n31[4] ,n155);
    nor g865(n1310 ,n1267 ,n1280);
    xnor g866(n2229 ,n2125 ,n2165);
    nand g867(n2073 ,n1954 ,n2009);
    or g868(n2414 ,n2396 ,n1566);
    buf g869(n13[8], 1'b0);
    nor g870(n452 ,n186 ,n444);
    nand g871(n405 ,n229 ,n303);
    nand g872(n1278 ,n2678 ,n23[6]);
    nand g873(n952 ,n866 ,n891);
    nand g874(n831 ,n2718 ,n820);
    nor g875(n33 ,n30[1] ,n30[0]);
    nand g876(n1694 ,n21[7] ,n23[3]);
    nand g877(n2642 ,n2592 ,n2617);
    xnor g878(n2104 ,n1995 ,n1929);
    nor g879(n2519 ,n2482 ,n2518);
    nor g880(n1354 ,n1267 ,n1304);
    nor g881(n2233 ,n2159 ,n2189);
    or g882(n2265 ,n2183 ,n2229);
    nor g883(n469 ,n252 ,n455);
    xnor g884(n1205 ,n1171 ,n1103);
    nor g885(n86 ,n5[7] ,n5[6]);
    nor g886(n1162 ,n973 ,n1131);
    xnor g887(n2716 ,n2461 ,n2445);
    or g888(n1752 ,n1676 ,n1576);
    nand g889(n781 ,n21[2] ,n763);
    nand g890(n853 ,n2712 ,n824);
    xnor g891(n1451 ,n1401 ,n1382);
    nor g892(n726 ,n636 ,n677);
    nand g893(n2270 ,n2180 ,n2232);
    dff g894(.RN(n1), .SN(1'b1), .CK(n0), .D(n407), .Q(n25[6]));
    nand g895(n1304 ,n1279 ,n1274);
    not g896(n1309 ,n1308);
    nand g897(n365 ,n192 ,n276);
    nand g898(n2599 ,n2684 ,n2546);
    nor g899(n1260 ,n1259 ,n1229);
    xnor g900(n1185 ,n1150 ,n1121);
    nor g901(n161 ,n116 ,n98);
    nor g902(n1295 ,n1269 ,n1282);
    nand g903(n1301 ,n1281 ,n1277);
    nand g904(n352 ,n261 ,n167);
    buf g905(n9[12], 1'b0);
    nand g906(n691 ,n434 ,n620);
    nand g907(n311 ,n750 ,n141);
    nand g908(n2616 ,n2708 ,n2547);
    nor g909(n1337 ,n1267 ,n1298);
    or g910(n1755 ,n1582 ,n1651);
    xnor g911(n1819 ,n1607 ,n1578);
    nor g912(n1807 ,n1619 ,n1616);
    xnor g913(n939 ,n818 ,n826);
    dff g914(.RN(n1), .SN(1'b1), .CK(n0), .D(n416), .Q(n10[13]));
    xor g915(n814 ,n796 ,n785);
    nor g916(n1894 ,n1629 ,n1813);
    not g917(n2185 ,n2184);
    nand g918(n948 ,n870 ,n916);
    nand g919(n658 ,n550 ,n508);
    nand g920(n596 ,n20[6] ,n468);
    xnor g921(n2362 ,n2324 ,n2321);
    nand g922(n72 ,n25[3] ,n71);
    nand g923(n2159 ,n2062 ,n2113);
    nand g924(n325 ,n10[4] ,n156);
    or g925(n1498 ,n1413 ,n1474);
    nand g926(n228 ,n28[15] ,n140);
    xor g927(n2712 ,n23[0] ,n22[0]);
    nand g928(n404 ,n9[6] ,n252);
    nand g929(n566 ,n23[6] ,n474);
    nand g930(n2212 ,n2074 ,n2151);
    nand g931(n677 ,n421 ,n609);
    buf g932(n12[0], 1'b0);
    not g933(n2259 ,n2258);
    or g934(n1727 ,n1574 ,n1683);
    xnor g935(n805 ,n766 ,n777);
    nand g936(n1589 ,n20[3] ,n22[6]);
    nand g937(n276 ,n31[10] ,n141);
    nand g938(n1258 ,n1230 ,n1257);
    nor g939(n751 ,n62 ,n64);
    nand g940(n650 ,n544 ,n504);
    xnor g941(n1476 ,n1436 ,n1381);
    nand g942(n2242 ,n2212 ,n2188);
    nand g943(n2578 ,n2690 ,n2546);
    nor g944(n1092 ,n960 ,n1077);
    dff g945(.RN(n1), .SN(1'b1), .CK(n0), .D(n419), .Q(n10[10]));
    nand g946(n337 ,n755 ,n141);
    nand g947(n248 ,n30[7] ,n140);
    nor g948(n55 ,n30[1] ,n30[0]);
    nand g949(n981 ,n816 ,n936);
    nand g950(n2267 ,n2246 ,n2234);
    nand g951(n381 ,n208 ,n284);
    buf g952(n13[28], n10[4]);
    nor g953(n2539 ,n2728 ,n32[5]);
    nor g954(n67 ,n25[1] ,n25[0]);
    nand g955(n2581 ,n32[7] ,n2561);
    or g956(n444 ,n155 ,n350);
    dff g957(.RN(n1), .SN(1'b1), .CK(n0), .D(n410), .Q(n25[3]));
    nor g958(n62 ,n30[5] ,n61);
    nand g959(n1893 ,n1724 ,n1789);
    nand g960(n432 ,n249 ,n311);
    nor g961(n111 ,n26[6] ,n26[7]);
    xnor g962(n2302 ,n2172 ,n2274);
    xor g963(n783 ,n21[0] ,n20[0]);
    nand g964(n1682 ,n20[0] ,n22[6]);
    xnor g965(n2711 ,n1206 ,n1262);
    nand g966(n896 ,n2715 ,n848);
    dff g967(.RN(n1), .SN(1'b1), .CK(n0), .D(n422), .Q(n10[8]));
    nor g968(n1217 ,n1203 ,n1191);
    nand g969(n2442 ,n22[3] ,n23[3]);
    nand g970(n2423 ,n2406 ,n2422);
    xnor g971(n2670 ,n2529 ,n2490);
    dff g972(.RN(n1), .SN(1'b1), .CK(n0), .D(n737), .Q(n9[1]));
    nand g973(n2659 ,n2590 ,n2640);
    nand g974(n796 ,n776 ,n779);
    nand g975(n1940 ,n1731 ,n1896);
    nand g976(n646 ,n540 ,n500);
    nand g977(n956 ,n873 ,n917);
    nand g978(n1781 ,n1670 ,n1674);
    buf g979(n9[11], 1'b0);
    not g980(n1948 ,n1947);
    xnor g981(n818 ,n801 ,n775);
    nand g982(n285 ,n29[4] ,n140);
    buf g983(n13[2], 1'b0);
    nand g984(n619 ,n24[2] ,n482);
    nand g985(n947 ,n869 ,n918);
    xnor g986(n1849 ,n1697 ,n1575);
    nand g987(n250 ,n29[15] ,n140);
    xnor g988(n2484 ,n2711 ,n2695);
    nand g989(n1653 ,n21[2] ,n23[0]);
    nand g990(n954 ,n867 ,n888);
    not g991(n345 ,n253);
    nand g992(n1691 ,n20[0] ,n22[2]);
    or g993(n1751 ,n1584 ,n1677);
    nor g994(n761 ,n20[7] ,n21[7]);
    buf g995(n9[8], 1'b0);
    not g996(n636 ,n610);
    nand g997(n348 ,n170 ,n169);
    nand g998(n2277 ,n2209 ,n2241);
    xnor g999(n2014 ,n1819 ,n1613);
    nand g1000(n540 ,n20[7] ,n465);
    or g1001(n2204 ,n2109 ,n2165);
    or g1002(n1464 ,n1431 ,n1449);
    or g1003(n2057 ,n1935 ,n1964);
    xnor g1004(n1069 ,n817 ,n995);
    nor g1005(n1375 ,n1289 ,n1335);
    buf g1006(n13[30], n10[6]);
    nand g1007(n769 ,n20[4] ,n20[3]);
    nor g1008(n1757 ,n1596 ,n1690);
    nand g1009(n2059 ,n1930 ,n1999);
    nor g1010(n1186 ,n1136 ,n1169);
    nor g1011(n108 ,n18[1] ,n18[2]);
    nand g1012(n226 ,n26[2] ,n87);
    nor g1013(n728 ,n638 ,n691);
    buf g1014(n9[22], 1'b0);
    nand g1015(n328 ,n10[1] ,n156);
    nand g1016(n197 ,n28[14] ,n140);
    nand g1017(n837 ,n2714 ,n821);
    nand g1018(n496 ,n6[5] ,n464);
    xnor g1019(n2324 ,n2284 ,n2272);
    nand g1020(n280 ,n28[12] ,n141);
    nand g1021(n1942 ,n1744 ,n1895);
    or g1022(n1739 ,n1605 ,n1671);
    nand g1023(n703 ,n572 ,n492);
    not g1024(n1116 ,n1115);
    nand g1025(n379 ,n207 ,n307);
    nand g1026(n2444 ,n22[5] ,n23[5]);
    xnor g1027(n2688 ,n2411 ,n2422);
    or g1028(n167 ,n87 ,n131);
    nand g1029(n643 ,n537 ,n499);
    nor g1030(n2512 ,n2502 ,n2511);
    nand g1031(n1085 ,n1020 ,n1047);
    xnor g1032(n1441 ,n1347 ,n1400);
    nand g1033(n663 ,n556 ,n488);
    nand g1034(n2232 ,n2123 ,n2179);
    nand g1035(n869 ,n2720 ,n819);
    nor g1036(n1082 ,n1000 ,n1061);
    or g1037(n1733 ,n1684 ,n1606);
    nand g1038(n275 ,n31[12] ,n141);
    nand g1039(n2238 ,n2167 ,n2205);
    nand g1040(n576 ,n22[4] ,n478);
    nand g1041(n597 ,n20[0] ,n468);
    xnor g1042(n2352 ,n2298 ,n2286);
    nor g1043(n2513 ,n2475 ,n2512);
    xnor g1044(n2378 ,n2304 ,n2350);
    nand g1045(n2629 ,n2578 ,n2609);
    nor g1046(n1761 ,n1725 ,n1649);
    or g1047(n1271 ,n2677 ,n23[5]);
    nor g1048(n1212 ,n1168 ,n1197);
    nand g1049(n2633 ,n2583 ,n2612);
    nand g1050(n563 ,n24[1] ,n461);
    xnor g1051(n1529 ,n1505 ,n1483);
    nor g1052(n1232 ,n1152 ,n1207);
    xnor g1053(n1842 ,n1574 ,n1683);
    xnor g1054(n822 ,n808 ,n761);
    xnor g1055(n2146 ,n2033 ,n1954);
    nand g1056(n593 ,n21[6] ,n467);
    nand g1057(n789 ,n2715 ,n783);
    nor g1058(n472 ,n252 ,n454);
    xnor g1059(n1183 ,n1148 ,n1115);
    xnor g1060(n1122 ,n1065 ,n757);
    xnor g1061(n2137 ,n2030 ,n1964);
    nand g1062(n701 ,n571 ,n491);
    xnor g1063(n2282 ,n2218 ,n2143);
    nand g1064(n671 ,n404 ,n596);
    buf g1065(n11[14], 1'b0);
    not g1066(n1452 ,n1451);
    nand g1067(n2162 ,n2041 ,n2118);
    nand g1068(n919 ,n844 ,n884);
    nand g1069(n702 ,n628 ,n627);
    nand g1070(n1769 ,n1597 ,n1669);
    xnor g1071(n1838 ,n1648 ,n1690);
    nor g1072(n1196 ,n1150 ,n1176);
    not g1073(n633 ,n591);
    xnor g1074(n1475 ,n1434 ,n1379);
    xnor g1075(n2502 ,n2701 ,n2685);
    xnor g1076(n1188 ,n1139 ,n1161);
    nand g1077(n249 ,n30[6] ,n140);
    nor g1078(n1292 ,n1268 ,n1283);
    nand g1079(n1785 ,n1696 ,n1664);
    xnor g1080(n2296 ,n2261 ,n2270);
    nand g1081(n416 ,n315 ,n230);
    not g1082(n1718 ,n1717);
    nor g1083(n2365 ,n2304 ,n2350);
    dff g1084(.RN(n1), .SN(1'b1), .CK(n0), .D(n355), .Q(n29[6]));
    nand g1085(n230 ,n31[13] ,n155);
    nand g1086(n2582 ,n2687 ,n2546);
    nand g1087(n1799 ,n1687 ,n1591);
    buf g1088(n13[23], 1'b0);
    nor g1089(n1043 ,n1016 ,n983);
    nand g1090(n227 ,n26[1] ,n87);
    nand g1091(n1673 ,n20[1] ,n22[3]);
    nand g1092(n384 ,n339 ,n255);
    nand g1093(n1580 ,n20[0] ,n22[5]);
    nand g1094(n2660 ,n2619 ,n2646);
    nand g1095(n271 ,n28[10] ,n141);
    buf g1096(n11[29], n10[13]);
    nand g1097(n601 ,n24[5] ,n482);
    nand g1098(n1513 ,n1483 ,n1495);
    nor g1099(n1376 ,n1320 ,n1340);
    nand g1100(n2600 ,n2665 ,n2561);
    or g1101(n1050 ,n994 ,n989);
    nand g1102(n2426 ,n2425 ,n2416);
    nand g1103(n431 ,n329 ,n247);
    nand g1104(n2291 ,n2270 ,n2261);
    nand g1105(n1230 ,n1212 ,n1188);
    dff g1106(.RN(n1), .SN(1'b1), .CK(n0), .D(n364), .Q(n28[9]));
    nand g1107(n2606 ,n2671 ,n2559);
    nand g1108(n1668 ,n21[4] ,n23[1]);
    buf g1109(n12[1], 1'b0);
    nand g1110(n2395 ,n2371 ,n2383);
    nor g1111(n1453 ,n1405 ,n1445);
    nor g1112(n103 ,n5[25] ,n5[24]);
    xnor g1113(n32[11] ,n1518 ,n1561);
    xnor g1114(n2704 ,n1222 ,n1246);
    nor g1115(n2535 ,n2725 ,n32[8]);
    xnor g1116(n1164 ,n1122 ,n1098);
    xor g1117(n820 ,n804 ,n810);
    nor g1118(n2566 ,n2560 ,n2540);
    nand g1119(n164 ,n107 ,n85);
    xnor g1120(n1825 ,n1692 ,n1587);
    nand g1121(n800 ,n768 ,n781);
    nand g1122(n2527 ,n2480 ,n2526);
    nand g1123(n414 ,n313 ,n233);
    xnor g1124(n771 ,n21[6] ,n21[5]);
    not g1125(n1586 ,n1585);
    or g1126(n1534 ,n1493 ,n1525);
    nand g1127(n705 ,n573 ,n524);
    xnor g1128(n1831 ,n1663 ,n1662);
    nor g1129(n1519 ,n1489 ,n1507);
    nand g1130(n32[12] ,n1511 ,n1562);
    nor g1131(n468 ,n252 ,n459);
    nand g1132(n375 ,n204 ,n332);
    nand g1133(n2243 ,n2162 ,n2182);
    not g1134(n1622 ,n1571);
    nor g1135(n1166 ,n1114 ,n1146);
    or g1136(n31[13] ,n2584 ,n2637);
    nand g1137(n383 ,n287 ,n338);
    xnor g1138(n2682 ,n2170 ,n2122);
    xnor g1139(n1860 ,n1710 ,n1698);
    xnor g1140(n1820 ,n1661 ,n1693);
    xnor g1141(n32[4] ,n1526 ,n1524);
    not g1142(n1432 ,n1424);
    dff g1143(.RN(n1), .SN(1'b1), .CK(n0), .D(n377), .Q(n28[4]));
    nand g1144(n2651 ,n2558 ,n2571);
    not g1145(n2347 ,n2346);
    nand g1146(n36 ,n34 ,n33);
    nand g1147(n791 ,n2714 ,n783);
    not g1148(n1009 ,n1008);
    xnor g1149(n1193 ,n1142 ,n1117);
    nand g1150(n652 ,n545 ,n505);
    xnor g1151(n824 ,n803 ,n795);
    nand g1152(n244 ,n28[13] ,n140);
    nor g1153(n1765 ,n1643 ,n1636);
    nand g1154(n287 ,n740 ,n141);
    nand g1155(n2384 ,n2322 ,n2359);
    nand g1156(n430 ,n328 ,n187);
    nand g1157(n309 ,n746 ,n143);
    or g1158(n1931 ,n1873 ,n1863);
    nand g1159(n259 ,n27[1] ,n155);
    nor g1160(n1020 ,n967 ,n979);
    xnor g1161(n1970 ,n1829 ,n1632);
    xnor g1162(n1539 ,n1517 ,n1515);
    nand g1163(n1246 ,n1209 ,n1245);
    nor g1164(n721 ,n706 ,n702);
    dff g1165(.RN(n1), .SN(1'b1), .CK(n0), .D(n353), .Q(n29[3]));
    xnor g1166(n2093 ,n1985 ,n1936);
    nand g1167(n2645 ,n2553 ,n2568);
    nand g1168(n150 ,n118 ,n111);
    nor g1169(n1446 ,n1381 ,n1430);
    nor g1170(n1081 ,n996 ,n1060);
    nand g1171(n353 ,n301 ,n168);
    nand g1172(n1782 ,n1596 ,n1690);
    xnor g1173(n2220 ,n2129 ,n2141);
    xnor g1174(n1437 ,n1388 ,n1370);
    nand g1175(n1615 ,n20[6] ,n22[0]);
    not g1176(n1106 ,n1105);
    nand g1177(n247 ,n31[0] ,n155);
    nor g1178(n171 ,n151 ,n153);
    nand g1179(n810 ,n784 ,n802);
    nand g1180(n793 ,n2717 ,n783);
    xnor g1181(n2494 ,n2707 ,n2691);
    nand g1182(n1795 ,n1605 ,n1671);
    buf g1183(n12[27], 1'b0);
    nand g1184(n258 ,n30[1] ,n87);
    nand g1185(n1591 ,n21[4] ,n23[3]);
    nand g1186(n1929 ,n1768 ,n1904);
    nand g1187(n854 ,n2719 ,n821);
    nand g1188(n2412 ,n2393 ,n2404);
    nand g1189(n1514 ,n1444 ,n1497);
    nor g1190(n1180 ,n1040 ,n1156);
    xnor g1191(n2215 ,n2146 ,n1962);
    nand g1192(n1521 ,n1481 ,n1508);
    xnor g1193(n2694 ,n2376 ,n2434);
    nand g1194(n395 ,n266 ,n342);
    nand g1195(n682 ,n558 ,n512);
    nor g1196(n1449 ,n1387 ,n1416);
    nor g1197(n1407 ,n1371 ,n1376);
    nand g1198(n920 ,n854 ,n914);
    nor g1199(n1254 ,n1253 ,n1239);
    nand g1200(n68 ,n25[1] ,n25[0]);
    nand g1201(n1688 ,n21[1] ,n23[0]);
    or g1202(n1497 ,n1442 ,n1475);
    nand g1203(n1628 ,n20[6] ,n22[1]);
    nor g1204(n1293 ,n1268 ,n1282);
    nand g1205(n293 ,n29[10] ,n141);
    nor g1206(n119 ,n93 ,n18[1]);
    nand g1207(n2577 ,n2686 ,n2546);
    nand g1208(n447 ,n156 ,n359);
    nand g1209(n491 ,n6[1] ,n475);
    dff g1210(.RN(n1), .SN(1'b1), .CK(n0), .D(n428), .Q(n10[2]));
    nand g1211(n246 ,n31[2] ,n155);
    not g1212(n1723 ,n1722);
    not g1213(n2375 ,n2366);
    nand g1214(n901 ,n790 ,n856);
    xnor g1215(n2410 ,n2388 ,n2395);
    nor g1216(n1250 ,n1213 ,n1249);
    xnor g1217(n2307 ,n2253 ,n2162);
    not g1218(n929 ,n930);
    nand g1219(n534 ,n21[5] ,n463);
    nand g1220(n2604 ,n32[12] ,n2561);
    not g1221(n140 ,n141);
    nand g1222(n202 ,n28[8] ,n87);
    dff g1223(.RN(n1), .SN(1'b1), .CK(n0), .D(n370), .Q(n29[8]));
    or g1224(n2437 ,n22[1] ,n23[1]);
    nor g1225(n1098 ,n1030 ,n1078);
    not g1226(n1203 ,n1202);
    xor g1227(n1843 ,n1724 ,n1678);
    nand g1228(n2422 ,n2392 ,n2418);
    nor g1229(n96 ,n5[5] ,n5[4]);
    xnor g1230(n2342 ,n2268 ,n2301);
    xnor g1231(n2261 ,n2173 ,n2133);
    not g1232(n1667 ,n1666);
    nand g1233(n1678 ,n20[5] ,n22[5]);
    xor g1234(n2675 ,n20[3] ,n21[3]);
    xnor g1235(n1961 ,n1828 ,n1634);
    nor g1236(n39 ,n30[7] ,n38);
    nor g1237(n170 ,n26[0] ,n154);
    not g1238(n1266 ,n24[2]);
    nor g1239(n1174 ,n1157 ,n1160);
    nand g1240(n2430 ,n2429 ,n2417);
    nand g1241(n2579 ,n2693 ,n2546);
    xnor g1242(n969 ,n807 ,n907);
    buf g1243(n10[16], 1'b0);
    xnor g1244(n1850 ,n1582 ,n1651);
    nand g1245(n198 ,n25[5] ,n142);
    nand g1246(n2463 ,n2441 ,n2462);
    nand g1247(n272 ,n31[8] ,n141);
    or g1248(n2330 ,n2271 ,n2306);
    xor g1249(n2676 ,n20[4] ,n21[4]);
    xnor g1250(n1455 ,n1402 ,n1380);
    nor g1251(n1324 ,n1268 ,n1284);
    or g1252(n1527 ,n1514 ,n1516);
    nand g1253(n2590 ,n2682 ,n2546);
    xor g1254(n2022 ,n1851 ,n1705);
    nand g1255(n267 ,n28[13] ,n141);
    nand g1256(n512 ,n6[7] ,n462);
    xnor g1257(n2032 ,n1852 ,n1947);
    xnor g1258(n1457 ,n1403 ,n1378);
    or g1259(n1996 ,n1955 ,n1914);
    or g1260(n2245 ,n2196 ,n2193);
    xnor g1261(n1985 ,n1826 ,n1608);
    xnor g1262(n988 ,n921 ,n816);
    nand g1263(n2241 ,n2021 ,n2198);
    nand g1264(n507 ,n6[6] ,n477);
    dff g1265(.RN(n1), .SN(1'b1), .CK(n0), .D(n443), .Q(n18[1]));
    xnor g1266(n1187 ,n1141 ,n1125);
    nor g1267(n106 ,n5[29] ,n5[28]);
    nor g1268(n1724 ,n1567 ,n1568);
    buf g1269(n10[20], 1'b0);
    nor g1270(n1157 ,n1058 ,n1118);
    nand g1271(n2049 ,n1913 ,n2007);
    nand g1272(n504 ,n6[3] ,n466);
    nand g1273(n2157 ,n2054 ,n2105);
    buf g1274(n12[5], 1'b0);
    nand g1275(n187 ,n31[1] ,n155);
    nor g1276(n1045 ,n1007 ,n993);
    nand g1277(n1546 ,n1521 ,n1535);
    xnor g1278(n32[3] ,n1504 ,n1501);
    nand g1279(n2465 ,n2444 ,n2464);
    dff g1280(.RN(n1), .SN(1'b1), .CK(n0), .D(n649), .Q(n20[4]));
    not g1281(n1038 ,n756);
    nand g1282(n1933 ,n1691 ,n1860);
    nand g1283(n200 ,n28[11] ,n87);
    nand g1284(n2530 ,n2491 ,n2529);
    nand g1285(n602 ,n23[5] ,n480);
    dff g1286(.RN(n1), .SN(1'b1), .CK(n0), .D(n693), .Q(n23[7]));
    buf g1287(n10[23], 1'b0);
    nand g1288(n149 ,n109 ,n110);
    buf g1289(n12[19], n10[11]);
    nand g1290(n1777 ,n1582 ,n1651);
    nor g1291(n2514 ,n2503 ,n2513);
    nand g1292(n2351 ,n2316 ,n2337);
    or g1293(n1759 ,n1588 ,n1601);
    xnor g1294(n2248 ,n2157 ,n2213);
    dff g1295(.RN(n1), .SN(1'b1), .CK(n0), .D(n354), .Q(n29[1]));
    or g1296(n31[8] ,n2643 ,n2664);
    nand g1297(n2034 ,n1921 ,n1987);
    nand g1298(n607 ,n24[4] ,n482);
    nand g1299(n1562 ,n1510 ,n1561);
    not g1300(n759 ,n2716);
    nand g1301(n628 ,n21[1] ,n467);
    not g1302(n2534 ,n2669);
    nand g1303(n1679 ,n20[1] ,n22[0]);
    not g1304(n774 ,n773);
    or g1305(n2045 ,n1944 ,n1963);
    nor g1306(n1208 ,n1181 ,n1187);
    xnor g1307(n2102 ,n1958 ,n1766);
    xnor g1308(n2132 ,n2023 ,n1982);
    xnor g1309(n807 ,n773 ,n770);
    nand g1310(n148 ,n125 ,n104);
    xnor g1311(n816 ,n802 ,n784);
    xnor g1312(n2170 ,n1565 ,n1979);
    nand g1313(n548 ,n19[7] ,n476);
    buf g1314(n13[15], 1'b0);
    nor g1315(n1809 ,n1647 ,n1715);
    nor g1316(n122 ,n91 ,n5[5]);
    nor g1317(n143 ,n18[1] ,n128);
    nand g1318(n915 ,n2712 ,n876);
    xnor g1319(n2103 ,n1994 ,n1955);
    nand g1320(n2331 ,n2247 ,n2313);
    buf g1321(n10[30], 1'b0);
    nand g1322(n1409 ,n1326 ,n1397);
    nand g1323(n153 ,n115 ,n103);
    xnor g1324(n990 ,n946 ,n818);
    buf g1325(n12[30], 1'b0);
    xnor g1326(n2260 ,n2174 ,n2161);
    xnor g1327(n997 ,n818 ,n948);
    or g1328(n1052 ,n1015 ,n984);
    xnor g1329(n2189 ,n2085 ,n2018);
    or g1330(n2332 ,n2278 ,n2307);
    nand g1331(n951 ,n868 ,n892);
    dff g1332(.RN(n1), .SN(1'b1), .CK(n0), .D(n714), .Q(n22[0]));
    nor g1333(n2511 ,n2473 ,n2510);
    xnor g1334(n1226 ,n1185 ,n1145);
    nor g1335(n2106 ,n1991 ,n2077);
    nand g1336(n237 ,n31[11] ,n155);
    buf g1337(n9[28], 1'b0);
    nand g1338(n413 ,n9[5] ,n252);
    nand g1339(n2429 ,n2428 ,n2415);
    nand g1340(n570 ,n23[2] ,n474);
    nor g1341(n727 ,n637 ,n681);
    xnor g1342(n995 ,n941 ,n818);
    nor g1343(n113 ,n5[31] ,n5[30]);
    nand g1344(n710 ,n577 ,n528);
    xnor g1345(n2725 ,n2503 ,n2513);
    xnor g1346(n2719 ,n2448 ,n2467);
    nand g1347(n2006 ,n1928 ,n1911);
    xnor g1348(n2703 ,n1228 ,n1244);
    nand g1349(n1424 ,n1395 ,n1372);
    xnor g1350(n2503 ,n2702 ,n2686);
    nand g1351(n572 ,n23[0] ,n474);
    nand g1352(n269 ,n28[9] ,n141);
    dff g1353(.RN(n1), .SN(1'b1), .CK(n0), .D(n398), .Q(n26[5]));
    nand g1354(n152 ,n100 ,n101);
    buf g1355(n13[7], 1'b0);
    nand g1356(n845 ,n2715 ,n821);
    dff g1357(.RN(n1), .SN(1'b1), .CK(n0), .D(n644), .Q(n21[1]));
    nand g1358(n1035 ,n1006 ,n988);
    nand g1359(n1866 ,n1595 ,n1761);
    nand g1360(n714 ,n580 ,n494);
    not g1361(n2455 ,n2454);
    or g1362(n31[2] ,n2642 ,n2659);
    nand g1363(n307 ,n31[2] ,n141);
    nor g1364(n1135 ,n756 ,n1106);
    nor g1365(n1477 ,n1454 ,n1455);
    nand g1366(n1683 ,n20[7] ,n22[5]);
    nand g1367(n879 ,n2717 ,n848);
    nand g1368(n242 ,n28[5] ,n87);
    nand g1369(n797 ,n778 ,n771);
    nor g1370(n1388 ,n1318 ,n1344);
    dff g1371(.RN(n1), .SN(1'b1), .CK(n0), .D(n351), .Q(n29[7]));
    nand g1372(n1930 ,n1739 ,n1901);
    nor g1373(n2720 ,n2438 ,n2468);
    nand g1374(n552 ,n19[3] ,n476);
    nand g1375(n675 ,n606 ,n605);
    nand g1376(n698 ,n569 ,n522);
    nand g1377(n2396 ,n2360 ,n2384);
    not g1378(n1859 ,n1858);
    nand g1379(n2266 ,n2214 ,n2223);
    buf g1380(n11[3], 1'b0);
    nand g1381(n2441 ,n22[4] ,n23[4]);
    xnor g1382(n2402 ,n2349 ,n2382);
    dff g1383(.RN(n1), .SN(1'b1), .CK(n0), .D(n713), .Q(n22[1]));
    nand g1384(n310 ,n747 ,n143);
    xnor g1385(n1832 ,n1605 ,n1671);
    nand g1386(n672 ,n600 ,n599);
    nand g1387(n1693 ,n21[2] ,n23[3]);
    dff g1388(.RN(n1), .SN(1'b1), .CK(n0), .D(n442), .Q(n26[7]));
    buf g1389(n12[22], n10[14]);
    buf g1390(n13[16], 1'b0);
    nand g1391(n1919 ,n1742 ,n1891);
    nand g1392(n1788 ,n1672 ,n1577);
    dff g1393(.RN(n1), .SN(1'b1), .CK(n0), .D(n438), .Q(n28[14]));
    nand g1394(n391 ,n248 ,n341);
    nand g1395(n376 ,n242 ,n281);
    buf g1396(n12[14], n10[6]);
    nor g1397(n61 ,n54 ,n60);
    xnor g1398(n970 ,n902 ,n816);
    nand g1399(n1789 ,n1678 ,n1694);
    nand g1400(n924 ,n835 ,n882);
    xnor g1401(n1962 ,n1850 ,n1717);
    xnor g1402(n2219 ,n2166 ,n2140);
    nand g1403(n500 ,n6[7] ,n466);
    nor g1404(n1372 ,n1314 ,n1342);
    buf g1405(n11[4], 1'b0);
    nor g1406(n347 ,n180 ,n184);
    nand g1407(n917 ,n2719 ,n846);
    nor g1408(n1370 ,n1321 ,n1350);
    not g1409(n637 ,n616);
    nand g1410(n1897 ,n1718 ,n1777);
    xnor g1411(n32[7] ,n1547 ,n1553);
    not g1412(n1938 ,n1937);
    not g1413(n1946 ,n1945);
    nand g1414(n1612 ,n21[3] ,n23[3]);
    nor g1415(n102 ,n5[11] ,n5[10]);
    nand g1416(n273 ,n31[11] ,n141);
    nor g1417(n127 ,n92 ,n18[0]);
    nand g1418(n583 ,n19[0] ,n481);
    buf g1419(n13[24], n10[0]);
    not g1420(n1813 ,n1791);
    dff g1421(.RN(n1), .SN(1'b1), .CK(n0), .D(n372), .Q(n29[13]));
    nand g1422(n670 ,n632 ,n594);
    xnor g1423(n2339 ,n2053 ,n2308);
    not g1424(n1646 ,n1572);
    xnor g1425(n2046 ,n1822 ,n1957);
    xnor g1426(n2192 ,n2093 ,n2104);
    nand g1427(n394 ,n171 ,n177);
    dff g1428(.RN(n1), .SN(1'b1), .CK(n0), .D(n664), .Q(n27[0]));
    xnor g1429(n1148 ,n1003 ,n1108);
    nand g1430(n270 ,n28[8] ,n141);
    nand g1431(n910 ,n2713 ,n876);
    nand g1432(n1167 ,n1109 ,n1144);
    xnor g1433(n1433 ,n1375 ,n1373);
    nand g1434(n1722 ,n21[6] ,n23[2]);
    nand g1435(n1665 ,n20[4] ,n22[3]);
    nand g1436(n382 ,n286 ,n259);
    nor g1437(n2518 ,n2485 ,n2517);
    xnor g1438(n1840 ,n1642 ,n1653);
    or g1439(n2224 ,n2212 ,n2188);
    nor g1440(n1312 ,n1269 ,n1285);
    not g1441(n66 ,n25[4]);
    nand g1442(n2078 ,n1909 ,n2011);
    nand g1443(n291 ,n29[12] ,n141);
    or g1444(n1348 ,n1268 ,n1305);
    nand g1445(n2624 ,n2556 ,n2572);
    nand g1446(n1587 ,n21[6] ,n23[0]);
    xnor g1447(n752 ,n30[4] ,n60);
    nand g1448(n547 ,n20[0] ,n465);
    nor g1449(n2666 ,n1426 ,n1414);
    xnor g1450(n1851 ,n1696 ,n1664);
    dff g1451(.RN(n1), .SN(1'b1), .CK(n0), .D(n363), .Q(n29[10]));
    nand g1452(n906 ,n793 ,n861);
    nor g1453(n1443 ,n1399 ,n1418);
    xnor g1454(n1006 ,n949 ,n817);
    xnor g1455(n2253 ,n2181 ,n2149);
    not g1456(n1060 ,n1042);
    nand g1457(n567 ,n23[5] ,n474);
    nor g1458(n1339 ,n1267 ,n1307);
    xnor g1459(n2024 ,n1919 ,n1939);
    nand g1460(n736 ,n722 ,n715);
    not g1461(n1853 ,n1852);
    dff g1462(.RN(n1), .SN(1'b1), .CK(n0), .D(n391), .Q(n30[7]));
    dff g1463(.RN(n1), .SN(1'b1), .CK(n0), .D(n690), .Q(n24[1]));
    nand g1464(n1422 ,n1371 ,n1376);
    nand g1465(n339 ,n17[3] ,n156);
    nand g1466(n1647 ,n20[6] ,n22[3]);
    nand g1467(n2555 ,n2727 ,n32[6]);
    nand g1468(n513 ,n6[6] ,n462);
    or g1469(n2151 ,n2066 ,n2104);
    xnor g1470(n2448 ,n23[7] ,n22[7]);
    nand g1471(n2122 ,n1866 ,n2071);
    nor g1472(n1351 ,n1266 ,n1298);
    nand g1473(n1421 ,n1373 ,n1375);
    not g1474(n1721 ,n1720);
    nand g1475(n2556 ,n2721 ,n32[12]);
    dff g1476(.RN(n1), .SN(1'b1), .CK(n0), .D(n448), .Q(n15));
    xnor g1477(n2251 ,n2160 ,n2189);
    nand g1478(n627 ,n22[1] ,n469);
    nand g1479(n2167 ,n2044 ,n2115);
    nand g1480(n458 ,n83 ,n80);
    xnor g1481(n998 ,n816 ,n936);
    nand g1482(n1585 ,n21[5] ,n23[0]);
    nor g1483(n2165 ,n2035 ,n2112);
    nand g1484(n412 ,n262 ,n312);
    nor g1485(n180 ,n740 ,n140);
    or g1486(n1744 ,n1697 ,n1575);
    nor g1487(n719 ,n688 ,n685);
    nand g1488(n422 ,n320 ,n239);
    or g1489(n82 ,n157 ,n394);
    nand g1490(n2208 ,n2122 ,n2152);
    xnor g1491(n1821 ,n1672 ,n1577);
    buf g1492(n10[17], 1'b0);
    or g1493(n1520 ,n1481 ,n1508);
    nand g1494(n1042 ,n1016 ,n983);
    nor g1495(n1448 ,n1368 ,n1412);
    nor g1496(n1318 ,n1269 ,n1280);
    nand g1497(n1054 ,n931 ,n990);
    nand g1498(n316 ,n10[12] ,n156);
    nor g1499(n2111 ,n1992 ,n2082);
    nand g1500(n575 ,n22[5] ,n478);
    nand g1501(n1579 ,n21[1] ,n23[5]);
    nand g1502(n900 ,n791 ,n857);
    nand g1503(n302 ,n29[1] ,n141);
    xnor g1504(n2487 ,n2705 ,n2689);
    xnor g1505(n1976 ,n1827 ,n1722);
    nand g1506(n2335 ,n2276 ,n2312);
    nand g1507(n222 ,n29[13] ,n140);
    dff g1508(.RN(n1), .SN(1'b1), .CK(n0), .D(n689), .Q(n24[2]));
    nand g1509(n1710 ,n20[1] ,n22[1]);
    nand g1510(n434 ,n9[2] ,n252);
    nand g1511(n2348 ,n2275 ,n2327);
    xnor g1512(n1528 ,n1502 ,n1482);
    nor g1513(n1953 ,n1740 ,n1894);
    dff g1514(.RN(n1), .SN(1'b1), .CK(n0), .D(n657), .Q(n19[6]));
    xor g1515(n2729 ,n2496 ,n2505);
    nor g1516(n717 ,n676 ,n675);
    nand g1517(n1662 ,n21[4] ,n23[2]);
    nand g1518(n126 ,n18[1] ,n18[2]);
    nand g1519(n1896 ,n1703 ,n1783);
    nor g1520(n80 ,n164 ,n82);
    nor g1521(n762 ,n20[1] ,n21[1]);
    nand g1522(n2634 ,n2600 ,n2613);
    nand g1523(n886 ,n2713 ,n847);
    nor g1524(n2546 ,n2533 ,n27[1]);
    nand g1525(n2409 ,n2356 ,n2400);
    nand g1526(n255 ,n27[0] ,n155);
    nand g1527(n1717 ,n21[6] ,n23[7]);
    nand g1528(n1957 ,n1749 ,n1886);
    or g1529(n1768 ,n1603 ,n1665);
    nand g1530(n858 ,n2715 ,n825);
    nand g1531(n1573 ,n21[7] ,n23[0]);
    nor g1532(n2472 ,n2702 ,n2686);
    or g1533(n2054 ,n1921 ,n1987);
    or g1534(n1425 ,n1394 ,n1391);
    nor g1535(n912 ,n759 ,n875);
    xnor g1536(n1120 ,n1064 ,n1090);
    buf g1537(n11[7], 1'b0);
    or g1538(n2128 ,n2119 ,n2052);
    not g1539(n471 ,n470);
    nand g1540(n2117 ,n1975 ,n2046);
    not g1541(n2187 ,n2186);
    nor g1542(n479 ,n344 ,n455);
    nand g1543(n802 ,n769 ,n782);
    or g1544(n1545 ,n1519 ,n1528);
    nand g1545(n2079 ,n1867 ,n2008);
    nand g1546(n893 ,n2712 ,n847);
    nor g1547(n1057 ,n1004 ,n1018);
    nand g1548(n890 ,n2716 ,n846);
    nor g1549(n1004 ,n850 ,n964);
    dff g1550(.RN(n1), .SN(1'b1), .CK(n0), .D(n697), .Q(n23[4]));
    or g1551(n183 ,n3 ,n138);
    nand g1552(n1558 ,n1543 ,n1557);
    nor g1553(n34 ,n30[3] ,n30[2]);
    nand g1554(n305 ,n743 ,n143);
    xnor g1555(n1982 ,n1834 ,n1699);
    dff g1556(.RN(n1), .SN(1'b1), .CK(n0), .D(n710), .Q(n22[3]));
    nand g1557(n355 ,n191 ,n173);
    dff g1558(.RN(n1), .SN(1'b1), .CK(n0), .D(n733), .Q(n9[5]));
    nor g1559(n2568 ,n2560 ,n2539);
    nor g1560(n2109 ,n2015 ,n2047);
    nand g1561(n439 ,n264 ,n330);
    or g1562(n31[4] ,n2649 ,n2662);
    xnor g1563(n1112 ,n1076 ,n960);
    xnor g1564(n2707 ,n1241 ,n1253);
    xnor g1565(n1505 ,n1447 ,n1471);
    nand g1566(n2213 ,n2117 ,n2150);
    not g1567(n1763 ,n1762);
    nand g1568(n1623 ,n21[0] ,n23[4]);
    nor g1569(n1107 ,n1037 ,n1088);
    buf g1570(n11[0], 1'b0);
    or g1571(n31[3] ,n2647 ,n2661);
    nand g1572(n397 ,n9[7] ,n252);
    xnor g1573(n784 ,n20[5] ,n21[5]);
    not g1574(n69 ,n68);
    dff g1575(.RN(n1), .SN(1'b1), .CK(n0), .D(n374), .Q(n28[7]));
    nand g1576(n403 ,n227 ,n302);
    not g1577(n1943 ,n1942);
    buf g1578(n11[28], n10[12]);
    nand g1579(n2158 ,n2057 ,n2095);
    not g1580(n1569 ,n21[4]);
    nand g1581(n2200 ,n2120 ,n2158);
    nand g1582(n1630 ,n21[4] ,n23[4]);
    xnor g1583(n1024 ,n849 ,n964);
    nor g1584(n2035 ,n1978 ,n1977);
    nand g1585(n1363 ,n24[0] ,n1297);
    nand g1586(n2596 ,n2683 ,n2546);
    nor g1587(n748 ,n69 ,n67);
    nand g1588(n327 ,n10[2] ,n156);
    nor g1589(n1625 ,n1567 ,n1570);
    xnor g1590(n1436 ,n1376 ,n1371);
    dff g1591(.RN(n1), .SN(1'b1), .CK(n0), .D(n654), .Q(n20[0]));
    xnor g1592(n1140 ,n1089 ,n1110);
    not g1593(n1268 ,n24[0]);
    nand g1594(n1648 ,n21[4] ,n23[6]);
    nand g1595(n1626 ,n20[3] ,n22[0]);
    not g1596(n38 ,n37);
    nand g1597(n1783 ,n1661 ,n1693);
    nor g1598(n2570 ,n2560 ,n2542);
    nand g1599(n1551 ,n1531 ,n1550);
    buf g1600(n12[15], n10[7]);
    nand g1601(n693 ,n565 ,n518);
    nand g1602(n1564 ,n21[0] ,n23[1]);
    nand g1603(n1707 ,n20[6] ,n22[2]);
    nand g1604(n923 ,n829 ,n881);
    nand g1605(n529 ,n6[2] ,n479);
    xnor g1606(n2447 ,n23[6] ,n22[6]);
    xnor g1607(n987 ,n919 ,n818);
    nor g1608(n2567 ,n2560 ,n2541);
    nand g1609(n147 ,n123 ,n85);
    nand g1610(n239 ,n31[8] ,n155);
    nand g1611(n2003 ,n1919 ,n1939);
    nand g1612(n950 ,n863 ,n887);
    nor g1613(n2076 ,n1940 ,n1984);
    xnor g1614(n1530 ,n1503 ,n1484);
    dff g1615(.RN(n1), .SN(1'b1), .CK(n0), .D(n373), .Q(n28[8]));
    nand g1616(n2456 ,n2440 ,n2450);
    xnor g1617(n2445 ,n23[4] ,n22[4]);
    not g1618(n1181 ,n1180);
    nor g1619(n2072 ,n1943 ,n1980);
    nand g1620(n613 ,n24[3] ,n482);
    nand g1621(n511 ,n6[2] ,n477);
    buf g1622(n12[18], n10[10]);
    not g1623(n1366 ,n1365);
    xnor g1624(n1117 ,n1070 ,n1020);
    nand g1625(n303 ,n29[0] ,n141);
    nor g1626(n931 ,n834 ,n912);
    nand g1627(n1506 ,n1482 ,n1490);
    nor g1628(n1413 ,n1332 ,n1398);
    xnor g1629(n1833 ,n1673 ,n1600);
    xnor g1630(n1171 ,n1068 ,n1124);
    nand g1631(n684 ,n559 ,n514);
    or g1632(n173 ,n87 ,n139);
    nand g1633(n2271 ,n2201 ,n2245);
    nand g1634(n282 ,n31[3] ,n141);
    xnor g1635(n2135 ,n2027 ,n1963);
    not g1636(n1075 ,n1074);
    not g1637(n1302 ,n1303);
    xnor g1638(n2126 ,n2080 ,n1966);
    not g1639(n876 ,n875);
    xnor g1640(n1989 ,n1848 ,n1688);
    xnor g1641(n785 ,n20[3] ,n21[3]);
    nand g1642(n1103 ,n1052 ,n1086);
    nand g1643(n877 ,n2712 ,n848);
    nand g1644(n1774 ,n1607 ,n1578);
    nand g1645(n688 ,n621 ,n619);
    nand g1646(n2021 ,n1868 ,n1932);
    or g1647(n2194 ,n2051 ,n2161);
    nand g1648(n443 ,n165 ,n347);
    or g1649(n1540 ,n1522 ,n1529);
    nand g1650(n304 ,n742 ,n143);
    nand g1651(n2205 ,n1962 ,n2146);
    or g1652(n2470 ,n2697 ,n2681);
    or g1653(n181 ,n739 ,n142);
    not g1654(n2320 ,n2319);
    not g1655(n1808 ,n1807);
    xnor g1656(n2303 ,n2254 ,n2214);
    not g1657(n927 ,n928);
    nand g1658(n1905 ,n1633 ,n1805);
    nand g1659(n1525 ,n1492 ,n1512);
    dff g1660(.RN(n1), .SN(1'b1), .CK(n0), .D(n346), .Q(n30[0]));
    xnor g1661(n772 ,n21[4] ,n21[3]);
    xnor g1662(n2133 ,n2026 ,n1983);
    nor g1663(n1028 ,n962 ,n1011);
    not g1664(n1211 ,n1210);
    xnor g1665(n1063 ,n996 ,n1016);
    nand g1666(n417 ,n316 ,n236);
    nand g1667(n862 ,n2719 ,n820);
    nand g1668(n517 ,n6[2] ,n462);
    or g1669(n1741 ,n1599 ,n1590);
    or g1670(n460 ,n179 ,n78);
    xnor g1671(n2700 ,n1165 ,n1160);
    or g1672(n1750 ,n1673 ,n1600);
    nand g1673(n1790 ,n1675 ,n1668);
    nor g1674(n1095 ,n1031 ,n1079);
    xnor g1675(n2323 ,n2292 ,n2285);
    nand g1676(n1890 ,n1700 ,n1792);
    xnor g1677(n938 ,n817 ,n853);
    or g1678(n1411 ,n1390 ,n1374);
    xnor g1679(n2346 ,n2297 ,n2303);
    or g1680(n178 ,n87 ,n130);
    nand g1681(n1698 ,n20[2] ,n22[0]);
    or g1682(n1273 ,n2672 ,n23[0]);
    not g1683(n1041 ,n1035);
    not g1684(n964 ,n963);
    nor g1685(n1286 ,n1266 ,n1282);
    not g1686(n1611 ,n1610);
    not g1687(n966 ,n965);
    xnor g1688(n994 ,n924 ,n818);
    nand g1689(n216 ,n26[13] ,n87);
    nand g1690(n2038 ,n1918 ,n1965);
    nand g1691(n1775 ,n1603 ,n1665);
    nand g1692(n861 ,n2716 ,n825);
    xnor g1693(n2127 ,n2046 ,n1974);
    nand g1694(n1034 ,n958 ,n1012);
    nand g1695(n2531 ,n2479 ,n2530);
    nand g1696(n2528 ,n2498 ,n2527);
    nand g1697(n367 ,n199 ,n275);
    nor g1698(n1489 ,n1458 ,n1472);
    nand g1699(n300 ,n29[2] ,n141);
    nor g1700(n79 ,n147 ,n82);
    not g1701(n1014 ,n1013);
    nor g1702(n1210 ,n1170 ,n1186);
    nor g1703(n722 ,n678 ,n651);
    xnor g1704(n2403 ,n2377 ,n2363);
    buf g1705(n9[20], 1'b0);
    xnor g1706(n2686 ,n2380 ,n2390);
    not g1707(n1633 ,n1632);
    xnor g1708(n1018 ,n817 ,n950);
    nand g1709(n622 ,n19[2] ,n481);
    buf g1710(n13[11], 1'b0);
    buf g1711(n11[18], n10[2]);
    nand g1712(n620 ,n20[2] ,n468);
    xnor g1713(n2388 ,n2342 ,n2354);
    not g1714(n1362 ,n1361);
    nand g1715(n2206 ,n2051 ,n2161);
    not g1716(n1621 ,n1620);
    nand g1717(n219 ,n26[10] ,n87);
    xor g1718(n1848 ,n1563 ,n1679);
    nand g1719(n312 ,n748 ,n143);
    nand g1720(n1696 ,n20[2] ,n22[6]);
    xnor g1721(n1823 ,n1689 ,n1654);
    nand g1722(n402 ,n9[0] ,n252);
    nand g1723(n494 ,n6[0] ,n479);
    nand g1724(n695 ,n567 ,n520);
    dff g1725(.RN(n1), .SN(1'b1), .CK(n0), .D(n396), .Q(n26[6]));
    xnor g1726(n2217 ,n2120 ,n2158);
    buf g1727(n13[10], 1'b0);
    nor g1728(n1745 ,n1589 ,n1652);
    nor g1729(n1252 ,n1251 ,n1238);
    nor g1730(n49 ,n25[6] ,n25[5]);
    nor g1731(n1108 ,n1055 ,n1083);
    not g1732(n1811 ,n1778);
    xnor g1733(n32[10] ,n1537 ,n1559);
    xnor g1734(n1822 ,n1684 ,n1606);
    xnor g1735(n346 ,n140 ,n30[0]);
    nand g1736(n588 ,n24[7] ,n482);
    nor g1737(n976 ,n807 ,n927);
    nand g1738(n1787 ,n1695 ,n1686);
    xnor g1739(n750 ,n30[6] ,n63);
    xnor g1740(n1861 ,n1643 ,n1636);
    xnor g1741(n2306 ,n2251 ,n2262);
    nand g1742(n1282 ,n2672 ,n23[0]);
    nand g1743(n782 ,n21[4] ,n764);
    xor g1744(n1818 ,n1646 ,n1598);
    xnor g1745(n1988 ,n1849 ,n1630);
    nand g1746(n1307 ,n1283 ,n1270);
    or g1747(n176 ,n87 ,n135);
    dff g1748(.RN(n1), .SN(1'b1), .CK(n0), .D(n358), .Q(n29[4]));
    xnor g1749(n1016 ,n956 ,n817);
    nand g1750(n578 ,n22[2] ,n478);
    or g1751(n2113 ,n2020 ,n2083);
    not g1752(n1941 ,n1940);
    nand g1753(n1032 ,n817 ,n992);
    not g1754(n2160 ,n2159);
    or g1755(n2368 ,n2280 ,n2352);
    nor g1756(n2473 ,n2700 ,n2684);
    nand g1757(n386 ,n214 ,n289);
    nand g1758(n488 ,n6[0] ,n477);
    nand g1759(n406 ,n212 ,n304);
    not g1760(n1595 ,n1594);
    dff g1761(.RN(n1), .SN(1'b1), .CK(n0), .D(n703), .Q(n23[0]));
    nor g1762(n1358 ,n1269 ,n1303);
    xnor g1763(n2727 ,n2500 ,n2509);
    nand g1764(n1772 ,n1673 ,n1600);
    dff g1765(.RN(n1), .SN(1'b1), .CK(n0), .D(n684), .Q(n24[5]));
    xnor g1766(n1978 ,n1832 ,n1644);
    not g1767(n64 ,n63);
    nand g1768(n686 ,n560 ,n515);
    xnor g1769(n749 ,n65 ,n30[7]);
    not g1770(n89 ,n5[2]);
    nor g1771(n1315 ,n1269 ,n1279);
    nand g1772(n2526 ,n2489 ,n2525);
    nor g1773(n1168 ,n1113 ,n1147);
    not g1774(n2138 ,n2137);
    nand g1775(n2656 ,n2611 ,n2631);
    nand g1776(n490 ,n6[0] ,n462);
    nand g1777(n1719 ,n20[7] ,n22[1]);
    nor g1778(n112 ,n26[14] ,n26[15]);
    nand g1779(n2610 ,n2702 ,n2547);
    nand g1780(n852 ,n2720 ,n825);
    nand g1781(n1607 ,n20[6] ,n22[4]);
    xnor g1782(n2699 ,n1112 ,n1107);
    nand g1783(n289 ,n29[14] ,n141);
    nand g1784(n711 ,n578 ,n529);
    nor g1785(n177 ,n152 ,n149);
    nand g1786(n1672 ,n21[3] ,n23[1]);
    nand g1787(n930 ,n845 ,n909);
    xnor g1788(n2250 ,n2144 ,n2184);
    or g1789(n2228 ,n2168 ,n2195);
    xnor g1790(n1139 ,n1095 ,n1097);
    xnor g1791(n135 ,n19[7] ,n28[7]);
    nand g1792(n1283 ,n2675 ,n23[3]);
    nand g1793(n1899 ,n1609 ,n1787);
    nor g1794(n1445 ,n1379 ,n1432);
    not g1795(n1568 ,n23[7]);
    nand g1796(n1598 ,n20[0] ,n22[3]);
    nor g1797(n723 ,n633 ,n668);
    nor g1798(n1158 ,n1059 ,n1119);
    not g1799(n1659 ,n1658);
    nor g1800(n99 ,n5[15] ,n5[14]);
    dff g1801(.RN(n1), .SN(1'b1), .CK(n0), .D(n426), .Q(n10[4]));
    nand g1802(n1954 ,n1737 ,n1890);
    nand g1803(n1550 ,n1527 ,n1546);
    nand g1804(n2443 ,n22[2] ,n23[2]);
    or g1805(n1729 ,n1581 ,n1650);
    buf g1806(n11[10], 1'b0);
    dff g1807(.RN(n1), .SN(1'b1), .CK(n0), .D(n378), .Q(n28[3]));
    buf g1808(n12[23], n10[15]);
    dff g1809(.RN(n1), .SN(1'b1), .CK(n0), .D(n473), .Q(n16));
    nand g1810(n1871 ,n1658 ,n1810);
    not g1811(n1972 ,n1971);
    nand g1812(n679 ,n612 ,n611);
    nand g1813(n2549 ,n2731 ,n32[2]);
    nand g1814(n284 ,n31[0] ,n141);
    nand g1815(n360 ,n15 ,n345);
    nand g1816(n944 ,n841 ,n897);
    xnor g1817(n129 ,n19[1] ,n28[1]);
    nand g1818(n538 ,n21[1] ,n463);
    xnor g1819(n2382 ,n2323 ,n2343);
    or g1820(n2311 ,n2272 ,n2284);
    nor g1821(n2161 ,n2072 ,n2106);
    xnor g1822(n1137 ,n1074 ,n1109);
    or g1823(n1128 ,n1094 ,n1097);
    nand g1824(n324 ,n10[5] ,n156);
    buf g1825(n9[15], 1'b0);
    nor g1826(n1025 ,n1022 ,n997);
    nand g1827(n2322 ,n2265 ,n2288);
    nor g1828(n847 ,n812 ,n819);
    nand g1829(n235 ,n31[14] ,n155);
    nand g1830(n424 ,n323 ,n241);
    nand g1831(n741 ,n35 ,n39);
    nand g1832(n2529 ,n2478 ,n2528);
    not g1833(n1431 ,n1423);
    nand g1834(n2618 ,n2699 ,n2547);
    not g1835(n88 ,n5[3]);
    nand g1836(n2576 ,n32[6] ,n2561);
    nand g1837(n598 ,n19[6] ,n481);
    nor g1838(n1389 ,n1295 ,n1352);
    xor g1839(n2299 ,n2269 ,n2247);
    nor g1840(n1398 ,n1325 ,n1334);
    buf g1841(n13[13], 1'b0);
    nand g1842(n694 ,n566 ,n519);
    nand g1843(n1875 ,n1635 ,n1769);
    nand g1844(n573 ,n22[7] ,n478);
    xnor g1845(n2690 ,n2421 ,n2426);
    nand g1846(n2004 ,n1764 ,n1920);
    nand g1847(n1616 ,n20[5] ,n22[0]);
    dff g1848(.RN(n1), .SN(1'b1), .CK(n0), .D(n387), .Q(n26[13]));
    nand g1849(n656 ,n548 ,n506);
    nor g1850(n2563 ,n2560 ,n2536);
    nand g1851(n453 ,n155 ,n449);
    buf g1852(n11[13], 1'b0);
    nand g1853(n647 ,n541 ,n501);
    dff g1854(.RN(n1), .SN(1'b1), .CK(n0), .D(n653), .Q(n20[1]));
    nand g1855(n536 ,n21[3] ,n463);
    nor g1856(n1316 ,n1266 ,n1283);
    nand g1857(n2005 ,n1657 ,n1945);
    nand g1858(n1916 ,n1738 ,n1905);
    nand g1859(n2649 ,n2602 ,n2621);
    nand g1860(n673 ,n602 ,n601);
    nand g1861(n1773 ,n1679 ,n1688);
    dff g1862(.RN(n1), .SN(1'b1), .CK(n0), .D(n659), .Q(n19[4]));
    nand g1863(n483 ,n6[1] ,n464);
    xnor g1864(n2134 ,n2031 ,n1920);
    nor g1865(n2168 ,n2055 ,n2111);
    buf g1866(n9[26], 1'b0);
    nand g1867(n516 ,n6[3] ,n462);
    xnor g1868(n2254 ,n2135 ,n2186);
    nand g1869(n1804 ,n1599 ,n1590);
    xnor g1870(n1470 ,n1437 ,n1264);
    nand g1871(n251 ,n29[10] ,n140);
    nand g1872(n1924 ,n1736 ,n1879);
    not g1873(n1104 ,n1103);
    nor g1874(n47 ,n25[1] ,n25[0]);
    buf g1875(n13[14], 1'b0);
    xnor g1876(n2052 ,n1823 ,n1956);
    xnor g1877(n2139 ,n2032 ,n1930);
    nand g1878(n2098 ,n1924 ,n2038);
    or g1879(n1731 ,n1661 ,n1693);
    or g1880(n1758 ,n1679 ,n1688);
    xnor g1881(n743 ,n25[6] ,n75);
    nand g1882(n421 ,n9[4] ,n252);
    nor g1883(n1288 ,n1266 ,n1281);
    not g1884(n1259 ,n1258);
    nand g1885(n2639 ,n2597 ,n2616);
    nor g1886(n48 ,n25[3] ,n25[2]);
    xnor g1887(n2184 ,n2087 ,n1988);
    nand g1888(n2019 ,n1869 ,n1931);
    nor g1889(n2509 ,n2471 ,n2508);
    nor g1890(n1327 ,n1267 ,n1281);
    xnor g1891(n1991 ,n1845 ,n1617);
    nand g1892(n1144 ,n1075 ,n1120);
    nand g1893(n641 ,n535 ,n497);
    nand g1894(n532 ,n6[0] ,n470);
    nand g1895(n2623 ,n2574 ,n2573);
    or g1896(n1056 ,n931 ,n990);
    nand g1897(n660 ,n552 ,n510);
    nor g1898(n1914 ,n1806 ,n1855);
    xnor g1899(n1508 ,n1265 ,n1475);
    xnor g1900(n1486 ,n1455 ,n1453);
    nand g1901(n645 ,n539 ,n484);
    nand g1902(n2553 ,n2728 ,n32[5]);
    xnor g1903(n983 ,n944 ,n816);
    or g1904(n2060 ,n2014 ,n2016);
    buf g1905(n17[6], 1'b0);
    nor g1906(n1391 ,n1317 ,n1351);
    xnor g1907(n2454 ,n23[3] ,n22[3]);
    not g1908(n1172 ,n1171);
    xnor g1909(n999 ,n926 ,n818);
    buf g1910(n12[31], 1'b0);
    nor g1911(n125 ,n26[8] ,n26[9]);
    nand g1912(n587 ,n21[7] ,n467);
    nand g1913(n1046 ,n994 ,n989);
    not g1914(n1981 ,n1980);
    nand g1915(n868 ,n2714 ,n824);
    or g1916(n1748 ,n1678 ,n1694);
    not g1917(n638 ,n622);
    nand g1918(n1620 ,n21[5] ,n23[1]);
    nand g1919(n1462 ,n1389 ,n1441);
    nor g1920(n1385 ,n1327 ,n1364);
    nand g1921(n65 ,n30[6] ,n64);
    not g1922(n2163 ,n2162);
    nand g1923(n1792 ,n1583 ,n1681);
    nand g1924(n828 ,n2718 ,n821);
    nand g1925(n579 ,n22[1] ,n478);
    dff g1926(.RN(n1), .SN(1'b1), .CK(n0), .D(n700), .Q(n23[2]));
    nor g1927(n480 ,n252 ,n460);
    or g1928(n457 ,n166 ,n78);
    xnor g1929(n823 ,n807 ,n786);
    nor g1930(n2474 ,n2706 ,n2690);
    or g1931(n2040 ,n1918 ,n1965);
    xnor g1932(n986 ,n923 ,n818);
    nor g1933(n715 ,n655 ,n704);
    nor g1934(n1083 ,n935 ,n1053);
    xnor g1935(n1994 ,n1854 ,n1806);
    nor g1936(n848 ,n813 ,n820);
    nor g1937(n1080 ,n999 ,n1041);
    dff g1938(.RN(n1), .SN(1'b1), .CK(n0), .D(n436), .Q(n30[2]));
    nand g1939(n1669 ,n21[2] ,n23[1]);
    nor g1940(n1132 ,n1038 ,n1105);
    not g1941(n1815 ,n1800);
    nor g1942(n467 ,n252 ,n456);
    xnor g1943(n961 ,n806 ,n903);
    nand g1944(n2648 ,n2555 ,n2570);
    nand g1945(n668 ,n397 ,n590);
    buf g1946(n11[26], n10[10]);
    nand g1947(n678 ,n402 ,n597);
    xnor g1948(n1828 ,n1597 ,n1669);
    buf g1949(n13[21], 1'b0);
    nor g1950(n1333 ,n1267 ,n1282);
    buf g1951(n13[20], 1'b0);
    nand g1952(n2069 ,n1968 ,n1961);
    or g1953(n31[7] ,n2635 ,n2656);
    nand g1954(n2640 ,n2552 ,n2567);
    dff g1955(.RN(n1), .SN(1'b1), .CK(n0), .D(n417), .Q(n10[12]));
    nand g1956(n2619 ,n2705 ,n2547);
    nand g1957(n2369 ,n2320 ,n2346);
    nor g1958(n1055 ,n934 ,n1013);
    nand g1959(n318 ,n10[10] ,n156);
    buf g1960(n17[0], n17[2]);
    xnor g1961(n2453 ,n22[2] ,n23[2]);
    nand g1962(n841 ,n2718 ,n819);
    nand g1963(n611 ,n22[3] ,n469);
    or g1964(n2406 ,n2398 ,n2381);
    nand g1965(n945 ,n874 ,n885);
    not g1966(n1706 ,n1705);
    xnor g1967(n936 ,n816 ,n827);
    nand g1968(n735 ,n727 ,n718);
    nor g1969(n2466 ,n2447 ,n2465);
    nand g1970(n913 ,n2717 ,n876);
    not g1971(n2169 ,n2155);
    nor g1972(n2211 ,n2058 ,n2169);
    nor g1973(n1079 ,n995 ,n1039);
    nand g1974(n1415 ,n1394 ,n1391);
    nand g1975(n2626 ,n2606 ,n2588);
    xnor g1976(n2695 ,n2339 ,n2436);
    nand g1977(n2585 ,n32[11] ,n2561);
    nand g1978(n798 ,n777 ,n772);
    xor g1979(n2674 ,n20[2] ,n21[2]);
    nand g1980(n2587 ,n2681 ,n2546);
    nand g1981(n615 ,n20[3] ,n468);
    nand g1982(n667 ,n589 ,n588);
    nand g1983(n1937 ,n1760 ,n1906);
    or g1984(n2333 ,n2268 ,n2301);
    xnor g1985(n137 ,n19[2] ,n28[2]);
    nor g1986(n104 ,n26[10] ,n26[11]);
    nand g1987(n685 ,n617 ,n618);
    xnor g1988(n1841 ,n1603 ,n1665);
    nand g1989(n888 ,n2714 ,n846);
    xnor g1990(n2380 ,n2345 ,n2318);
    nand g1991(n1926 ,n1759 ,n1889);
    xnor g1992(n1960 ,n1864 ,n1585);
    nor g1993(n1319 ,n1266 ,n1279);
    nand g1994(n2661 ,n2618 ,n2645);
    nand g1995(n317 ,n10[11] ,n156);
    xnor g1996(n2020 ,n1821 ,n1861);
    not g1997(n2446 ,n2445);
    nand g1998(n2631 ,n2550 ,n2563);
    not g1999(n91 ,n5[4]);
    not g2000(n1248 ,n1247);
    nor g2001(n2290 ,n2233 ,n2262);
    nand g2002(n313 ,n10[15] ,n156);
    nand g2003(n937 ,n828 ,n913);
    nand g2004(n322 ,n31[15] ,n141);
    nor g2005(n2516 ,n2486 ,n2515);
    nand g2006(n697 ,n568 ,n521);
    nand g2007(n580 ,n22[0] ,n478);
    not g2008(n1810 ,n1809);
    dff g2009(.RN(n1), .SN(1'b1), .CK(n0), .D(n411), .Q(n25[2]));
    nand g2010(n1713 ,n20[4] ,n22[7]);
    not g2011(n1099 ,n1098);
    nor g2012(n110 ,n5[17] ,n5[16]);
    nand g2013(n2225 ,n2136 ,n2186);
    or g2014(n1737 ,n1583 ,n1681);
    nor g2015(n766 ,n20[3] ,n21[3]);
    nor g2016(n1037 ,n965 ,n1008);
    or g2017(n2314 ,n2211 ,n2281);
    xnor g2018(n2345 ,n2296 ,n2307);
    nand g2019(n420 ,n319 ,n211);
    nand g2020(n2370 ,n2333 ,n2354);
    or g2021(n2391 ,n2349 ,n2382);
    nor g2022(n120 ,n26[12] ,n26[13]);
    nand g2023(n860 ,n2714 ,n825);
    nand g2024(n314 ,n10[14] ,n156);
    nand g2025(n767 ,n20[6] ,n20[5]);
    nand g2026(n323 ,n10[6] ,n156);
    nor g2027(n825 ,n783 ,n811);
    nand g2028(n2483 ,n2696 ,n2680);
    nand g2029(n501 ,n6[6] ,n466);
    or g2030(n182 ,n17[2] ,n155);
    nand g2031(n857 ,n2713 ,n825);
    nand g2032(n1178 ,n1121 ,n1145);
    nor g2033(n730 ,n670 ,n669);
    nand g2034(n256 ,n26[9] ,n87);
    nand g2035(n2118 ,n2018 ,n2063);
    buf g2036(n12[13], n10[5]);
    xnor g2037(n2726 ,n2502 ,n2511);
    nor g2038(n2166 ,n2075 ,n2107);
    nor g2039(n2385 ,n2365 ,n2364);
    xnor g2040(n1073 ,n968 ,n994);
    xnor g2041(n1243 ,n1219 ,n1231);
    nand g2042(n1868 ,n1586 ,n1765);
    nand g2043(n1110 ,n1056 ,n1084);
    nand g2044(n368 ,n228 ,n322);
    nand g2045(n1915 ,n1752 ,n1878);
    dff g2046(.RN(n1), .SN(1'b1), .CK(n0), .D(n641), .Q(n21[4]));
    nand g2047(n614 ,n23[3] ,n480);
    nand g2048(n1884 ,n1611 ,n1779);
    nand g2049(n2121 ,n2002 ,n2042);
    nand g2050(n594 ,n24[6] ,n482);
    nor g2051(n2269 ,n2203 ,n2235);
    not g2052(n1163 ,n1154);
    dff g2053(.RN(n1), .SN(1'b1), .CK(n0), .D(n441), .Q(n30[3]));
    nor g2054(n2058 ,n1968 ,n1961);
    nand g2055(n2625 ,n2605 ,n2604);
    nor g2056(n1357 ,n1269 ,n1296);
    not g2057(n1269 ,n24[1]);
    not g2058(n2493 ,n2492);
    nand g2059(n2601 ,n32[9] ,n2561);
    nand g2060(n336 ,n31[14] ,n141);
    dff g2061(.RN(n1), .SN(1'b1), .CK(n0), .D(n395), .Q(n30[5]));
    xnor g2062(n971 ,n806 ,n906);
    nand g2063(n485 ,n6[1] ,n466);
    nand g2064(n1776 ,n1598 ,n1593);
    nand g2065(n2061 ,n1944 ,n1963);
    nand g2066(n2636 ,n2551 ,n2565);
    nand g2067(n2276 ,n2194 ,n2240);
    nand g2068(n1481 ,n1419 ,n1465);
    nand g2069(n1715 ,n20[7] ,n22[2]);
    nor g2070(n1197 ,n1162 ,n1166);
    nor g2071(n795 ,n770 ,n774);
    nand g2072(n585 ,n21[0] ,n467);
    not g2073(n815 ,n816);
    not g2074(n962 ,n961);
    nor g2075(n2545 ,n2722 ,n32[11]);
    nand g2076(n2334 ,n2294 ,n2315);
    or g2077(n1495 ,n1447 ,n1471);
    not g2078(n1119 ,n1118);
    nand g2079(n1644 ,n21[2] ,n23[4]);
    buf g2080(n11[8], 1'b0);
    not g2081(n1147 ,n1146);
    nor g2082(n2571 ,n2560 ,n2543);
    xnor g2083(n1118 ,n1072 ,n1010);
    nand g2084(n1888 ,n1714 ,n1804);
    nand g2085(n870 ,n2720 ,n820);
    nand g2086(n1501 ,n1461 ,n1478);
    nand g2087(n542 ,n20[5] ,n465);
    nand g2088(n553 ,n19[2] ,n476);
    nor g2089(n1330 ,n1267 ,n1285);
    nor g2090(n2467 ,n2439 ,n2466);
    xor g2091(n2174 ,n2051 ,n2124);
    not g2092(n1306 ,n1307);
    nand g2093(n889 ,n2716 ,n847);
    nand g2094(n2043 ,n1938 ,n1982);
    nand g2095(n2240 ,n2124 ,n2206);
    or g2096(n1270 ,n2675 ,n23[3]);
    nand g2097(n2433 ,n2432 ,n2394);
    dff g2098(.RN(n1), .SN(1'b1), .CK(n0), .D(n440), .Q(n30[1]));
    nor g2099(n1344 ,n1266 ,n1305);
    nand g2100(n612 ,n21[3] ,n467);
    nand g2101(n2000 ,n1801 ,n1956);
    nand g2102(n874 ,n2719 ,n819);
    nand g2103(n209 ,n29[12] ,n87);
    nor g2104(n1244 ,n1194 ,n1234);
    nor g2105(n1341 ,n1267 ,n1301);
    nand g2106(n410 ,n254 ,n309);
    nand g2107(n2214 ,n2094 ,n2154);
    nand g2108(n277 ,n31[9] ,n141);
    nor g2109(n1090 ,n1005 ,n1057);
    not g2110(n465 ,n466);
    nand g2111(n473 ,n288 ,n453);
    nor g2112(n1764 ,n1716 ,n1626);
    nor g2113(n94 ,n7[2] ,n7[1]);
    nand g2114(n770 ,n20[0] ,n21[0]);
    nand g2115(n786 ,n2712 ,n783);
    nand g2116(n1161 ,n978 ,n1130);
    nand g2117(n1491 ,n1451 ,n1469);
    nand g2118(n229 ,n26[0] ,n87);
    dff g2119(.RN(n1), .SN(1'b1), .CK(n0), .D(n385), .Q(n26[15]));
    nand g2120(n2583 ,n2691 ,n2546);
    xnor g2121(n1141 ,n756 ,n1105);
    nand g2122(n2558 ,n2726 ,n32[7]);
    nand g2123(n344 ,n2 ,n144);
    not g2124(n2489 ,n2488);
    xnor g2125(n1967 ,n1844 ,n1708);
    nand g2126(n571 ,n23[1] ,n474);
    xnor g2127(n1242 ,n1225 ,n1200);
    nor g2128(n1459 ,n1407 ,n1446);
    nand g2129(n1695 ,n20[1] ,n22[7]);
    nand g2130(n1922 ,n1732 ,n1874);
    nand g2131(n56 ,n30[1] ,n30[0]);
    xnor g2132(n1965 ,n1817 ,n1629);
    nor g2133(n1881 ,n1612 ,n1815);
    nand g2134(n2505 ,n2470 ,n2504);
    nor g2135(n744 ,n74 ,n76);
    nand g2136(n2274 ,n2176 ,n2238);
    nand g2137(n794 ,n2719 ,n783);
    not g2138(n1220 ,n1219);
    xnor g2139(n2683 ,n2252 ,n2246);
    dff g2140(.RN(n1), .SN(1'b1), .CK(n0), .D(n408), .Q(n25[5]));
    nand g2141(n217 ,n26[12] ,n87);
    nand g2142(n849 ,n2712 ,n821);
    nand g2143(n509 ,n6[4] ,n477);
    nand g2144(n1636 ,n20[4] ,n22[0]);
    nand g2145(n706 ,n437 ,n629);
    nand g2146(n1684 ,n21[5] ,n23[6]);
    not g2147(n1712 ,n1711);
    xnor g2148(n2286 ,n2220 ,n2164);
    nand g2149(n396 ,n223 ,n296);
    or g2150(n1998 ,n1764 ,n1920);
    nor g2151(n1131 ,n974 ,n1100);
    xnor g2152(n2691 ,n2419 ,n2428);
    nand g2153(n1512 ,n1484 ,n1498);
    or g2154(n1756 ,n1682 ,n1579);
    xnor g2155(n1992 ,n1847 ,n1687);
    xor g2156(n1264 ,n1377 ,n1367);
    nand g2157(n2440 ,n22[0] ,n23[0]);
    nand g2158(n459 ,n84 ,n80);
    nor g2159(n2221 ,n2160 ,n2190);
    nand g2160(n2595 ,n32[3] ,n2561);
    nand g2161(n2387 ,n2353 ,n2369);
    nor g2162(n729 ,n667 ,n666);
    nand g2163(n2573 ,n32[5] ,n2561);
    buf g2164(n9[23], 1'b0);
    dff g2165(.RN(n1), .SN(1'b1), .CK(n0), .D(n432), .Q(n30[6]));
    nand g2166(n2418 ,n2391 ,n2409);
    or g2167(n977 ,n932 ,n930);
    dff g2168(.RN(n1), .SN(1'b1), .CK(n0), .D(n642), .Q(n21[3]));
    not g2169(n1458 ,n1457);
    xnor g2170(n1977 ,n1831 ,n1612);
    nand g2171(n832 ,n2715 ,n819);
    nand g2172(n922 ,n842 ,n880);
    xnor g2173(n1401 ,n1361 ,n1329);
    nor g2174(n109 ,n5[19] ,n5[18]);
    not g2175(n2142 ,n2141);
    buf g2176(n12[17], n10[9]);
    xnor g2177(n1471 ,n1438 ,n1450);
    xnor g2178(n1089 ,n1021 ,n997);
    xor g2179(n2087 ,n1976 ,n2022);
    buf g2180(n9[27], 1'b0);
    nand g2181(n908 ,n2720 ,n846);
    nand g2182(n692 ,n564 ,n490);
    nand g2183(n2108 ,n1925 ,n2061);
    xnor g2184(n1963 ,n1838 ,n1596);
    nand g2185(n642 ,n536 ,n498);
    nor g2186(n1159 ,n1096 ,n1117);
    buf g2187(n10[29], 1'b0);
    nand g2188(n2609 ,n2706 ,n2547);
    nand g2189(n2065 ,n1978 ,n1977);
    xnor g2190(n776 ,n20[2] ,n21[2]);
    xor g2191(n1846 ,n1622 ,n1576);
    xnor g2192(n1074 ,n1002 ,n1013);
    or g2193(n168 ,n87 ,n132);
    not g2194(n1618 ,n1617);
    nand g2195(n2480 ,n2708 ,n2692);
    not g2196(n1429 ,n1421);
    xnor g2197(n2285 ,n2219 ,n2137);
    buf g2198(n11[25], n10[9]);
    nand g2199(n1882 ,n1712 ,n1770);
    or g2200(n1275 ,n2678 ,n23[6]);
    nand g2201(n595 ,n24[6] ,n461);
    nand g2202(n1671 ,n20[4] ,n22[2]);
    xnor g2203(n2449 ,n23[1] ,n22[1]);
    nand g2204(n561 ,n24[3] ,n461);
    buf g2205(n11[22], n10[6]);
    nand g2206(n864 ,n2717 ,n824);
    nand g2207(n2120 ,n2001 ,n2059);
    xnor g2208(n1845 ,n1670 ,n1674);
    nor g2209(n2680 ,n1814 ,n1761);
    nand g2210(n2525 ,n2477 ,n2524);
    nand g2211(n2593 ,n2701 ,n2547);
    nand g2212(n1650 ,n21[6] ,n23[3]);
    or g2213(n1997 ,n1915 ,n1916);
    nand g2214(n157 ,n99 ,n114);
    xnor g2215(n746 ,n25[3] ,n70);
    nand g2216(n58 ,n30[2] ,n57);
    dff g2217(.RN(n1), .SN(1'b1), .CK(n0), .D(n452), .Q(n18[0]));
    nand g2218(n731 ,n723 ,n729);
    nand g2219(n2373 ,n2330 ,n2355);
    nor g2220(n95 ,n5[9] ,n5[8]);
    xnor g2221(n2086 ,n1989 ,n1594);
    xnor g2222(n958 ,n901 ,n807);
    nor g2223(n1251 ,n1218 ,n1250);
    nand g2224(n189 ,n28[9] ,n87);
    xnor g2225(n996 ,n943 ,n818);
    nand g2226(n739 ,n49 ,n53);
    nand g2227(n713 ,n579 ,n493);
    nor g2228(n2521 ,n2476 ,n2520);
    nand g2229(n527 ,n6[4] ,n479);
    buf g2230(n12[25], 1'b0);
    xnor g2231(n2340 ,n2271 ,n2306);
    or g2232(n166 ,n146 ,n158);
    xnor g2233(n1537 ,n1493 ,n1525);
    nor g2234(n2197 ,n2121 ,n2143);
    nor g2235(n1239 ,n1211 ,n1227);
    nand g2236(n1951 ,n1748 ,n1893);
    nor g2237(n2475 ,n2701 ,n2685);
    nand g2238(n454 ,n83 ,n79);
    nand g2239(n1670 ,n20[2] ,n22[7]);
    nand g2240(n492 ,n6[0] ,n475);
    nand g2241(n2464 ,n2452 ,n2463);
    xnor g2242(n959 ,n806 ,n905);
    xnor g2243(n1233 ,n1188 ,n1212);
    nand g2244(n320 ,n10[8] ,n156);
    not g2245(n1975 ,n1974);
    nand g2246(n2481 ,n2698 ,n2682);
    nor g2247(n73 ,n66 ,n72);
    buf g2248(n11[20], n10[4]);
    nor g2249(n2561 ,n2532 ,n27[0]);
    nand g2250(n1685 ,n20[3] ,n22[4]);
    nand g2251(n342 ,n751 ,n141);
    nand g2252(n438 ,n197 ,n336);
    xor g2253(n1565 ,n1959 ,n1950);
    nor g2254(n477 ,n344 ,n457);
    nand g2255(n2432 ,n2408 ,n2431);
    xnor g2256(n1516 ,n1486 ,n1476);
    nor g2257(n1428 ,n1347 ,n1400);
    nand g2258(n1285 ,n2679 ,n23[7]);
    nand g2259(n2063 ,n1969 ,n1967);
    nor g2260(n846 ,n814 ,n824);
    nor g2261(n1033 ,n958 ,n1012);
    nand g2262(n790 ,n2718 ,n783);
    nor g2263(n2112 ,n1990 ,n2081);
    xnor g2264(n2033 ,n1656 ,n1945);
    nand g2265(n2424 ,n2423 ,n2407);
    nor g2266(n1395 ,n1291 ,n1355);
    nand g2267(n162 ,n94 ,n105);
    not g2268(n850 ,n849);
    nand g2269(n903 ,n788 ,n858);
    nand g2270(n326 ,n10[3] ,n156);
    nand g2271(n329 ,n10[0] ,n156);
    nor g2272(n43 ,n30[1] ,n41);
    xnor g2273(n2100 ,n1960 ,n1765);
    nand g2274(n286 ,n17[4] ,n156);
    nand g2275(n2647 ,n2596 ,n2595);
    or g2276(n2458 ,n2453 ,n2457);
    not g2277(n2182 ,n2181);
    xnor g2278(n1856 ,n1701 ,n1615);
    nor g2279(n2508 ,n2499 ,n2507);
    nor g2280(n1387 ,n1311 ,n1365);
    buf g2281(n11[1], 1'b0);
    not g2282(n1123 ,n1122);
    dff g2283(.RN(n1), .SN(1'b1), .CK(n0), .D(n367), .Q(n28[12]));
    buf g2284(n10[28], 1'b0);
    nor g2285(n105 ,n7[3] ,n7[0]);
    xnor g2286(n985 ,n925 ,n816);
    xnor g2287(n2301 ,n2248 ,n2230);
    nand g2288(n201 ,n29[0] ,n140);
    nand g2289(n2272 ,n2210 ,n2237);
    xnor g2290(n1206 ,n1173 ,n1138);
    nand g2291(n926 ,n840 ,n877);
    nor g2292(n1412 ,n1385 ,n1378);
    nand g2293(n829 ,n2714 ,n820);
    xnor g2294(n2420 ,n2396 ,n1566);
    nor g2295(n133 ,n127 ,n108);
    xnor g2296(n1019 ,n817 ,n953);
    nand g2297(n332 ,n31[6] ,n141);
    nand g2298(n842 ,n2716 ,n819);
    dff g2299(.RN(n1), .SN(1'b1), .CK(n0), .D(n393), .Q(n25[0]));
    nand g2300(n429 ,n9[3] ,n252);
    xnor g2301(n1450 ,n1331 ,n1398);
    or g2302(n1730 ,n1692 ,n1587);
    not g2303(n2148 ,n2147);
    nand g2304(n2179 ,n2101 ,n2131);
    buf g2305(n9[16], 1'b0);
    nand g2306(n895 ,n2718 ,n848);
    nand g2307(n657 ,n549 ,n507);
    nand g2308(n662 ,n553 ,n511);
    nand g2309(n498 ,n6[3] ,n464);
    or g2310(n1276 ,n2673 ,n23[1]);
    nand g2311(n2047 ,n1910 ,n2006);
    nand g2312(n1770 ,n1574 ,n1683);
    or g2313(n1909 ,n1691 ,n1860);
    nand g2314(n1689 ,n20[7] ,n22[7]);
    not g2315(n1192 ,n1191);
    dff g2316(.RN(n1), .SN(1'b1), .CK(n0), .D(n412), .Q(n25[1]));
    nand g2317(n117 ,n18[1] ,n93);
    nor g2318(n1417 ,n1326 ,n1397);
    xnor g2319(n753 ,n30[3] ,n58);
    nand g2320(n1878 ,n1622 ,n1802);
    nand g2321(n455 ,n84 ,n451);
    nor g2322(n1384 ,n1329 ,n1362);
    buf g2323(n10[18], 1'b0);
    xnor g2324(n1863 ,n1647 ,n1715);
    nand g2325(n1466 ,n1415 ,n1450);
    nand g2326(n655 ,n583 ,n582);
    nor g2327(n2077 ,n1942 ,n1981);
    nor g2328(n1371 ,n1322 ,n1345);
    xnor g2329(n1518 ,n1500 ,n1330);
    dff g2330(.RN(n1), .SN(1'b1), .CK(n0), .D(n420), .Q(n10[9]));
    nand g2331(n734 ,n724 ,n730);
    xnor g2332(n1493 ,n1440 ,n1460);
    nand g2333(n495 ,n6[6] ,n464);
    nand g2334(n2434 ,n2399 ,n2433);
    nand g2335(n2124 ,n2003 ,n2039);
    nand g2336(n617 ,n21[2] ,n467);
    nor g2337(n1392 ,n1294 ,n1337);
    nand g2338(n855 ,n2718 ,n825);
    xnor g2339(n742 ,n25[7] ,n77);
    xnor g2340(n2698 ,n1071 ,n1017);
    nand g2341(n1956 ,n1755 ,n1897);
    nand g2342(n1560 ,n1534 ,n1559);
    nand g2343(n510 ,n6[3] ,n477);
    or g2344(n2360 ,n2305 ,n2344);
    nand g2345(n399 ,n225 ,n298);
    nand g2346(n1654 ,n21[7] ,n23[7]);
    buf g2347(n13[17], 1'b0);
    nand g2348(n215 ,n25[4] ,n142);
    xnor g2349(n1474 ,n1439 ,n1399);
    nand g2350(n205 ,n28[4] ,n87);
    dff g2351(.RN(n1), .SN(1'b1), .CK(n0), .D(n356), .Q(n29[0]));
    nor g2352(n1743 ,n1663 ,n1662);
    xnor g2353(n1146 ,n982 ,n1111);
    nand g2354(n737 ,n721 ,n720);
    xor g2355(n2730 ,n2492 ,n2483);
    nor g2356(n1379 ,n1292 ,n1338);
    buf g2357(n13[9], 1'b0);
    xnor g2358(n777 ,n20[4] ,n21[4]);
    nor g2359(n834 ,n758 ,n822);
    nand g2360(n2425 ,n2414 ,n2424);
    not g2361(n1149 ,n1148);
    nand g2362(n1556 ,n1540 ,n1555);
    xnor g2363(n1241 ,n1226 ,n1211);
    xnor g2364(n1097 ,n1026 ,n990);
    nand g2365(n2289 ,n2213 ,n2257);
    xnor g2366(n2671 ,n2484 ,n2531);
    nand g2367(n2279 ,n2224 ,n2273);
    nor g2368(n2510 ,n2500 ,n2509);
    nand g2369(n502 ,n6[5] ,n466);
    buf g2370(n11[2], 1'b0);
    xnor g2371(n1115 ,n1063 ,n983);
    nor g2372(n724 ,n634 ,n671);
    nor g2373(n35 ,n30[6] ,n30[5]);
    nand g2374(n808 ,n775 ,n801);
    xnor g2375(n1165 ,n1119 ,n1058);
    xor g2376(n2731 ,n2696 ,n2680);
    nor g2377(n2543 ,n2726 ,n32[7]);
    nand g2378(n499 ,n6[2] ,n464);
    xnor g2379(n1003 ,n928 ,n807);
    xnor g2380(n132 ,n19[3] ,n28[3]);
    nand g2381(n283 ,n31[1] ,n141);
    nand g2382(n1600 ,n21[2] ,n23[2]);
    nor g2383(n1219 ,n1182 ,n1196);
    buf g2384(n9[21], 1'b0);
    xnor g2385(n2186 ,n2088 ,n2019);
    nor g2386(n2562 ,n2560 ,n2535);
    nand g2387(n387 ,n216 ,n290);
    nand g2388(n866 ,n2716 ,n824);
    nand g2389(n436 ,n203 ,n340);
    nand g2390(n1151 ,n1110 ,n1129);
    nand g2391(n2461 ,n2442 ,n2460);
    nor g2392(n1418 ,n1308 ,n1393);
    or g2393(n174 ,n140 ,n129);
    nor g2394(n185 ,n160 ,n163);
    dff g2395(.RN(n1), .SN(1'b1), .CK(n0), .D(n390), .Q(n26[10]));
    nand g2396(n2607 ,n2710 ,n2547);
    not g2397(n93 ,n18[0]);
    dff g2398(.RN(n1), .SN(1'b1), .CK(n0), .D(n439), .Q(n30[4]));
    nand g2399(n836 ,n2716 ,n820);
    not g2400(n1703 ,n1702);
    nand g2401(n925 ,n838 ,n889);
    nand g2402(n2268 ,n2177 ,n2239);
    nand g2403(n2164 ,n2060 ,n2116);
    nand g2404(n2316 ,n2272 ,n2284);
    nand g2405(n1044 ,n1007 ,n993);
    nand g2406(n1634 ,n21[1] ,n23[2]);
    xnor g2407(n2501 ,n2706 ,n2690);
    xnor g2408(n2488 ,n2708 ,n2692);
    buf g2409(n9[30], 1'b0);
    nand g2410(n2550 ,n2724 ,n32[9]);
    nand g2411(n341 ,n749 ,n141);
    nand g2412(n1901 ,n1645 ,n1795);
    nand g2413(n1716 ,n20[2] ,n22[1]);
    xnor g2414(n2687 ,n2402 ,n2409);
    xnor g2415(n1070 ,n991 ,n986);
    nand g2416(n1175 ,n1161 ,n1126);
    xnor g2417(n1834 ,n1583 ,n1681);
    nor g2418(n1488 ,n1457 ,n1473);
    nand g2419(n1017 ,n851 ,n969);
    nand g2420(n2312 ,n2231 ,n2286);
    buf g2421(n12[24], 1'b0);
    not g2422(n1986 ,n1985);
    xnor g2423(n1002 ,n935 ,n933);
    nor g2424(n2537 ,n2731 ,n32[2]);
    nand g2425(n426 ,n325 ,n243);
    nand g2426(n433 ,n250 ,n333);
    xnor g2427(n2379 ,n2319 ,n2346);
    dff g2428(.RN(n1), .SN(1'b1), .CK(n0), .D(n376), .Q(n28[5]));
    nor g2429(n2540 ,n2723 ,n32[10]);
    nand g2430(n949 ,n864 ,n890);
    xnor g2431(n2486 ,n2703 ,n2687);
    or g2432(n1048 ,n986 ,n991);
    buf g2433(n10[24], 1'b0);
    nor g2434(n2476 ,n2705 ,n2689);
    nand g2435(n1913 ,n1762 ,n1859);
    nand g2436(n1945 ,n1727 ,n1882);
    nor g2437(n1031 ,n817 ,n992);
    nor g2438(n1255 ,n1240 ,n1254);
    nand g2439(n1523 ,n1487 ,n1513);
    nand g2440(n933 ,n843 ,n915);
    nand g2441(n809 ,n785 ,n800);
    xnor g2442(n1973 ,n1841 ,n1640);
    not g2443(n145 ,n144);
    xnor g2444(n32[8] ,n1548 ,n1555);
    xnor g2445(n2026 ,n1941 ,n1953);
    xnor g2446(n2258 ,n2171 ,n2049);
    nand g2447(n203 ,n30[2] ,n140);
    not g2448(n1570 ,n23[4]);
    nand g2449(n844 ,n2715 ,n820);
    xnor g2450(n989 ,n945 ,n816);
    nand g2451(n2462 ,n2446 ,n2461);
    xnor g2452(n2216 ,n2134 ,n2048);
    xnor g2453(n2175 ,n2100 ,n2123);
    nand g2454(n159 ,n86 ,n96);
    nor g2455(n1944 ,n1745 ,n1877);
    dff g2456(.RN(n1), .SN(1'b1), .CK(n0), .D(n424), .Q(n10[6]));
    nand g2457(n2614 ,n2697 ,n2547);
    nor g2458(n1806 ,n1710 ,n1698);
    nand g2459(n199 ,n28[12] ,n140);
    nand g2460(n624 ,n23[1] ,n480);
    not g2461(n1814 ,n1797);
    nand g2462(n295 ,n29[7] ,n141);
    nand g2463(n2110 ,n2015 ,n2047);
    nand g2464(n665 ,n555 ,n531);
    xnor g2465(n1189 ,n1137 ,n1120);
    xnor g2466(n1231 ,n1184 ,n1162);
    xnor g2467(n992 ,n947 ,n816);
    xor g2468(n2677 ,n20[5] ,n21[5]);
    nand g2469(n541 ,n20[6] ,n465);
    nand g2470(n1536 ,n1493 ,n1525);
    xnor g2471(n2231 ,n2127 ,n2079);
    nor g2472(n462 ,n344 ,n458);
    xnor g2473(n804 ,n760 ,n778);
    nand g2474(n600 ,n21[5] ,n467);
    nor g2475(n2055 ,n1973 ,n1970);
    nand g2476(n261 ,n29[5] ,n87);
    nand g2477(n2605 ,n2692 ,n2546);
    nand g2478(n1447 ,n1369 ,n1410);
    nand g2479(n1559 ,n1541 ,n1558);
    xnor g2480(n1980 ,n1836 ,n1610);
    nand g2481(n1596 ,n20[3] ,n22[7]);
    nand g2482(n942 ,n839 ,n893);
    xnor g2483(n2381 ,n2341 ,n2344);
    nand g2484(n780 ,n21[6] ,n765);
    nand g2485(n826 ,n2712 ,n820);
    not g2486(n1469 ,n1468);
    nand g2487(n608 ,n23[4] ,n480);
    not g2488(n2140 ,n2139);
    nor g2489(n1507 ,n1459 ,n1488);
    nand g2490(n2327 ,n2260 ,n2303);
    nor g2491(n1325 ,n1266 ,n1284);
    buf g2492(n13[27], n10[3]);
    xnor g2493(n2421 ,n2404 ,n2393);
    nand g2494(n830 ,n2716 ,n821);
    nor g2495(n1374 ,n1315 ,n1353);
    nor g2496(n1515 ,n1479 ,n1494);
    xnor g2497(n1502 ,n1468 ,n1451);
    nand g2498(n2431 ,n2430 ,n2405);
    nand g2499(n2198 ,n2099 ,n2133);
    buf g2500(n11[21], n10[5]);
    nand g2501(n932 ,n830 ,n911);
    or g2502(n2357 ,n2285 ,n2343);
    nand g2503(n373 ,n202 ,n272);
    nand g2504(n1561 ,n1536 ,n1560);
    or g2505(n1461 ,n1389 ,n1441);
    nand g2506(n1923 ,n1729 ,n1884);
    dff g2507(.RN(n1), .SN(1'b1), .CK(n0), .D(n389), .Q(n26[11]));
    nor g2508(n1133 ,n976 ,n1108);
    nand g2509(n524 ,n6[7] ,n479);
    nand g2510(n592 ,n22[6] ,n469);
    nor g2511(n100 ,n5[23] ,n5[22]);
    nor g2512(n1331 ,n1267 ,n1279);
    nand g2513(n2207 ,n1966 ,n2132);
    xnor g2514(n2188 ,n2089 ,n1980);
    nor g2515(n1156 ,n1033 ,n1124);
    not g2516(n1454 ,n1453);
    nand g2517(n288 ,n16 ,n156);
    xnor g2518(n1145 ,n1001 ,n1100);
    buf g2519(n13[26], n10[2]);
    nand g2520(n497 ,n6[4] ,n464);
    buf g2521(n12[29], 1'b0);
    nor g2522(n1036 ,n1006 ,n988);
    nand g2523(n44 ,n42 ,n43);
    nor g2524(n755 ,n57 ,n55);
    nand g2525(n2239 ,n2164 ,n2178);
    nor g2526(n1336 ,n1269 ,n1298);
    nand g2527(n557 ,n27[0] ,n471);
    nand g2528(n1584 ,n21[1] ,n23[6]);
    nand g2529(n1947 ,n1730 ,n1887);
    dff g2530(.RN(n1), .SN(1'b1), .CK(n0), .D(n366), .Q(n29[12]));
    nor g2531(n2538 ,n2730 ,n32[3]);
    nand g2532(n214 ,n26[14] ,n87);
    nand g2533(n616 ,n19[3] ,n481);
    nand g2534(n625 ,n27[1] ,n472);
    nor g2535(n2547 ,n27[1] ,n27[0]);
    nand g2536(n2417 ,n2397 ,n2403);
    dff g2537(.RN(n1), .SN(1'b1), .CK(n0), .D(n405), .Q(n26[0]));
    buf g2538(n13[29], n10[5]);
    nand g2539(n37 ,n30[4] ,n36);
    nand g2540(n1613 ,n20[4] ,n22[6]);
    dff g2541(.RN(n1), .SN(1'b1), .CK(n0), .D(n643), .Q(n21[2]));
    nand g2542(n1780 ,n1682 ,n1579);
    not g2543(n2559 ,n2560);
    nand g2544(n1880 ,n1721 ,n1772);
    nand g2545(n2074 ,n1936 ,n1986);
    buf g2546(n11[5], 1'b0);
    nand g2547(n238 ,n31[10] ,n155);
    nand g2548(n586 ,n22[7] ,n469);
    nand g2549(n839 ,n2713 ,n819);
    nand g2550(n278 ,n29[15] ,n141);
    nand g2551(n649 ,n543 ,n503);
    nand g2552(n2654 ,n2580 ,n2632);
    nand g2553(n2123 ,n2004 ,n2037);
    nand g2554(n299 ,n29[3] ,n141);
    xor g2555(n2672 ,n20[0] ,n21[0]);
    xor g2556(n1566 ,n2378 ,n2364);
    or g2557(n1753 ,n1689 ,n1654);
    nand g2558(n1531 ,n1514 ,n1516);
    xnor g2559(n2710 ,n1223 ,n1260);
    nand g2560(n696 ,n624 ,n623);
    nand g2561(n1680 ,n20[3] ,n22[2]);
    nor g2562(n2318 ,n2221 ,n2290);
    nor g2563(n1237 ,n1201 ,n1225);
    nand g2564(n231 ,n25[6] ,n142);
    nand g2565(n1687 ,n20[1] ,n22[6]);
    xnor g2566(n1854 ,n1716 ,n1626);
    nor g2567(n1214 ,n1179 ,n1193);
    nand g2568(n1681 ,n21[6] ,n23[6]);
    nand g2569(n1303 ,n1284 ,n1271);
    xnor g2570(n2500 ,n2700 ,n2684);
    buf g2571(n13[5], 1'b0);
    nand g2572(n1677 ,n21[2] ,n23[5]);
    not g2573(n1227 ,n1226);
    nand g2574(n378 ,n206 ,n282);
    or g2575(n31[9] ,n2650 ,n2660);
    nand g2576(n292 ,n29[11] ,n141);
    nand g2577(n543 ,n20[4] ,n465);
    nand g2578(n257 ,n29[9] ,n140);
    xnor g2579(n2419 ,n2403 ,n2397);
    nand g2580(n266 ,n30[5] ,n140);
    nor g2581(n1030 ,n961 ,n1010);
    nor g2582(n1204 ,n1158 ,n1174);
    nand g2583(n1305 ,n1280 ,n1276);
    nor g2584(n451 ,n136 ,n82);
    nor g2585(n975 ,n806 ,n928);
    or g2586(n1742 ,n1696 ,n1664);
    nand g2587(n2150 ,n2079 ,n2096);
    xnor g2588(n2089 ,n1991 ,n1942);
    nor g2589(n1136 ,n1051 ,n1102);
    xnor g2590(n2326 ,n2281 ,n2211);
    nand g2591(n411 ,n232 ,n310);
    nand g2592(n1674 ,n20[5] ,n22[4]);
    nand g2593(n2504 ,n2483 ,n2493);
    xnor g2594(n1067 ,n988 ,n1006);
    dff g2595(.RN(n1), .SN(1'b1), .CK(n0), .D(n401), .Q(n26[2]));
    xnor g2596(n1091 ,n1023 ,n972);
    xnor g2597(n2218 ,n2121 ,n2147);
    not g2598(n1328 ,n1327);
    nand g2599(n51 ,n25[4] ,n50);
    nand g2600(n894 ,n2718 ,n846);
    nand g2601(n2141 ,n2045 ,n2108);
    nand g2602(n2105 ,n1951 ,n2034);
    nand g2603(n2355 ,n2314 ,n2334);
    nand g2604(n60 ,n30[3] ,n59);
    nand g2605(n1800 ,n1663 ,n1662);
    nor g2606(n1150 ,n975 ,n1133);
    nor g2607(n1334 ,n1267 ,n1303);
    nand g2608(n1247 ,n1215 ,n1246);
    dff g2609(.RN(n1), .SN(1'b1), .CK(n0), .D(n403), .Q(n26[1]));
    nor g2610(n2199 ,n2140 ,n2138);
    xnor g2611(n2283 ,n2217 ,n2168);
    nand g2612(n589 ,n23[7] ,n480);
    buf g2613(n9[13], 1'b0);
    nand g2614(n487 ,n6[1] ,n477);
    nand g2615(n2114 ,n2022 ,n2064);
    dff g2616(.RN(n1), .SN(1'b1), .CK(n0), .D(n369), .Q(n28[13]));
    xnor g2617(n1836 ,n1581 ,n1650);
    not g2618(n2050 ,n2049);
    not g2619(n40 ,n30[7]);
    or g2620(n1932 ,n1870 ,n1864);
    dff g2621(.RN(n1), .SN(1'b1), .CK(n0), .D(n645), .Q(n21[0]));
    nand g2622(n2056 ,n1935 ,n1964);
    nor g2623(n1207 ,n1153 ,n1204);
    nand g2624(n75 ,n25[5] ,n73);
    buf g2625(n9[9], 1'b0);
    nor g2626(n1373 ,n1287 ,n1336);
    nand g2627(n330 ,n752 ,n141);
    xnor g2628(n134 ,n19[0] ,n28[0]);
    nand g2629(n2436 ,n2374 ,n2435);
    xnor g2630(n1113 ,n1069 ,n992);
    xnor g2631(n2669 ,n2497 ,n2527);
    nand g2632(n188 ,n29[11] ,n140);
    xnor g2633(n2051 ,n1907 ,n1923);
    nand g2634(n2628 ,n2577 ,n2610);
    nor g2635(n1903 ,n1642 ,n1816);
    nand g2636(n661 ,n554 ,n487);
    xnor g2637(n1852 ,n1628 ,n1704);
    nor g2638(n107 ,n5[3] ,n5[2]);
    xnor g2639(n1971 ,n1824 ,n1639);
    nor g2640(n1386 ,n1310 ,n1366);
    nor g2641(n1383 ,n1293 ,n1357);
    not g2642(n71 ,n70);
    nand g2643(n331 ,n31[4] ,n141);
    nand g2644(n2080 ,n1733 ,n2010);
    nand g2645(n550 ,n19[5] ,n476);
    buf g2646(n11[6], 1'b0);
    nand g2647(n1911 ,n1808 ,n1856);
    nand g2648(n2428 ,n2413 ,n2427);
    nor g2649(n1170 ,n1149 ,n1115);
    dff g2650(.RN(n1), .SN(1'b1), .CK(n0), .D(n640), .Q(n21[5]));
    nand g2651(n2011 ,n1950 ,n1933);
    xnor g2652(n2029 ,n1915 ,n1916);
    xnor g2653(n1547 ,n1528 ,n1519);
    nand g2654(n1663 ,n20[2] ,n22[4]);
    xnor g2655(n2721 ,n2501 ,n2521);
    xnor g2656(n993 ,n940 ,n816);
    dff g2657(.RN(n1), .SN(1'b1), .CK(n0), .D(n695), .Q(n23[5]));
    nand g2658(n1606 ,n21[6] ,n23[5]);
    xnor g2659(n1403 ,n1363 ,n1327);
    nand g2660(n1420 ,n1370 ,n1388);
    nand g2661(n450 ,n181 ,n446);
    xnor g2662(n2281 ,n2216 ,n2193);
    nand g2663(n1690 ,n21[5] ,n23[5]);
    dff g2664(.RN(n1), .SN(1'b1), .CK(n0), .D(n418), .Q(n10[11]));
    buf g2665(n11[9], 1'b0);
    or g2666(n2180 ,n2101 ,n2131);
    nor g2667(n1093 ,n959 ,n1076);
    not g2668(n1456 ,n1455);
    nand g2669(n709 ,n576 ,n527);
    nor g2670(n1762 ,n1628 ,n1704);
    nand g2671(n2591 ,n32[8] ,n2561);
    nand g2672(n551 ,n19[4] ,n476);
    nor g2673(n1198 ,n1163 ,n1177);
    xnor g2674(n1065 ,n984 ,n1015);
    not g2675(n1201 ,n1200);
    xnor g2676(n1504 ,n1470 ,n1428);
    xor g2677(n1839 ,n1627 ,n1604);
    nand g2678(n599 ,n22[5] ,n469);
    not g2679(n1624 ,n1623);
    nor g2680(n973 ,n927 ,n930);
    xor g2681(n2025 ,n1951 ,n1921);
    nand g2682(n907 ,n792 ,n859);
    nand g2683(n338 ,n741 ,n144);
    not g2684(n52 ,n51);
    nand g2685(n1601 ,n21[7] ,n23[1]);
    nand g2686(n2397 ,n2372 ,n2387);
    nand g2687(n1895 ,n1631 ,n1794);
    nor g2688(n1289 ,n1269 ,n1284);
    xnor g2689(n2667 ,n2523 ,n2494);
    or g2690(n1129 ,n1089 ,n1094);
    nand g2691(n190 ,n29[8] ,n87);
    or g2692(n2044 ,n1938 ,n1982);
    not g2693(n821 ,n822);
    nand g2694(n208 ,n28[0] ,n87);
    or g2695(n31[5] ,n2623 ,n2663);
    nor g2696(n1346 ,n1268 ,n1304);
    nand g2697(n2594 ,n2694 ,n2546);
    nand g2698(n1666 ,n21[7] ,n23[2]);
    not g2699(n1857 ,n1856);
    xnor g2700(n2496 ,n2698 ,n2682);
    buf g2701(n17[7], 1'b0);
    or g2702(n2036 ,n1988 ,n1976);
    or g2703(n2096 ,n1975 ,n2046);
    nand g2704(n1898 ,n1638 ,n1780);
    dff g2705(.RN(n1), .SN(1'b1), .CK(n0), .D(n388), .Q(n26[12]));
    nand g2706(n252 ,n3 ,n155);
    nand g2707(n669 ,n593 ,n592);
    nand g2708(n801 ,n767 ,n780);
    nand g2709(n2551 ,n2730 ,n32[3]);
    nand g2710(n2602 ,n32[4] ,n2561);
    nand g2711(n408 ,n198 ,n306);
    xor g2712(n2678 ,n20[6] ,n21[6]);
    nor g2713(n1294 ,n1266 ,n1278);
    nand g2714(n366 ,n209 ,n280);
    buf g2715(n10[19], 1'b0);
    buf g2716(n11[19], n10[3]);
    buf g2717(n10[25], 1'b0);
    xor g2718(n2713 ,n2449 ,n2440);
    nand g2719(n1554 ,n1544 ,n1553);
    nand g2720(n2459 ,n2443 ,n2458);
    not g2721(n1267 ,n24[3]);
    nand g2722(n2155 ,n2069 ,n2103);
    nand g2723(n2329 ,n2271 ,n2306);
    nor g2724(n1262 ,n1217 ,n1261);
    nand g2725(n909 ,n2714 ,n876);
    nor g2726(n1249 ,n1248 ,n1214);
    nand g2727(n385 ,n213 ,n278);
    nand g2728(n681 ,n429 ,n615);
    xnor g2729(n2172 ,n2052 ,n2119);
    xnor g2730(n2295 ,n2183 ,n2277);
    buf g2731(n13[0], 1'b0);
    nor g2732(n2107 ,n1953 ,n2076);
    nor g2733(n1101 ,n1036 ,n1080);
    nand g2734(n1779 ,n1581 ,n1650);
    nor g2735(n1027 ,n966 ,n1009);
    xnor g2736(n2088 ,n2016 ,n2014);
    nor g2737(n1872 ,n1595 ,n1761);
    xnor g2738(n2085 ,n1967 ,n1969);
    nand g2739(n878 ,n2714 ,n847);
    not g2740(n1635 ,n1634);
    nand g2741(n603 ,n20[5] ,n468);
    or g2742(n2394 ,n2362 ,n2389);
    dff g2743(.RN(n1), .SN(1'b1), .CK(n0), .D(n371), .Q(n28[11]));
    nand g2744(n897 ,n2717 ,n847);
    nand g2745(n654 ,n547 ,n486);
    xnor g2746(n1824 ,n1589 ,n1652);
    nor g2747(n2235 ,n2166 ,n2199);
    nand g2748(n1049 ,n987 ,n985);
    nand g2749(n1904 ,n1641 ,n1775);
    nand g2750(n369 ,n244 ,n274);
    dff g2751(.RN(n1), .SN(1'b1), .CK(n0), .D(n661), .Q(n19[1]));
    nand g2752(n2371 ,n2280 ,n2352);
    nand g2753(n978 ,n932 ,n930);
    nand g2754(n415 ,n314 ,n235);
    xnor g2755(n2490 ,n2710 ,n2694);
    nor g2756(n2520 ,n2487 ,n2519);
    nor g2757(n464 ,n344 ,n456);
    xnor g2758(n2343 ,n2295 ,n2229);
    or g2759(n31[12] ,n2625 ,n2639);
    nand g2760(n1920 ,n1746 ,n1875);
    xnor g2761(n2171 ,n1971 ,n2102);
    nand g2762(n2247 ,n2110 ,n2204);
    xnor g2763(n1000 ,n818 ,n939);
    nand g2764(n265 ,n28[7] ,n87);
    xnor g2765(n1979 ,n1840 ,n1602);
    xnor g2766(n1983 ,n1825 ,n1620);
    nand g2767(n1492 ,n1413 ,n1474);
    nand g2768(n2598 ,n2670 ,n2559);
    dff g2769(.RN(n1), .SN(1'b1), .CK(n0), .D(n450), .Q(n18[2]));
    nand g2770(n315 ,n10[13] ,n156);
    nand g2771(n1465 ,n1420 ,n1264);
    nand g2772(n1652 ,n21[4] ,n23[5]);
    nand g2773(n359 ,n14 ,n345);
    nand g2774(n437 ,n9[1] ,n252);
    xnor g2775(n2404 ,n2379 ,n2353);
    not g2776(n2452 ,n2451);
    nand g2777(n827 ,n2712 ,n819);
    nand g2778(n232 ,n25[2] ,n142);
    nand g2779(n1643 ,n20[3] ,n22[1]);
    nand g2780(n2622 ,n2688 ,n2546);
    nand g2781(n526 ,n6[5] ,n479);
    not g2782(n476 ,n477);
    nand g2783(n687 ,n561 ,n516);
    nand g2784(n31[15] ,n2620 ,n2638);
    buf g2785(n9[17], 1'b0);
    not g2786(n2638 ,n2626);
    xnor g2787(n2693 ,n2401 ,n2432);
    nand g2788(n343 ,n29[5] ,n141);
    nand g2789(n2657 ,n2575 ,n2624);
    nor g2790(n1236 ,n1220 ,n1231);
    nand g2791(n2663 ,n2593 ,n2651);
    nor g2792(n2564 ,n2560 ,n2537);
    nand g2793(n1619 ,n20[4] ,n22[1]);
    nand g2794(n1797 ,n1725 ,n1649);
    nand g2795(n1928 ,n1754 ,n1892);
    nor g2796(n1460 ,n1404 ,n1443);
    xnor g2797(n1007 ,n952 ,n817);
    nand g2798(n493 ,n6[1] ,n479);
    nand g2799(n1047 ,n986 ,n991);
    xnor g2800(n745 ,n25[4] ,n72);
    nand g2801(n154 ,n120 ,n112);
    nand g2802(n206 ,n28[3] ,n87);
    not g2803(n1297 ,n1298);
    xnor g2804(n775 ,n21[7] ,n20[7]);
    nand g2805(n1444 ,n1427 ,n1263);
    not g2806(n960 ,n959);
    nand g2807(n2288 ,n2277 ,n2256);
    nand g2808(n407 ,n231 ,n305);
    xnor g2809(n2718 ,n2447 ,n2465);
    or g2810(n2310 ,n2231 ,n2286);
    nand g2811(n621 ,n23[2] ,n480);
    nand g2812(n448 ,n142 ,n360);
    nand g2813(n537 ,n21[2] ,n463);
    nand g2814(n294 ,n29[8] ,n141);
    xnor g2815(n1503 ,n1474 ,n1413);
    nand g2816(n565 ,n23[7] ,n474);
    nand g2817(n212 ,n25[7] ,n142);
    nand g2818(n306 ,n744 ,n143);
    nand g2819(n362 ,n188 ,n268);
    xnor g2820(n2341 ,n2305 ,n2322);
    nand g2821(n1702 ,n21[1] ,n23[4]);
    buf g2822(n10[27], 1'b0);
    nand g2823(n319 ,n10[9] ,n156);
    nand g2824(n1487 ,n1447 ,n1471);
    nand g2825(n980 ,n817 ,n938);
    or g2826(n31[11] ,n2641 ,n2633);
    or g2827(n1760 ,n1655 ,n1604);
    buf g2828(n17[1], 1'b0);
    nand g2829(n1640 ,n21[0] ,n23[7]);
    nand g2830(n1664 ,n20[5] ,n22[3]);
    nand g2831(n788 ,n2716 ,n783);
    nor g2832(n470 ,n344 ,n454);
    nand g2833(n2457 ,n2437 ,n2456);
    xnor g2834(n1817 ,n1580 ,n1680);
    nand g2835(n955 ,n872 ,n894);
    or g2836(n41 ,n30[4] ,n30[3]);
    dff g2837(.RN(n1), .SN(1'b1), .CK(n0), .D(n414), .Q(n10[15]));
    nor g2838(n2572 ,n2560 ,n2544);
    xnor g2839(n1124 ,n1066 ,n993);
    nand g2840(n610 ,n19[4] ,n481);
    nand g2841(n356 ,n201 ,n172);
    buf g2842(n11[23], n10[7]);
    nor g2843(n81 ,n157 ,n394);
    buf g2844(n12[11], n10[3]);
    or g2845(n1510 ,n1330 ,n1500);
    nand g2846(n2095 ,n1949 ,n2056);
    nand g2847(n240 ,n31[7] ,n155);
    not g2848(n163 ,n162);
    dff g2849(.RN(n1), .SN(1'b1), .CK(n0), .D(n409), .Q(n25[4]));
    or g2850(n1532 ,n1515 ,n1517);
    nand g2851(n523 ,n6[2] ,n475);
    nand g2852(n340 ,n754 ,n141);
    xnor g2853(n2091 ,n1977 ,n1990);
    or g2854(n2156 ,n1979 ,n1565);
    nand g2855(n1577 ,n21[4] ,n23[0]);
    xnor g2856(n1096 ,n1024 ,n1018);
    nand g2857(n1891 ,n1706 ,n1785);
    xnor g2858(n2252 ,n2078 ,n2191);
    nand g2859(n1798 ,n1692 ,n1587);
    nand g2860(n2256 ,n2183 ,n2229);
    nand g2861(n2655 ,n2576 ,n2627);
    xnor g2862(n2262 ,n2175 ,n2131);
    nand g2863(n2338 ,n2293 ,n2300);
    xnor g2864(n2183 ,n2090 ,n1992);
    xnor g2865(n130 ,n19[4] ,n28[4]);
    nand g2866(n279 ,n31[7] ,n141);
    xnor g2867(n2451 ,n23[5] ,n22[5]);
    nor g2868(n2196 ,n2048 ,n2134);
    nand g2869(n210 ,n28[1] ,n140);
    nor g2870(n1404 ,n1309 ,n1392);
    nor g2871(n1234 ,n1195 ,n1232);
    xnor g2872(n1990 ,n1830 ,n1637);
    not g2873(n1816 ,n1803);
    nand g2874(n2552 ,n2729 ,n32[4]);
    xnor g2875(n1066 ,n1000 ,n1007);
    xnor g2876(n2401 ,n2389 ,n2362);
    nand g2877(n2478 ,n2709 ,n2693);
    nand g2878(n2039 ,n1926 ,n2012);
    or g2879(n740 ,n30[6] ,n46);
    nand g2880(n979 ,n818 ,n939);
    nand g2881(n2018 ,n1728 ,n1934);
    not g2882(n1061 ,n1044);
    nor g2883(n2523 ,n2474 ,n2522);
    or g2884(n2012 ,n1919 ,n1939);
    nand g2885(n296 ,n29[6] ,n141);
    nand g2886(n506 ,n6[7] ,n477);
    buf g2887(n17[5], 1'b0);
    nand g2888(n885 ,n2718 ,n847);
    nor g2889(n2075 ,n1941 ,n1983);
    not g2890(n76 ,n75);
    xnor g2891(n2702 ,n1205 ,n1232);
    nand g2892(n2154 ,n2102 ,n2097);
    nand g2893(n46 ,n40 ,n45);
    not g2894(n1397 ,n1396);
    nand g2895(n2363 ,n2328 ,n2348);
    dff g2896(.RN(n1), .SN(1'b1), .CK(n0), .D(n734), .Q(n9[6]));
    nand g2897(n2407 ,n2398 ,n2381);
    xnor g2898(n1023 ,n920 ,n957);
    nand g2899(n1720 ,n21[1] ,n23[3]);
    xnor g2900(n1995 ,n1858 ,n1762);
    nand g2901(n1661 ,n20[1] ,n22[4]);
    nand g2902(n2592 ,n32[2] ,n2561);
    nand g2903(n2557 ,n2723 ,n32[10]);
    nand g2904(n441 ,n263 ,n297);
    nand g2905(n484 ,n6[0] ,n464);
    nand g2906(n1284 ,n2677 ,n23[5]);
    nand g2907(n738 ,n728 ,n719);
    nand g2908(n370 ,n190 ,n270);
    xnor g2909(n2376 ,n2302 ,n2351);
    nand g2910(n2374 ,n2302 ,n2351);
    dff g2911(.RN(n1), .SN(1'b1), .CK(n0), .D(n687), .Q(n24[3]));
    or g2912(n1277 ,n2674 ,n23[2]);
    nor g2913(n124 ,n88 ,n5[2]);
    xnor g2914(n1138 ,n1091 ,n1025);
    or g2915(n31[10] ,n2629 ,n2657);
    nand g2916(n631 ,n24[0] ,n482);
    nand g2917(n236 ,n31[12] ,n155);
    not g2918(n141 ,n87);
    nor g2919(n85 ,n5[1] ,n5[0]);
    nor g2920(n1873 ,n1667 ,n1766);
    buf g2921(n11[16], n10[0]);
    nand g2922(n918 ,n2719 ,n847);
    nand g2923(n902 ,n2720 ,n847);
    nand g2924(n2408 ,n2388 ,n2395);
    nand g2925(n632 ,n23[6] ,n480);
    nand g2926(n1365 ,n24[0] ,n1302);
    not g2927(n1062 ,n1049);
    or g2928(n87 ,n18[2] ,n121);
    nand g2929(n840 ,n2713 ,n820);
    nor g2930(n1152 ,n1098 ,n1123);
    nand g2931(n388 ,n217 ,n291);
    buf g2932(n11[12], 1'b0);
    not g2933(n155 ,n156);
    xnor g2934(n2668 ,n2488 ,n2525);
    nor g2935(n1179 ,n1132 ,n1155);
    nand g2936(n843 ,n2713 ,n821);
    nand g2937(n1524 ,n1496 ,n1509);
    not g2938(n635 ,n604);
    or g2939(n1274 ,n2676 ,n23[4]);
    nor g2940(n84 ,n158 ,n159);
    nand g2941(n562 ,n24[2] ,n461);
    nand g2942(n364 ,n189 ,n277);
    nand g2943(n521 ,n6[4] ,n475);
    nand g2944(n427 ,n326 ,n245);
    dff g2945(.RN(n1), .SN(1'b1), .CK(n0), .D(n686), .Q(n24[4]));
    nand g2946(n435 ,n193 ,n334);
    nor g2947(n1380 ,n1288 ,n1341);
    nand g2948(n268 ,n28[11] ,n141);
    nor g2949(n1261 ,n1216 ,n1260);
    dff g2950(.RN(n1), .SN(1'b1), .CK(n0), .D(n182), .Q(n17[2]));
    nand g2951(n712 ,n581 ,n530);
    nand g2952(n2280 ,n2225 ,n2266);
    xnor g2953(n2031 ,n1922 ,n1764);
    nand g2954(n1572 ,n21[0] ,n23[3]);
    nand g2955(n1111 ,n1050 ,n1087);
    xnor g2956(n2284 ,n2215 ,n2167);
    nand g2957(n1900 ,n1563 ,n1773);
    xnor g2958(n2191 ,n2084 ,n2103);
    nand g2959(n1637 ,n21[0] ,n23[6]);
    nor g2960(n184 ,n741 ,n145);
    buf g2961(n12[3], 1'b0);
    nand g2962(n674 ,n413 ,n603);
    dff g2963(.RN(n1), .SN(1'b1), .CK(n0), .D(n427), .Q(n10[3]));
    nand g2964(n508 ,n6[5] ,n477);
    nor g2965(n1360 ,n1269 ,n1305);
    nand g2966(n354 ,n195 ,n174);
    xnor g2967(n1467 ,n1441 ,n1389);
    nor g2968(n2203 ,n2139 ,n2137);
    nand g2969(n732 ,n726 ,n717);
    or g2970(n165 ,n160 ,n162);
    nor g2971(n1355 ,n1266 ,n1301);
    nand g2972(n584 ,n22[0] ,n469);
    xor g2973(n2027 ,n1925 ,n1944);
    nand g2974(n2627 ,n2548 ,n2562);
    nand g2975(n914 ,n2718 ,n876);
    not g2976(n634 ,n598);
    nand g2977(n1581 ,n20[4] ,n22[5]);
    xnor g2978(n2705 ,n1221 ,n1249);
    xnor g2979(n393 ,n142 ,n25[0]);
    nand g2980(n308 ,n745 ,n143);
    nand g2981(n1173 ,n1127 ,n1151);
    nand g2982(n2319 ,n2242 ,n2279);
    xnor g2983(n1008 ,n817 ,n938);
    not g2984(n1638 ,n1637);
    nand g2985(n574 ,n22[6] ,n478);
    nand g2986(n2315 ,n2211 ,n2281);
    nand g2987(n2223 ,n2135 ,n2187);
    xnor g2988(n1125 ,n1067 ,n999);
    xnor g2989(n754 ,n30[2] ,n56);
    xnor g2990(n1844 ,n1675 ,n1668);
    nand g2991(n690 ,n563 ,n489);
    nand g2992(n1553 ,n1532 ,n1552);
    xnor g2993(n965 ,n806 ,n900);
    nand g2994(n363 ,n251 ,n271);
    buf g2995(n11[17], n10[1]);
    nor g2996(n2517 ,n2469 ,n2516);
    not g2997(n1918 ,n1917);
    nand g2998(n350 ,n160 ,n183);
    nand g2999(n409 ,n215 ,n308);
    nand g3000(n700 ,n570 ,n523);
    xnor g3001(n963 ,n806 ,n899);
    buf g3002(n13[22], 1'b0);
    nand g3003(n1029 ,n1015 ,n984);
    nand g3004(n1511 ,n1330 ,n1500);
    nand g3005(n676 ,n608 ,n607);
    nor g3006(n1238 ,n1200 ,n1224);
    or g3007(n2234 ,n2078 ,n2191);
    nand g3008(n1602 ,n21[1] ,n23[1]);
    nand g3009(n321 ,n10[7] ,n156);
    xnor g3010(n2723 ,n2485 ,n2517);
    nand g3011(n873 ,n2720 ,n824);
    nand g3012(n2641 ,n2589 ,n2585);
    nor g3013(n1317 ,n1269 ,n1278);
endmodule
