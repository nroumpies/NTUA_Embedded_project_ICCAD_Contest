module top (n0, n1, n2, n3, n4, n5, n6, n8, n9, n7, n10, n11, n12, n13, n14, n15);
    input n0, n1;
    input [7:0] n2, n3, n4, n5, n6, n7;
    input [2:0] n8;
    input [3:0] n9;
    output [15:0] n10, n11, n12, n13, n14;
    output [7:0] n15;
    wire n0, n1;
    wire [7:0] n2, n3, n4, n5, n6, n7;
    wire [2:0] n8;
    wire [3:0] n9;
    wire [15:0] n10, n11, n12, n13, n14;
    wire [7:0] n15;
    wire [15:0] n16;
    wire [15:0] n17;
    wire [3:0] n18;
    wire [7:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [15:0] n22;
    wire [15:0] n23;
    wire [7:0] n24;
    wire [2:0] n25;
    wire [15:0] n26;
    wire [15:0] n27;
    wire [15:0] n28;
    wire [15:0] n29;
    wire [15:0] n30;
    wire [15:0] n31;
    wire [7:0] n32;
    wire [15:0] n33;
    wire [15:0] n34;
    wire [15:0] n35;
    wire [7:0] n36;
    wire [7:0] n37;
    wire [15:0] n38;
    wire [15:0] n39;
    wire [15:0] n40;
    wire [15:0] n41;
    wire n42, n43, n44, n45, n46, n47, n48, n49;
    wire n50, n51, n52, n53, n54, n55, n56, n57;
    wire n58, n59, n60, n61, n62, n63, n64, n65;
    wire n66, n67, n68, n69, n70, n71, n72, n73;
    wire n74, n75, n76, n77, n78, n79, n80, n81;
    wire n82, n83, n84, n85, n86, n87, n88, n89;
    wire n90, n91, n92, n93, n94, n95, n96, n97;
    wire n98, n99, n100, n101, n102, n103, n104, n105;
    wire n106, n107, n108, n109, n110, n111, n112, n113;
    wire n114, n115, n116, n117, n118, n119, n120, n121;
    wire n122, n123, n124, n125, n126, n127, n128, n129;
    wire n130, n131, n132, n133, n134, n135, n136, n137;
    wire n138, n139, n140, n141, n142, n143, n144, n145;
    wire n146, n147, n148, n149, n150, n151, n152, n153;
    wire n154, n155, n156, n157, n158, n159, n160, n161;
    wire n162, n163, n164, n165, n166, n167, n168, n169;
    wire n170, n171, n172, n173, n174, n175, n176, n177;
    wire n178, n179, n180, n181, n182, n183, n184, n185;
    wire n186, n187, n188, n189, n190, n191, n192, n193;
    wire n194, n195, n196, n197, n198, n199, n200, n201;
    wire n202, n203, n204, n205, n206, n207, n208, n209;
    wire n210, n211, n212, n213, n214, n215, n216, n217;
    wire n218, n219, n220, n221, n222, n223, n224, n225;
    wire n226, n227, n228, n229, n230, n231, n232, n233;
    wire n234, n235, n236, n237, n238, n239, n240, n241;
    wire n242, n243, n244, n245, n246, n247, n248, n249;
    wire n250, n251, n252, n253, n254, n255, n256, n257;
    wire n258, n259, n260, n261, n262, n263, n264, n265;
    wire n266, n267, n268, n269, n270, n271, n272, n273;
    wire n274, n275, n276, n277, n278, n279, n280, n281;
    wire n282, n283, n284, n285, n286, n287, n288, n289;
    wire n290, n291, n292, n293, n294, n295, n296, n297;
    wire n298, n299, n300, n301, n302, n303, n304, n305;
    wire n306, n307, n308, n309, n310, n311, n312, n313;
    wire n314, n315, n316, n317, n318, n319, n320, n321;
    wire n322, n323, n324, n325, n326, n327, n328, n329;
    wire n330, n331, n332, n333, n334, n335, n336, n337;
    wire n338, n339, n340, n341, n342, n343, n344, n345;
    wire n346, n347, n348, n349, n350, n351, n352, n353;
    wire n354, n355, n356, n357, n358, n359, n360, n361;
    wire n362, n363, n364, n365, n366, n367, n368, n369;
    wire n370, n371, n372, n373, n374, n375, n376, n377;
    wire n378, n379, n380, n381, n382, n383, n384, n385;
    wire n386, n387, n388, n389, n390, n391, n392, n393;
    wire n394, n395, n396, n397, n398, n399, n400, n401;
    wire n402, n403, n404, n405, n406, n407, n408, n409;
    wire n410, n411, n412, n413, n414, n415, n416, n417;
    wire n418, n419, n420, n421, n422, n423, n424, n425;
    wire n426, n427, n428, n429, n430, n431, n432, n433;
    wire n434, n435, n436, n437, n438, n439, n440, n441;
    wire n442, n443, n444, n445, n446, n447, n448, n449;
    wire n450, n451, n452, n453, n454, n455, n456, n457;
    wire n458, n459, n460, n461, n462, n463, n464, n465;
    wire n466, n467, n468, n469, n470, n471, n472, n473;
    wire n474, n475, n476, n477, n478, n479, n480, n481;
    wire n482, n483, n484, n485, n486, n487, n488, n489;
    wire n490, n491, n492, n493, n494, n495, n496, n497;
    wire n498, n499, n500, n501, n502, n503, n504, n505;
    wire n506, n507, n508, n509, n510, n511, n512, n513;
    wire n514, n515, n516, n517, n518, n519, n520, n521;
    wire n522, n523, n524, n525, n526, n527, n528, n529;
    wire n530, n531, n532, n533, n534, n535, n536, n537;
    wire n538, n539, n540, n541, n542, n543, n544, n545;
    wire n546, n547, n548, n549, n550, n551, n552, n553;
    wire n554, n555, n556, n557, n558, n559, n560, n561;
    wire n562, n563, n564, n565, n566, n567, n568, n569;
    wire n570, n571, n572, n573, n574, n575, n576, n577;
    wire n578, n579, n580, n581, n582, n583, n584, n585;
    wire n586, n587, n588, n589, n590, n591, n592, n593;
    wire n594, n595, n596, n597, n598, n599, n600, n601;
    wire n602, n603, n604, n605, n606, n607, n608, n609;
    wire n610, n611, n612, n613, n614, n615, n616, n617;
    wire n618, n619, n620, n621, n622, n623, n624, n625;
    wire n626, n627, n628, n629, n630, n631, n632, n633;
    wire n634, n635, n636, n637, n638, n639, n640, n641;
    wire n642, n643, n644, n645, n646, n647, n648, n649;
    wire n650, n651, n652, n653, n654, n655, n656, n657;
    wire n658, n659, n660, n661, n662, n663, n664, n665;
    wire n666, n667, n668, n669, n670, n671, n672, n673;
    wire n674, n675, n676, n677, n678, n679, n680, n681;
    wire n682, n683, n684, n685, n686, n687, n688, n689;
    wire n690, n691, n692, n693, n694, n695, n696, n697;
    wire n698, n699, n700, n701, n702, n703, n704, n705;
    wire n706, n707, n708, n709, n710, n711, n712, n713;
    wire n714, n715, n716, n717, n718, n719, n720, n721;
    wire n722, n723, n724, n725, n726, n727, n728, n729;
    wire n730, n731, n732, n733, n734, n735, n736, n737;
    wire n738, n739, n740, n741, n742, n743, n744, n745;
    wire n746, n747, n748, n749, n750, n751, n752, n753;
    wire n754, n755, n756, n757, n758, n759, n760, n761;
    wire n762, n763, n764, n765, n766, n767, n768, n769;
    wire n770, n771, n772, n773, n774, n775, n776, n777;
    wire n778, n779, n780, n781, n782, n783, n784, n785;
    wire n786, n787, n788, n789, n790, n791, n792, n793;
    wire n794, n795, n796, n797, n798, n799, n800, n801;
    wire n802, n803, n804, n805, n806, n807, n808, n809;
    wire n810, n811, n812, n813, n814, n815, n816, n817;
    wire n818, n819, n820, n821, n822, n823, n824, n825;
    wire n826, n827, n828, n829, n830, n831, n832, n833;
    wire n834, n835, n836, n837, n838, n839, n840, n841;
    wire n842, n843, n844, n845, n846, n847, n848, n849;
    wire n850, n851, n852, n853, n854, n855, n856, n857;
    wire n858, n859, n860, n861, n862, n863, n864, n865;
    wire n866, n867, n868, n869, n870, n871, n872, n873;
    wire n874, n875, n876, n877, n878, n879, n880, n881;
    wire n882, n883, n884, n885, n886, n887, n888, n889;
    wire n890, n891, n892, n893, n894, n895, n896, n897;
    wire n898, n899, n900, n901, n902, n903, n904, n905;
    wire n906, n907, n908, n909, n910, n911, n912, n913;
    wire n914, n915, n916, n917, n918, n919, n920, n921;
    wire n922, n923, n924, n925, n926, n927, n928, n929;
    wire n930, n931, n932, n933, n934, n935, n936, n937;
    wire n938, n939, n940, n941, n942, n943, n944, n945;
    wire n946, n947, n948, n949, n950, n951, n952, n953;
    wire n954, n955, n956, n957, n958, n959, n960, n961;
    wire n962, n963, n964, n965, n966, n967, n968, n969;
    wire n970, n971, n972, n973, n974, n975, n976, n977;
    wire n978, n979, n980, n981, n982, n983, n984, n985;
    wire n986, n987, n988, n989, n990, n991, n992, n993;
    wire n994, n995, n996, n997, n998, n999, n1000, n1001;
    wire n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009;
    wire n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017;
    wire n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
    wire n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
    wire n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041;
    wire n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049;
    wire n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057;
    wire n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065;
    wire n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073;
    wire n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081;
    wire n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089;
    wire n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097;
    wire n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105;
    wire n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113;
    wire n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121;
    wire n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129;
    wire n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137;
    wire n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145;
    wire n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153;
    wire n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161;
    wire n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169;
    wire n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177;
    wire n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185;
    wire n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193;
    wire n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201;
    wire n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209;
    wire n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217;
    wire n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225;
    wire n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233;
    wire n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241;
    wire n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249;
    wire n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257;
    wire n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265;
    wire n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273;
    wire n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281;
    wire n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289;
    wire n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297;
    wire n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305;
    wire n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313;
    wire n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321;
    wire n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329;
    wire n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;
    wire n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345;
    wire n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353;
    wire n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;
    wire n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369;
    wire n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377;
    wire n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385;
    wire n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393;
    wire n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401;
    wire n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409;
    wire n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417;
    wire n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425;
    wire n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433;
    wire n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441;
    wire n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449;
    wire n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457;
    wire n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465;
    wire n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473;
    wire n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481;
    wire n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489;
    wire n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497;
    wire n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505;
    wire n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513;
    wire n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521;
    wire n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529;
    wire n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537;
    wire n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545;
    wire n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553;
    wire n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561;
    wire n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569;
    wire n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577;
    wire n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585;
    wire n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593;
    wire n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601;
    wire n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609;
    wire n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617;
    wire n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625;
    wire n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633;
    wire n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641;
    wire n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649;
    wire n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657;
    wire n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665;
    wire n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673;
    wire n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681;
    wire n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689;
    wire n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697;
    wire n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705;
    wire n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713;
    wire n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721;
    wire n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729;
    wire n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737;
    wire n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745;
    wire n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753;
    wire n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761;
    wire n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769;
    wire n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777;
    wire n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785;
    wire n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793;
    wire n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801;
    wire n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809;
    wire n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817;
    wire n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825;
    wire n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833;
    wire n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;
    wire n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849;
    wire n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857;
    wire n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865;
    wire n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873;
    wire n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881;
    wire n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889;
    wire n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897;
    wire n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905;
    wire n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913;
    wire n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921;
    wire n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929;
    wire n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937;
    wire n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945;
    wire n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953;
    wire n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961;
    wire n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969;
    wire n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977;
    wire n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985;
    wire n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993;
    wire n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001;
    wire n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009;
    wire n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017;
    wire n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025;
    wire n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033;
    wire n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041;
    wire n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049;
    wire n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057;
    wire n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065;
    wire n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073;
    wire n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081;
    wire n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089;
    wire n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097;
    wire n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105;
    wire n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113;
    wire n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121;
    wire n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129;
    wire n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137;
    wire n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145;
    wire n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153;
    wire n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161;
    wire n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169;
    wire n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177;
    wire n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185;
    wire n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193;
    wire n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201;
    wire n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209;
    wire n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217;
    wire n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225;
    wire n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233;
    wire n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241;
    wire n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249;
    wire n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257;
    wire n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265;
    wire n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273;
    wire n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281;
    wire n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289;
    wire n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297;
    wire n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305;
    wire n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313;
    wire n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321;
    wire n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329;
    wire n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337;
    wire n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345;
    wire n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353;
    wire n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361;
    wire n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369;
    wire n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377;
    wire n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385;
    wire n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393;
    wire n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401;
    wire n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409;
    wire n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417;
    wire n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425;
    wire n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433;
    wire n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441;
    wire n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449;
    wire n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457;
    wire n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465;
    wire n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473;
    wire n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481;
    wire n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489;
    wire n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497;
    wire n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505;
    wire n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513;
    wire n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521;
    wire n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529;
    wire n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537;
    wire n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545;
    wire n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553;
    wire n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561;
    wire n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569;
    wire n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577;
    wire n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585;
    wire n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593;
    wire n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601;
    wire n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609;
    wire n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617;
    wire n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625;
    wire n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633;
    wire n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641;
    wire n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649;
    wire n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657;
    wire n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665;
    wire n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673;
    wire n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681;
    wire n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689;
    wire n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697;
    wire n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705;
    wire n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713;
    wire n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721;
    wire n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729;
    wire n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737;
    wire n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745;
    wire n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753;
    wire n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761;
    wire n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769;
    wire n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777;
    wire n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785;
    wire n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793;
    wire n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801;
    wire n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809;
    wire n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817;
    wire n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825;
    wire n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833;
    wire n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841;
    wire n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849;
    wire n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857;
    wire n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865;
    wire n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873;
    wire n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881;
    wire n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889;
    wire n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897;
    wire n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905;
    wire n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913;
    wire n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921;
    wire n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929;
    wire n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937;
    wire n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945;
    wire n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953;
    wire n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961;
    wire n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969;
    wire n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977;
    wire n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985;
    wire n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993;
    wire n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001;
    wire n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009;
    wire n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017;
    wire n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025;
    wire n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033;
    wire n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041;
    wire n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049;
    wire n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057;
    wire n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065;
    wire n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073;
    wire n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081;
    wire n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089;
    wire n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097;
    wire n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105;
    wire n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113;
    wire n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121;
    wire n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129;
    wire n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137;
    wire n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145;
    wire n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153;
    wire n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161;
    wire n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169;
    wire n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177;
    wire n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185;
    wire n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193;
    wire n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201;
    wire n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209;
    wire n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217;
    wire n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225;
    wire n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233;
    wire n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241;
    wire n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249;
    wire n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257;
    wire n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265;
    wire n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273;
    wire n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281;
    wire n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289;
    wire n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297;
    wire n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305;
    wire n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313;
    wire n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321;
    wire n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329;
    wire n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337;
    wire n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345;
    wire n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353;
    wire n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361;
    wire n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369;
    wire n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377;
    wire n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385;
    wire n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393;
    wire n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401;
    wire n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409;
    wire n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417;
    wire n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425;
    wire n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433;
    wire n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441;
    wire n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449;
    wire n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457;
    wire n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465;
    wire n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473;
    wire n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481;
    wire n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489;
    wire n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497;
    wire n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505;
    wire n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513;
    wire n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521;
    wire n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529;
    wire n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537;
    wire n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545;
    wire n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553;
    wire n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561;
    wire n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569;
    wire n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577;
    wire n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585;
    wire n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593;
    wire n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601;
    wire n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609;
    wire n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617;
    wire n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625;
    wire n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633;
    wire n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641;
    wire n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649;
    wire n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657;
    wire n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665;
    wire n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673;
    wire n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681;
    wire n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689;
    wire n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697;
    wire n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705;
    wire n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713;
    wire n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721;
    wire n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729;
    wire n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737;
    wire n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745;
    wire n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753;
    wire n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761;
    wire n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769;
    wire n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777;
    wire n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785;
    wire n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793;
    wire n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801;
    wire n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809;
    wire n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817;
    wire n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825;
    wire n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833;
    wire n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841;
    wire n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849;
    wire n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857;
    wire n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865;
    wire n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873;
    wire n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881;
    wire n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889;
    wire n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897;
    wire n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905;
    wire n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913;
    wire n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921;
    wire n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929;
    wire n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937;
    wire n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945;
    wire n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953;
    wire n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961;
    wire n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969;
    wire n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977;
    wire n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985;
    wire n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993;
    wire n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001;
    wire n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009;
    wire n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017;
    wire n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025;
    wire n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033;
    wire n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041;
    wire n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049;
    wire n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057;
    wire n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065;
    wire n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073;
    wire n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081;
    wire n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089;
    wire n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097;
    wire n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105;
    wire n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113;
    wire n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121;
    wire n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129;
    wire n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137;
    wire n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145;
    wire n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153;
    wire n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161;
    wire n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169;
    wire n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177;
    wire n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185;
    wire n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193;
    wire n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201;
    wire n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209;
    wire n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217;
    wire n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225;
    wire n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233;
    wire n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241;
    wire n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249;
    wire n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257;
    wire n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265;
    wire n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273;
    wire n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281;
    wire n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289;
    wire n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297;
    wire n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305;
    wire n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313;
    wire n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321;
    wire n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329;
    wire n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337;
    wire n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345;
    wire n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353;
    wire n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361;
    wire n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369;
    wire n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377;
    wire n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385;
    wire n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393;
    wire n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401;
    wire n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409;
    wire n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417;
    wire n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425;
    wire n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433;
    wire n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441;
    wire n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449;
    wire n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457;
    wire n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465;
    wire n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473;
    wire n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481;
    wire n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489;
    wire n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497;
    wire n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505;
    wire n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513;
    wire n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521;
    wire n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529;
    wire n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537;
    wire n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545;
    wire n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553;
    wire n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561;
    wire n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569;
    wire n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577;
    wire n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585;
    wire n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593;
    wire n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601;
    wire n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609;
    wire n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617;
    wire n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625;
    wire n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633;
    wire n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641;
    wire n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649;
    wire n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657;
    wire n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665;
    wire n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673;
    wire n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681;
    wire n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689;
    wire n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697;
    wire n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705;
    wire n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713;
    wire n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721;
    wire n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729;
    wire n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737;
    wire n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745;
    wire n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753;
    wire n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761;
    wire n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769;
    wire n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777;
    wire n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785;
    wire n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793;
    wire n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801;
    wire n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809;
    wire n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817;
    wire n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825;
    wire n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833;
    wire n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841;
    wire n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849;
    wire n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857;
    wire n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865;
    wire n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873;
    wire n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881;
    wire n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889;
    wire n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897;
    wire n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905;
    wire n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913;
    wire n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921;
    wire n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929;
    wire n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937;
    wire n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945;
    wire n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953;
    wire n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961;
    wire n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969;
    wire n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977;
    wire n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985;
    wire n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993;
    wire n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001;
    wire n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009;
    wire n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017;
    wire n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025;
    wire n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033;
    wire n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041;
    wire n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049;
    wire n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057;
    wire n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065;
    wire n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073;
    wire n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081;
    wire n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089;
    wire n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097;
    wire n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105;
    wire n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113;
    wire n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121;
    wire n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129;
    wire n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137;
    wire n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145;
    wire n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153;
    wire n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161;
    wire n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169;
    wire n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177;
    wire n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185;
    wire n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193;
    wire n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201;
    wire n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209;
    wire n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217;
    wire n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225;
    wire n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233;
    wire n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241;
    wire n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249;
    wire n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257;
    wire n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265;
    wire n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273;
    wire n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281;
    wire n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289;
    wire n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297;
    wire n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305;
    wire n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313;
    wire n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321;
    wire n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329;
    wire n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337;
    wire n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345;
    wire n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353;
    wire n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361;
    wire n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369;
    wire n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377;
    wire n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385;
    wire n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393;
    wire n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401;
    wire n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409;
    wire n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417;
    wire n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425;
    wire n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433;
    wire n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441;
    wire n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449;
    wire n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457;
    wire n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465;
    wire n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473;
    wire n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481;
    wire n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489;
    wire n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497;
    wire n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505;
    wire n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513;
    wire n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521;
    wire n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529;
    wire n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537;
    wire n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545;
    wire n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553;
    wire n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561;
    wire n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569;
    wire n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577;
    wire n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585;
    wire n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593;
    wire n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601;
    wire n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609;
    wire n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617;
    wire n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625;
    wire n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633;
    wire n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641;
    wire n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649;
    wire n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657;
    wire n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665;
    wire n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673;
    wire n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681;
    wire n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689;
    wire n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697;
    wire n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705;
    wire n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713;
    wire n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721;
    wire n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729;
    wire n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737;
    wire n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745;
    wire n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753;
    wire n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761;
    wire n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769;
    wire n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777;
    wire n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785;
    wire n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793;
    wire n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801;
    wire n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809;
    wire n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817;
    wire n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825;
    wire n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833;
    wire n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841;
    wire n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849;
    wire n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857;
    wire n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865;
    wire n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873;
    wire n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881;
    wire n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889;
    wire n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897;
    wire n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905;
    wire n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913;
    wire n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921;
    wire n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929;
    wire n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937;
    wire n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945;
    wire n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953;
    wire n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961;
    wire n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969;
    wire n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977;
    wire n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985;
    wire n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993;
    wire n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001;
    wire n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009;
    wire n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017;
    wire n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025;
    wire n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033;
    wire n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041;
    wire n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049;
    wire n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057;
    wire n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065;
    wire n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073;
    wire n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081;
    wire n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089;
    wire n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097;
    wire n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105;
    wire n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113;
    wire n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121;
    wire n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129;
    wire n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137;
    wire n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145;
    wire n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153;
    wire n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161;
    wire n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169;
    wire n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177;
    wire n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185;
    wire n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193;
    wire n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201;
    wire n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209;
    wire n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217;
    wire n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225;
    wire n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233;
    wire n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241;
    wire n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249;
    wire n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257;
    wire n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265;
    wire n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273;
    wire n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281;
    wire n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289;
    wire n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297;
    wire n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305;
    wire n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313;
    wire n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321;
    wire n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329;
    wire n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337;
    wire n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345;
    wire n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353;
    wire n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361;
    wire n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369;
    wire n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377;
    wire n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385;
    wire n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393;
    wire n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401;
    wire n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409;
    wire n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417;
    wire n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425;
    wire n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433;
    wire n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441;
    wire n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449;
    wire n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457;
    wire n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465;
    wire n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473;
    wire n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481;
    wire n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489;
    wire n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497;
    wire n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505;
    wire n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513;
    wire n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521;
    wire n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529;
    wire n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537;
    wire n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545;
    wire n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553;
    wire n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561;
    wire n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569;
    wire n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577;
    wire n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585;
    wire n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593;
    wire n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601;
    wire n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609;
    wire n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617;
    wire n6618;
    nand g0(n398 ,n264 ,n360);
    nor g1(n2967 ,n2837 ,n2932);
    nand g2(n3934 ,n3697 ,n3878);
    nand g3(n1144 ,n27[11] ,n718);
    nand g4(n3714 ,n3546 ,n3502);
    nand g5(n6214 ,n6213 ,n6205);
    nand g6(n4291 ,n4262 ,n4277);
    nor g7(n751 ,n594 ,n711);
    nand g8(n3377 ,n3343 ,n3376);
    nor g9(n3733 ,n3569 ,n3571);
    nand g10(n4871 ,n4428 ,n4438);
    xnor g11(n4310 ,n4266 ,n4276);
    nand g12(n5478 ,n5143 ,n5357);
    nand g13(n1708 ,n1588 ,n1675);
    nand g14(n846 ,n16[4] ,n714);
    nand g15(n2960 ,n2940 ,n2939);
    nand g16(n1376 ,n821 ,n1124);
    nand g17(n3567 ,n3482 ,n19[6]);
    nand g18(n6406 ,n6275 ,n6314);
    nand g19(n5465 ,n5191 ,n5350);
    nand g20(n1199 ,n613 ,n794);
    nor g21(n877 ,n608 ,n555);
    not g22(n4396 ,n4367);
    nor g23(n2010 ,n1974 ,n1991);
    nand g24(n3515 ,n3460 ,n3480);
    nand g25(n35[6] ,n6448 ,n6479);
    nand g26(n4999 ,n4658 ,n4818);
    nor g27(n6451 ,n6399 ,n6397);
    or g28(n6171 ,n6122 ,n6146);
    xor g29(n4946 ,n4510 ,n4459);
    nand g30(n3569 ,n3470 ,n3476);
    nand g31(n1009 ,n12[11] ,n555);
    nand g32(n4453 ,n21[5] ,n4367);
    nand g33(n5587 ,n5349 ,n5484);
    xnor g34(n4056 ,n3945 ,n3897);
    nand g35(n992 ,n34[8] ,n717);
    nand g36(n634 ,n22[4] ,n26[4]);
    nand g37(n6046 ,n6019 ,n6011);
    or g38(n4707 ,n4622 ,n4474);
    nor g39(n2968 ,n2844 ,n2935);
    nor g40(n4144 ,n4069 ,n4112);
    nor g41(n6453 ,n6407 ,n6403);
    nand g42(n479 ,n450 ,n465);
    not g43(n2568 ,n6530);
    xnor g44(n5459 ,n5231 ,n5147);
    not g45(n6068 ,n6062);
    or g46(n791 ,n1517 ,n715);
    nand g47(n811 ,n35[0] ,n712);
    nand g48(n4501 ,n4386 ,n20[7]);
    nand g49(n5844 ,n5806 ,n5783);
    xnor g50(n5184 ,n4897 ,n4586);
    nand g51(n3878 ,n3677 ,n3820);
    not g52(n5611 ,n5610);
    or g53(n3191 ,n3167 ,n3169);
    not g54(n710 ,n712);
    not g55(n3285 ,n3284);
    xnor g56(n4267 ,n4221 ,n4232);
    xnor g57(n2106 ,n2062 ,n2080);
    nand g58(n3524 ,n3464 ,n3478);
    nand g59(n5092 ,n4717 ,n4999);
    xnor g60(n3414 ,n6555 ,n39[6]);
    nand g61(n3603 ,n3462 ,n3481);
    not g62(n1560 ,n1559);
    nand g63(n1736 ,n1584 ,n1700);
    xnor g64(n2616 ,n6526 ,n6531);
    buf g65(n37[6] ,n1506);
    nor g66(n611 ,n33[3] ,n35[3]);
    nand g67(n876 ,n1508 ,n714);
    nor g68(n5588 ,n5401 ,n5448);
    nand g69(n3514 ,n3462 ,n3484);
    nand g70(n6385 ,n6263 ,n6312);
    nand g71(n2057 ,n2000 ,n2056);
    xor g72(n1540 ,n90 ,n94);
    nand g73(n3610 ,n3474 ,n3480);
    nand g74(n4581 ,n4388 ,n20[7]);
    nand g75(n2128 ,n6533 ,n2122);
    nor g76(n4156 ,n4068 ,n4111);
    xnor g77(n2912 ,n2873 ,n2789);
    xnor g78(n4175 ,n4107 ,n4066);
    nand g79(n4136 ,n3995 ,n4072);
    nand g80(n4803 ,n4581 ,n4586);
    dff g81(.RN(n1), .SN(1'b1), .CK(n0), .D(n1293), .Q(n11[10]));
    not g82(n4067 ,n4066);
    or g83(n5745 ,n5648 ,n5663);
    nand g84(n5065 ,n4790 ,n4957);
    nand g85(n2165 ,n6539 ,n2126);
    xnor g86(n4107 ,n4010 ,n3888);
    nor g87(n5373 ,n5122 ,n5291);
    nor g88(n4787 ,n4697 ,n4651);
    xnor g89(n4940 ,n4587 ,n4602);
    dff g90(.RN(n1), .SN(1'b1), .CK(n0), .D(n1241), .Q(n33[2]));
    nand g91(n227 ,n163 ,n152);
    xnor g92(n6036 ,n5960 ,n5856);
    nand g93(n4682 ,n21[7] ,n4378);
    not g94(n2854 ,n2846);
    nand g95(n1277 ,n858 ,n1041);
    xnor g96(n3904 ,n3769 ,n3633);
    nand g97(n5032 ,n4527 ,n4850);
    nand g98(n1008 ,n4[0] ,n557);
    nand g99(n3057 ,n3045 ,n3048);
    nor g100(n3673 ,n3597 ,n3520);
    nand g101(n6042 ,n5987 ,n6008);
    nand g102(n499 ,n473 ,n485);
    xnor g103(n3754 ,n3502 ,n3546);
    nand g104(n4091 ,n3964 ,n4040);
    nor g105(n1675 ,n1644 ,n1652);
    not g106(n3490 ,n36[5]);
    nor g107(n5714 ,n5541 ,n5630);
    or g108(n3193 ,n3165 ,n3180);
    nand g109(n475 ,n413 ,n452);
    nand g110(n3536 ,n3476 ,n19[4]);
    nor g111(n2452 ,n2277 ,n2435);
    xnor g112(n3181 ,n3134 ,n38[11]);
    xnor g113(n5460 ,n5233 ,n5092);
    nand g114(n1106 ,n33[0] ,n555);
    xnor g115(n3135 ,n6573 ,n6550);
    not g116(n219 ,n218);
    nor g117(n5061 ,n4781 ,n4959);
    xnor g118(n1547 ,n32[3] ,n136);
    not g119(n3255 ,n3254);
    nand g120(n2255 ,n2167 ,n2185);
    nand g121(n202 ,n163 ,n157);
    nand g122(n540 ,n525 ,n539);
    nor g123(n3988 ,n3864 ,n3894);
    dff g124(.RN(n1), .SN(1'b1), .CK(n0), .D(n1292), .Q(n1511));
    or g125(n3662 ,n3518 ,n3535);
    nor g126(n2981 ,n2923 ,n2948);
    dff g127(.RN(n1), .SN(1'b1), .CK(n0), .D(n1341), .Q(n33[12]));
    nand g128(n3575 ,n3468 ,n3486);
    nor g129(n6038 ,n5924 ,n6001);
    nand g130(n2143 ,n6539 ,n2121);
    not g131(n2748 ,n2747);
    not g132(n5929 ,n5928);
    nand g133(n5775 ,n5645 ,n5750);
    nand g134(n6471 ,n6317 ,n6387);
    xnor g135(n5865 ,n5801 ,n5616);
    not g136(n2089 ,n21[0]);
    nand g137(n3600 ,n3485 ,n19[3]);
    nand g138(n4348 ,n4347 ,n4336);
    nor g139(n3639 ,n3492 ,n3497);
    nor g140(n838 ,n565 ,n721);
    xnor g141(n6093 ,n6022 ,n6007);
    or g142(n257 ,n189 ,n191);
    nand g143(n2179 ,n6533 ,n2150);
    nand g144(n2349 ,n2288 ,n2293);
    nand g145(n5351 ,n5063 ,n5248);
    xnor g146(n1878 ,n1637 ,n1826);
    nand g147(n4862 ,n4445 ,n4470);
    nand g148(n629 ,n23[7] ,n34[7]);
    xnor g149(n5284 ,n4939 ,n4695);
    xnor g150(n3219 ,n3153 ,n3170);
    nor g151(n2557 ,n2542 ,n2556);
    nor g152(n2643 ,n2566 ,n2587);
    not g153(n1791 ,n1790);
    nor g154(n795 ,n22[0] ,n703);
    nand g155(n3160 ,n3116 ,n3149);
    nand g156(n6071 ,n6018 ,n6044);
    nand g157(n5038 ,n4550 ,n4858);
    xnor g158(n1871 ,n1801 ,n1802);
    nand g159(n4295 ,n4252 ,n4276);
    nor g160(n6461 ,n6421 ,n6418);
    nand g161(n3419 ,n3398 ,n3418);
    nand g162(n825 ,n17[5] ,n721);
    nor g163(n108 ,n24[6] ,n24[5]);
    nand g164(n2200 ,n2096 ,n2157);
    nand g165(n3932 ,n3708 ,n3851);
    xnor g166(n444 ,n418 ,n224);
    not g167(n70 ,n36[0]);
    nand g168(n1281 ,n638 ,n734);
    nor g169(n599 ,n9[1] ,n9[0]);
    nor g170(n785 ,n616 ,n715);
    not g171(n1571 ,n37[3]);
    nand g172(n2582 ,n40[8] ,n6519);
    nand g173(n4328 ,n4318 ,n4310);
    nand g174(n897 ,n24[6] ,n715);
    nor g175(n590 ,n16[6] ,n23[6]);
    nand g176(n3732 ,n3601 ,n3582);
    buf g177(n36[6] ,n1514);
    or g178(n727 ,n710 ,n675);
    nand g179(n2588 ,n40[11] ,n6522);
    nor g180(n4673 ,n4415 ,n4411);
    not g181(n3446 ,n36[2]);
    nand g182(n3859 ,n3660 ,n3804);
    nand g183(n1118 ,n1528 ,n716);
    nor g184(n6230 ,n41[4] ,n6596);
    nand g185(n2283 ,n2118 ,n2238);
    xnor g186(n5532 ,n5302 ,n5152);
    xnor g187(n6002 ,n5915 ,n5852);
    not g188(n293 ,n282);
    nand g189(n984 ,n20[3] ,n714);
    xor g190(n40[4] ,n6607 ,n38[5]);
    nand g191(n1716 ,n1582 ,n1677);
    nand g192(n6014 ,n5953 ,n5986);
    nor g193(n2330 ,n2264 ,n2313);
    nand g194(n6353 ,n6576 ,n6247);
    not g195(n4003 ,n3984);
    xnor g196(n2265 ,n2108 ,n2201);
    nand g197(n6472 ,n6286 ,n6388);
    not g198(n1568 ,n1567);
    xor g199(n4885 ,n4531 ,n4429);
    or g200(n741 ,n717 ,n699);
    nor g201(n660 ,n19[2] ,n27[2]);
    nand g202(n1601 ,n1566 ,n19[0]);
    xor g203(n3768 ,n3614 ,n3542);
    nand g204(n4629 ,n4389 ,n20[0]);
    xnor g205(n6506 ,n3071 ,n3083);
    or g206(n3654 ,n3578 ,n3540);
    nand g207(n3311 ,n3295 ,n3310);
    dff g208(.RN(n1), .SN(1'b1), .CK(n0), .D(n1289), .Q(n1512));
    not g209(n5112 ,n5111);
    nand g210(n983 ,n17[0] ,n721);
    nand g211(n2218 ,n6540 ,n2150);
    nand g212(n5735 ,n5568 ,n5611);
    xnor g213(n6487 ,n38[0] ,n3135);
    xor g214(n6527 ,n3445 ,n19[0]);
    xnor g215(n6562 ,n4332 ,n4352);
    nand g216(n1365 ,n644 ,n754);
    dff g217(.RN(n1), .SN(1'b1), .CK(n0), .D(n1249), .Q(n22[3]));
    nand g218(n1629 ,n1576 ,n1612);
    not g219(n5128 ,n5127);
    nand g220(n3112 ,n38[11] ,n6584);
    nand g221(n1237 ,n1093 ,n782);
    nand g222(n812 ,n34[7] ,n717);
    nand g223(n4586 ,n20[7] ,n4371);
    nand g224(n2100 ,n2079 ,n2074);
    nand g225(n1010 ,n1538 ,n557);
    xnor g226(n1538 ,n98 ,n82);
    nand g227(n4355 ,n4313 ,n4354);
    xnor g228(n3217 ,n3166 ,n3183);
    xor g229(n4225 ,n4171 ,n4200);
    nor g230(n774 ,n615 ,n717);
    not g231(n294 ,n284);
    or g232(n5320 ,n5178 ,n5177);
    nand g233(n4837 ,n4467 ,n4575);
    xnor g234(n3226 ,n38[1] ,n3197);
    xnor g235(n5609 ,n5439 ,n5226);
    nand g236(n6442 ,n6304 ,n6373);
    not g237(n1778 ,n1777);
    nand g238(n196 ,n163 ,n144);
    nand g239(n2049 ,n2048 ,n2036);
    xnor g240(n5634 ,n5420 ,n5225);
    nand g241(n4457 ,n21[6] ,n4376);
    nand g242(n4180 ,n4105 ,n4152);
    not g243(n2783 ,n2782);
    nor g244(n2824 ,n2661 ,n2745);
    xor g245(n6521 ,n6583 ,n6560);
    dff g246(.RN(n1), .SN(1'b1), .CK(n0), .D(n1431), .Q(n25[2]));
    nand g247(n4241 ,n4171 ,n4205);
    or g248(n2578 ,n40[3] ,n6514);
    xnor g249(n2325 ,n2222 ,n2259);
    or g250(n4203 ,n4194 ,n4184);
    nand g251(n6216 ,n6200 ,n6215);
    xnor g252(n4206 ,n4141 ,n4087);
    not g253(n4387 ,n36[0]);
    xnor g254(n2862 ,n2749 ,n2727);
    nand g255(n6122 ,n6069 ,n6102);
    nand g256(n2211 ,n6535 ,n2178);
    xnor g257(n1799 ,n1763 ,n1648);
    nand g258(n2003 ,n1935 ,n1977);
    nand g259(n1410 ,n650 ,n785);
    xnor g260(n4303 ,n4249 ,n4268);
    not g261(n3332 ,n3331);
    nand g262(n2805 ,n2727 ,n2750);
    nand g263(n2195 ,n6533 ,n2149);
    nand g264(n6063 ,n6025 ,n6034);
    nand g265(n3933 ,n3872 ,n3856);
    nand g266(n2132 ,n6537 ,n2123);
    nand g267(n5852 ,n5711 ,n5798);
    nand g268(n860 ,n16[0] ,n714);
    xor g269(n4931 ,n4530 ,n4574);
    nand g270(n958 ,n21[5] ,n714);
    nand g271(n3805 ,n3618 ,n3731);
    not g272(n1582 ,n1581);
    nand g273(n3814 ,n3552 ,n3724);
    nand g274(n4473 ,n21[6] ,n4382);
    nor g275(n4701 ,n4407 ,n4413);
    nor g276(n6448 ,n6386 ,n6385);
    xnor g277(n2260 ,n2203 ,n2109);
    xnor g278(n5414 ,n5176 ,n5173);
    nand g279(n2432 ,n2279 ,n2413);
    xnor g280(n5290 ,n4945 ,n4570);
    xnor g281(n5601 ,n5205 ,n5457);
    nor g282(n2097 ,n2072 ,n2076);
    buf g283(n36[3] ,n1511);
    xnor g284(n460 ,n388 ,n430);
    xnor g285(n4251 ,n4208 ,n4135);
    nor g286(n574 ,n16[2] ,n23[2]);
    not g287(n2705 ,n2704);
    nor g288(n2826 ,n2663 ,n2759);
    buf g289(n37[0] ,n1500);
    dff g290(.RN(n1), .SN(1'b1), .CK(n0), .D(n1301), .Q(n11[5]));
    xnor g291(n6131 ,n6088 ,n6038);
    not g292(n1190 ,n1101);
    nor g293(n779 ,n592 ,n720);
    nand g294(n4543 ,n21[5] ,n4371);
    nand g295(n1395 ,n958 ,n1152);
    xnor g296(n4297 ,n4226 ,n4273);
    nor g297(n2434 ,n2340 ,n2407);
    not g298(n4696 ,n4695);
    nand g299(n3822 ,n3564 ,n3712);
    nor g300(n3792 ,n3577 ,n3687);
    nor g301(n5882 ,n5721 ,n5821);
    or g302(n4727 ,n4481 ,n4432);
    xnor g303(n6195 ,n6177 ,n6174);
    xnor g304(n5509 ,n5402 ,n5288);
    nor g305(n2772 ,n2641 ,n2683);
    nand g306(n1128 ,n33[4] ,n555);
    nand g307(n244 ,n163 ,n150);
    nand g308(n4636 ,n21[4] ,n4380);
    nand g309(n3107 ,n38[2] ,n6575);
    nand g310(n1030 ,n12[3] ,n710);
    nand g311(n874 ,n33[8] ,n554);
    nand g312(n6212 ,n6211 ,n6198);
    nand g313(n1328 ,n992 ,n1083);
    not g314(n1822 ,n1821);
    nand g315(n5577 ,n5317 ,n5477);
    nand g316(n4281 ,n4209 ,n4268);
    or g317(n4035 ,n3912 ,n4007);
    nand g318(n6366 ,n6505 ,n6249);
    not g319(n554 ,n555);
    nand g320(n929 ,n29[5] ,n721);
    not g321(n5827 ,n5826);
    xnor g322(n5884 ,n5758 ,n5808);
    nand g323(n455 ,n399 ,n431);
    not g324(n168 ,n36[5]);
    nand g325(n4575 ,n21[4] ,n4386);
    xnor g326(n2856 ,n2760 ,n2786);
    nand g327(n3370 ,n3319 ,n3369);
    nand g328(n6346 ,n38[2] ,n6246);
    xnor g329(n1775 ,n1636 ,n1729);
    nor g330(n1484 ,n578 ,n1199);
    nor g331(n3843 ,n3673 ,n3802);
    nor g332(n4659 ,n4409 ,n4416);
    xnor g333(n3128 ,n6578 ,n6555);
    nand g334(n6363 ,n6499 ,n6249);
    nand g335(n473 ,n401 ,n455);
    nand g336(n6282 ,n6570 ,n6254);
    nand g337(n1388 ,n640 ,n779);
    nand g338(n1400 ,n963 ,n1156);
    nand g339(n2137 ,n6538 ,n2122);
    nand g340(n6331 ,n6575 ,n6247);
    nand g341(n1350 ,n904 ,n1103);
    xnor g342(n358 ,n311 ,n185);
    xnor g343(n6505 ,n3052 ,n3081);
    nand g344(n1301 ,n1057 ,n806);
    nand g345(n1188 ,n8[1] ,n713);
    nand g346(n5068 ,n4734 ,n4986);
    xnor g347(n5958 ,n5868 ,n5876);
    nand g348(n4213 ,n4137 ,n4182);
    nand g349(n5507 ,n5254 ,n5366);
    xnor g350(n3218 ,n3161 ,n3174);
    nand g351(n1440 ,n983 ,n1253);
    or g352(n4732 ,n4566 ,n4476);
    nand g353(n5664 ,n5581 ,n5573);
    nor g354(n1990 ,n1913 ,n1975);
    nand g355(n1362 ,n912 ,n1114);
    xnor g356(n3025 ,n2971 ,n2955);
    nand g357(n763 ,n724 ,n696);
    not g358(n4393 ,n21[1]);
    nor g359(n607 ,n23[7] ,n34[7]);
    nor g360(n773 ,n607 ,n717);
    nand g361(n4309 ,n4259 ,n4295);
    nor g362(n115 ,n32[2] ,n32[0]);
    nand g363(n1490 ,n722 ,n1484);
    nand g364(n796 ,n557 ,n705);
    xnor g365(n426 ,n390 ,n389);
    nand g366(n1058 ,n11[4] ,n711);
    xnor g367(n448 ,n392 ,n374);
    dff g368(.RN(n1), .SN(1'b1), .CK(n0), .D(n1322), .Q(n34[12]));
    xor g369(n6523 ,n6585 ,n6562);
    nand g370(n1694 ,n1584 ,n1654);
    nor g371(n1838 ,n1776 ,n1822);
    nand g372(n5508 ,n5258 ,n5341);
    nand g373(n3320 ,n6585 ,n41[12]);
    xnor g374(n5415 ,n5211 ,n5160);
    nand g375(n946 ,n27[15] ,n715);
    nand g376(n4618 ,n4384 ,n20[1]);
    xnor g377(n4248 ,n4206 ,n4192);
    xnor g378(n522 ,n495 ,n458);
    xnor g379(n699 ,n23[1] ,n34[1]);
    or g380(n3063 ,n3028 ,n3039);
    or g381(n1488 ,n720 ,n1483);
    nand g382(n4606 ,n4376 ,n20[6]);
    not g383(n5518 ,n5517);
    nand g384(n6052 ,n5979 ,n6014);
    nor g385(n3392 ,n6553 ,n39[4]);
    nand g386(n6475 ,n6363 ,n6429);
    not g387(n4436 ,n4435);
    nand g388(n1710 ,n1582 ,n1675);
    buf g389(n14[12], n11[12]);
    nand g390(n4214 ,n4196 ,n4183);
    nand g391(n6311 ,n6494 ,n6253);
    nand g392(n1311 ,n1069 ,n957);
    nand g393(n6047 ,n5967 ,n6007);
    xnor g394(n6030 ,n5961 ,n5853);
    nand g395(n5462 ,n5252 ,n5400);
    or g396(n752 ,n555 ,n684);
    nand g397(n467 ,n433 ,n445);
    nor g398(n2435 ,n2278 ,n2410);
    nor g399(n2800 ,n2657 ,n2677);
    nor g400(n2899 ,n2817 ,n2882);
    nor g401(n4981 ,n4436 ,n4787);
    xnor g402(n531 ,n507 ,n512);
    nand g403(n1196 ,n1072 ,n950);
    xor g404(n1612 ,n1566 ,n19[0]);
    nand g405(n631 ,n33[12] ,n35[12]);
    xnor g406(n5597 ,n5168 ,n5455);
    nand g407(n947 ,n27[14] ,n715);
    nand g408(n4838 ,n4492 ,n4434);
    xnor g409(n4173 ,n4136 ,n4103);
    xnor g410(n3000 ,n2918 ,n2967);
    not g411(n5619 ,n5618);
    nand g412(n5138 ,n4773 ,n5051);
    nand g413(n5737 ,n5687 ,n5624);
    nand g414(n3085 ,n3059 ,n3084);
    xnor g415(n3132 ,n6580 ,n6557);
    nand g416(n1623 ,n1582 ,n1612);
    nor g417(n4785 ,n4556 ,n4545);
    or g418(n733 ,n717 ,n667);
    nand g419(n352 ,n254 ,n327);
    xnor g420(n5873 ,n5772 ,n5756);
    nand g421(n4085 ,n3960 ,n4036);
    not g422(n62 ,n36[6]);
    nor g423(n2641 ,n2566 ,n2582);
    xnor g424(n2286 ,n2118 ,n2244);
    nand g425(n5371 ,n5152 ,n5242);
    buf g426(n14[7], n10[7]);
    xnor g427(n2105 ,n2064 ,n2078);
    nand g428(n3075 ,n3044 ,n3074);
    not g429(n3466 ,n3465);
    nand g430(n5966 ,n5900 ,n5919);
    xnor g431(n6548 ,n3335 ,n3384);
    not g432(n149 ,n37[5]);
    xor g433(n6024 ,n5972 ,n5993);
    nand g434(n6102 ,n6073 ,n6067);
    or g435(n747 ,n717 ,n690);
    or g436(n744 ,n717 ,n665);
    nand g437(n1684 ,n1579 ,n1655);
    nand g438(n3009 ,n2945 ,n2980);
    nand g439(n6300 ,n6561 ,n6251);
    nand g440(n3137 ,n38[7] ,n3098);
    nor g441(n2333 ,n2119 ,n2294);
    nand g442(n1235 ,n1032 ,n731);
    nand g443(n5867 ,n5797 ,n5836);
    buf g444(n37[1] ,n1501);
    nand g445(n1322 ,n883 ,n1078);
    nand g446(n875 ,n1509 ,n714);
    or g447(n5665 ,n5588 ,n5559);
    xnor g448(n1553 ,n24[4] ,n126);
    nor g449(n6253 ,n6227 ,n6224);
    xnor g450(n3003 ,n2957 ,n2929);
    nand g451(n998 ,n8[0] ,n713);
    nand g452(n895 ,n33[0] ,n712);
    nor g453(n600 ,n21[1] ,n30[1]);
    nand g454(n5809 ,n5677 ,n5745);
    nand g455(n944 ,n24[2] ,n715);
    xor g456(n5861 ,n5780 ,n5757);
    nand g457(n6424 ,n6287 ,n6355);
    nand g458(n3876 ,n3662 ,n3825);
    nand g459(n4676 ,n20[3] ,n4369);
    or g460(n3061 ,n3029 ,n3038);
    xor g461(n4928 ,n4667 ,n4423);
    nand g462(n1004 ,n1537 ,n557);
    xnor g463(n4052 ,n3935 ,n3969);
    or g464(n4771 ,n4602 ,n4587);
    xnor g465(n3784 ,n3619 ,n3612);
    nor g466(n3011 ,n2958 ,n2976);
    not g467(n4960 ,n4959);
    xor g468(n4908 ,n4650 ,n4421);
    nand g469(n1036 ,n2[6] ,n557);
    xnor g470(n3749 ,n3600 ,n3515);
    nor g471(n2606 ,n2567 ,n2596);
    xnor g472(n361 ,n296 ,n314);
    nand g473(n1018 ,n1539 ,n557);
    xnor g474(n2021 ,n1973 ,n1991);
    nand g475(n3161 ,n3117 ,n3148);
    nor g476(n1545 ,n140 ,n142);
    nor g477(n2730 ,n2567 ,n2626);
    nand g478(n1293 ,n1047 ,n871);
    nand g479(n1705 ,n1580 ,n1677);
    nand g480(n1299 ,n876 ,n1055);
    nand g481(n6193 ,n6171 ,n6185);
    not g482(n3155 ,n3154);
    xnor g483(n2928 ,n2869 ,n2770);
    nor g484(n2392 ,n2307 ,n2359);
    nand g485(n5976 ,n5902 ,n5945);
    not g486(n3488 ,n36[2]);
    xnor g487(n2310 ,n2119 ,n2240);
    dff g488(.RN(n1), .SN(1'b1), .CK(n0), .D(n1375), .Q(n30[7]));
    not g489(n2676 ,n2675);
    nand g490(n6315 ,n38[6] ,n6246);
    nor g491(n2700 ,n2565 ,n2632);
    dff g492(.RN(n1), .SN(1'b1), .CK(n0), .D(n1474), .Q(n27[2]));
    nor g493(n569 ,n34[5] ,n34[6]);
    nor g494(n594 ,n31[1] ,n35[1]);
    not g495(n66 ,n36[5]);
    nor g496(n2642 ,n2566 ,n2584);
    xnor g497(n6508 ,n3049 ,n3087);
    nor g498(n2702 ,n2567 ,n2623);
    nand g499(n4470 ,n4380 ,n20[0]);
    nand g500(n6320 ,n6546 ,n6248);
    xnor g501(n4286 ,n4248 ,n4246);
    nand g502(n110 ,n24[4] ,n109);
    nand g503(n4989 ,n4646 ,n4852);
    or g504(n3650 ,n3609 ,n3602);
    nand g505(n5090 ,n4722 ,n5052);
    nand g506(n5399 ,n5284 ,n5287);
    nand g507(n3074 ,n3041 ,n3073);
    nand g508(n3045 ,n2996 ,n3022);
    xnor g509(n5962 ,n5873 ,n5909);
    nand g510(n1061 ,n11[2] ,n711);
    nor g511(n2684 ,n2566 ,n2617);
    nor g512(n1971 ,n1924 ,n1953);
    not g513(n4400 ,n21[0]);
    not g514(n310 ,n309);
    nand g515(n4555 ,n21[6] ,n4373);
    xnor g516(n3745 ,n3506 ,n3588);
    xnor g517(n495 ,n463 ,n447);
    nand g518(n4466 ,n21[7] ,n4380);
    xnor g519(n3753 ,n3534 ,n3509);
    nand g520(n4666 ,n21[6] ,n4371);
    nand g521(n6417 ,n6310 ,n6346);
    nand g522(n1711 ,n1580 ,n1676);
    nand g523(n6347 ,n39[2] ,n6248);
    nand g524(n6050 ,n6015 ,n5974);
    nor g525(n3424 ,n3414 ,n3423);
    nand g526(n1397 ,n959 ,n1153);
    nor g527(n3685 ,n3622 ,n3610);
    nand g528(n4675 ,n21[7] ,n4371);
    xnor g529(n5300 ,n5136 ,n5124);
    nor g530(n2779 ,n2640 ,n2694);
    nand g531(n1019 ,n1531 ,n716);
    nand g532(n2945 ,n2827 ,n2926);
    or g533(n781 ,n720 ,n671);
    nand g534(n5382 ,n5178 ,n5177);
    nor g535(n4070 ,n3965 ,n4032);
    or g536(n524 ,n507 ,n512);
    nor g537(n6257 ,n6233 ,n6252);
    xnor g538(n5973 ,n5861 ,n5832);
    nand g539(n551 ,n487 ,n550);
    not g540(n3486 ,n3488);
    dff g541(.RN(n1), .SN(1'b1), .CK(n0), .D(n1448), .Q(n12[1]));
    nor g542(n783 ,n580 ,n715);
    xnor g543(n1831 ,n1771 ,n1645);
    nor g544(n6447 ,n6424 ,n6423);
    not g545(n4663 ,n4662);
    xnor g546(n3916 ,n3777 ,n3733);
    nand g547(n2628 ,n2587 ,n2578);
    or g548(n4744 ,n4574 ,n4468);
    or g549(n5241 ,n5118 ,n5107);
    nor g550(n2965 ,n2881 ,n2941);
    nand g551(n2623 ,n2593 ,n2572);
    nor g552(n2044 ,n2043 ,n2017);
    not g553(n171 ,n36[2]);
    xnor g554(n4051 ,n3973 ,n3902);
    nand g555(n1887 ,n1757 ,n1862);
    nand g556(n1498 ,n1481 ,n1497);
    nor g557(n2698 ,n2568 ,n2626);
    nand g558(n1133 ,n17[7] ,n722);
    xnor g559(n4971 ,n4606 ,n4466);
    xor g560(n6511 ,n6573 ,n6550);
    nor g561(n3558 ,n3489 ,n3498);
    nor g562(n4204 ,n4156 ,n4186);
    xnor g563(n3180 ,n3127 ,n38[6]);
    xnor g564(n2302 ,n2120 ,n2241);
    buf g565(n14[1], n11[1]);
    xnor g566(n297 ,n220 ,n221);
    not g567(n3498 ,n19[4]);
    nand g568(n456 ,n416 ,n435);
    nand g569(n4609 ,n4380 ,n20[6]);
    xor g570(n4899 ,n4507 ,n4578);
    xnor g571(n296 ,n189 ,n191);
    nand g572(n1375 ,n914 ,n1126);
    xnor g573(n3940 ,n3766 ,n3578);
    xnor g574(n5763 ,n5644 ,n5578);
    xnor g575(n421 ,n361 ,n363);
    nand g576(n96 ,n80 ,n95);
    nand g577(n1742 ,n1662 ,n1706);
    not g578(n3269 ,n3268);
    xnor g579(n3906 ,n3752 ,n3615);
    not g580(n4364 ,n37[5]);
    dff g581(.RN(n1), .SN(1'b1), .CK(n0), .D(n1482), .Q(n29[6]));
    nand g582(n77 ,n71 ,n53);
    not g583(n2567 ,n6527);
    nand g584(n982 ,n27[1] ,n715);
    or g585(n787 ,n717 ,n668);
    nand g586(n5977 ,n5857 ,n5939);
    nand g587(n1341 ,n1146 ,n954);
    nand g588(n3235 ,n3207 ,n3234);
    xor g589(n2059 ,n2283 ,n2273);
    nand g590(n5063 ,n4791 ,n4956);
    xnor g591(n4011 ,n3893 ,n3864);
    nand g592(n1234 ,n1027 ,n789);
    nand g593(n3308 ,n3292 ,n3307);
    nand g594(n2469 ,n2411 ,n2446);
    xnor g595(n5168 ,n4904 ,n4498);
    xnor g596(n1933 ,n1870 ,n1808);
    not g597(n2396 ,n2397);
    nand g598(n2235 ,n2145 ,n2217);
    not g599(n1903 ,n1904);
    xnor g600(n5595 ,n5180 ,n5461);
    xnor g601(n4010 ,n3887 ,n3911);
    nand g602(n5126 ,n4737 ,n5049);
    xnor g603(n2939 ,n2879 ,n2800);
    xnor g604(n335 ,n202 ,n236);
    nand g605(n506 ,n468 ,n483);
    or g606(n4147 ,n4136 ,n4103);
    nand g607(n2180 ,n6535 ,n2149);
    nand g608(n1182 ,n29[3] ,n724);
    nand g609(n3712 ,n3604 ,n3511);
    or g610(n4102 ,n4027 ,n4055);
    xnor g611(n4298 ,n4230 ,n4274);
    xnor g612(n5158 ,n4923 ,n4486);
    nand g613(n4563 ,n21[4] ,n4363);
    nor g614(n2689 ,n2566 ,n2632);
    nor g615(n1908 ,n1836 ,n1888);
    nand g616(n5922 ,n5785 ,n5878);
    dff g617(.RN(n1), .SN(1'b1), .CK(n0), .D(n1430), .Q(n26[0]));
    nand g618(n4088 ,n3958 ,n4042);
    nand g619(n4490 ,n21[0] ,n4380);
    nand g620(n2001 ,n1965 ,n1979);
    xnor g621(n2320 ,n2119 ,n2252);
    xnor g622(n2125 ,n2109 ,n2088);
    xnor g623(n2309 ,n2254 ,n2119);
    nand g624(n5086 ,n4726 ,n4991);
    nand g625(n4336 ,n4315 ,n4326);
    nand g626(n4502 ,n21[3] ,n4384);
    nand g627(n1766 ,n1681 ,n1738);
    or g628(n4794 ,n4642 ,n4464);
    nand g629(n2244 ,n2141 ,n2195);
    not g630(n2313 ,n2312);
    nor g631(n4086 ,n3956 ,n4034);
    nor g632(n2464 ,n2275 ,n2433);
    xnor g633(n389 ,n299 ,n270);
    nand g634(n1013 ,n10[0] ,n555);
    nand g635(n3559 ,n3470 ,n3485);
    nor g636(n2457 ,n2437 ,n2427);
    nand g637(n3290 ,n3273 ,n3259);
    not g638(n4368 ,n37[2]);
    nand g639(n4124 ,n3971 ,n4080);
    xnor g640(n302 ,n193 ,n217);
    nand g641(n3930 ,n3522 ,n3846);
    nand g642(n6322 ,n6585 ,n6247);
    nand g643(n332 ,n238 ,n280);
    nand g644(n2242 ,n2135 ,n2188);
    nand g645(n3059 ,n3032 ,n3037);
    nor g646(n4667 ,n4409 ,n4406);
    or g647(n746 ,n715 ,n676);
    nor g648(n754 ,n602 ,n720);
    xnor g649(n4299 ,n4271 ,n4218);
    nand g650(n327 ,n240 ,n276);
    or g651(n500 ,n473 ,n485);
    nand g652(n4997 ,n4674 ,n4870);
    not g653(n2920 ,n2919);
    xnor g654(n5762 ,n5643 ,n5532);
    nor g655(n3030 ,n2997 ,n3018);
    xnor g656(n2303 ,n2232 ,n2230);
    nand g657(n1407 ,n655 ,n784);
    not g658(n5971 ,n5970);
    not g659(n4514 ,n4513);
    nand g660(n6098 ,n6016 ,n6059);
    nand g661(n4043 ,n3927 ,n3993);
    nand g662(n6439 ,n6301 ,n6374);
    nand g663(n542 ,n528 ,n541);
    nor g664(n2150 ,n2115 ,n2122);
    not g665(n113 ,n32[7]);
    nand g666(n328 ,n209 ,n277);
    not g667(n3475 ,n36[7]);
    nand g668(n1670 ,n1582 ,n1649);
    nor g669(n2233 ,n2136 ,n2214);
    xnor g670(n3901 ,n3761 ,n3529);
    nand g671(n6276 ,n6569 ,n6254);
    nand g672(n5101 ,n4728 ,n4983);
    nand g673(n5051 ,n4681 ,n4851);
    nor g674(n2814 ,n2673 ,n2779);
    nand g675(n4045 ,n3929 ,n3998);
    nand g676(n2907 ,n2825 ,n2891);
    not g677(n2262 ,n2261);
    not g678(n159 ,n158);
    or g679(n3982 ,n3858 ,n3908);
    or g680(n4118 ,n3971 ,n4080);
    nand g681(n4849 ,n4483 ,n4595);
    xor g682(n5422 ,n5177 ,n5294);
    nor g683(n4077 ,n3884 ,n4023);
    nand g684(n3378 ,n3325 ,n3377);
    xor g685(n1541 ,n86 ,n77);
    nor g686(n583 ,n34[13] ,n34[14]);
    dff g687(.RN(n1), .SN(1'b1), .CK(n0), .D(n1408), .Q(n21[0]));
    xnor g688(n2272 ,n2204 ,n2118);
    xnor g689(n4264 ,n4193 ,n4231);
    nand g690(n3587 ,n3464 ,n3481);
    not g691(n4411 ,n20[2]);
    nand g692(n4680 ,n21[3] ,n4388);
    dff g693(.RN(n1), .SN(1'b1), .CK(n0), .D(n1443), .Q(n12[10]));
    nor g694(n6144 ,n6138 ,n6105);
    nand g695(n5380 ,n5160 ,n5211);
    nand g696(n325 ,n283 ,n270);
    nand g697(n2191 ,n6537 ,n2149);
    nand g698(n4813 ,n4618 ,n4427);
    nand g699(n918 ,n30[5] ,n723);
    nand g700(n1436 ,n930 ,n1210);
    or g701(n3194 ,n3160 ,n3171);
    dff g702(.RN(n1), .SN(1'b1), .CK(n0), .D(n1308), .Q(n10[14]));
    not g703(n3866 ,n3865);
    not g704(n4371 ,n4370);
    nand g705(n2625 ,n2594 ,n2579);
    nand g706(n6051 ,n5942 ,n6012);
    nand g707(n6118 ,n6107 ,n6063);
    nand g708(n855 ,n16[2] ,n714);
    nand g709(n1325 ,n934 ,n1080);
    nand g710(n547 ,n520 ,n546);
    nand g711(n1338 ,n1090 ,n956);
    nand g712(n3599 ,n3464 ,n3480);
    nand g713(n93 ,n77 ,n87);
    nand g714(n5251 ,n4793 ,n5067);
    nand g715(n2548 ,n2511 ,n2547);
    nand g716(n5142 ,n4794 ,n5019);
    nand g717(n1062 ,n11[1] ,n711);
    nand g718(n4089 ,n3982 ,n4031);
    nand g719(n5755 ,n5514 ,n5685);
    nand g720(n4645 ,n20[0] ,n4367);
    not g721(n2757 ,n2756);
    dff g722(.RN(n1), .SN(1'b1), .CK(n0), .D(n1325), .Q(n34[10]));
    xnor g723(n6088 ,n6031 ,n5966);
    not g724(n4529 ,n4528);
    nand g725(n418 ,n253 ,n381);
    nand g726(n5495 ,n5259 ,n5348);
    nand g727(n2532 ,n2514 ,n2490);
    nand g728(n6310 ,n6567 ,n6254);
    nand g729(n1042 ,n11[13] ,n711);
    dff g730(.RN(n1), .SN(1'b1), .CK(n0), .D(n1339), .Q(n24[3]));
    not g731(n1776 ,n1775);
    nand g732(n3167 ,n3110 ,n3144);
    xor g733(n4910 ,n4665 ,n4494);
    not g734(n3477 ,n36[3]);
    nand g735(n4211 ,n4150 ,n4190);
    nand g736(n1450 ,n832 ,n1333);
    nor g737(n784 ,n590 ,n715);
    or g738(n2354 ,n2317 ,n2286);
    nand g739(n3511 ,n3485 ,n19[1]);
    not g740(n4362 ,n37[6]);
    or g741(n4262 ,n4193 ,n4231);
    nor g742(n1591 ,n1572 ,n19[3]);
    nand g743(n6334 ,n6487 ,n6253);
    or g744(n254 ,n213 ,n214);
    dff g745(.RN(n1), .SN(1'b1), .CK(n0), .D(n1373), .Q(n23[2]));
    nand g746(n3796 ,n3561 ,n3703);
    or g747(n4163 ,n4100 ,n4115);
    nand g748(n4352 ,n4351 ,n4340);
    xnor g749(n1607 ,n1564 ,n19[4]);
    or g750(n4729 ,n4619 ,n4421);
    xnor g751(n4932 ,n4621 ,n4422);
    dff g752(.RN(n1), .SN(1'b1), .CK(n0), .D(n1480), .Q(n17[6]));
    nand g753(n2994 ,n2938 ,n2953);
    nor g754(n2597 ,n2565 ,n2586);
    nand g755(n280 ,n190 ,n181);
    xor g756(n6520 ,n6582 ,n6559);
    nand g757(n3087 ,n3061 ,n3086);
    nand g758(n1291 ,n1046 ,n870);
    dff g759(.RN(n1), .SN(1'b1), .CK(n0), .D(n1226), .Q(n27[3]));
    nand g760(n5264 ,n4979 ,n5094);
    xnor g761(n4249 ,n4209 ,n4219);
    nand g762(n5015 ,n4507 ,n4842);
    xnor g763(n1924 ,n1876 ,n1817);
    nand g764(n3716 ,n3598 ,n3593);
    not g765(n4004 ,n3985);
    nand g766(n4098 ,n4027 ,n4055);
    nand g767(n1430 ,n803 ,n1185);
    xnor g768(n5196 ,n4944 ,n4463);
    not g769(n4537 ,n4536);
    xnor g770(n6576 ,n1920 ,n1915);
    nand g771(n1411 ,n977 ,n1168);
    nand g772(n1283 ,n863 ,n1036);
    nand g773(n857 ,n1500 ,n714);
    nand g774(n5261 ,n5070 ,n5080);
    nand g775(n129 ,n24[5] ,n127);
    or g776(n739 ,n717 ,n666);
    nor g777(n2647 ,n2566 ,n2592);
    or g778(n253 ,n180 ,n222);
    nand g779(n864 ,n1513 ,n556);
    nand g780(n2098 ,n2078 ,n2081);
    nand g781(n5067 ,n4777 ,n5002);
    nand g782(n1258 ,n842 ,n1000);
    nor g783(n2601 ,n2567 ,n2592);
    nand g784(n3879 ,n3693 ,n3809);
    nand g785(n224 ,n159 ,n144);
    nand g786(n518 ,n481 ,n504);
    or g787(n5490 ,n5225 ,n5413);
    not g788(n71 ,n70);
    not g789(n1825 ,n1824);
    nor g790(n2384 ,n2302 ,n2363);
    nand g791(n648 ,n33[11] ,n35[11]);
    nand g792(n2225 ,n2131 ,n2183);
    nand g793(n5801 ,n5657 ,n5746);
    xnor g794(n41[5] ,n6109 ,n6124);
    xnor g795(n5440 ,n5159 ,n5140);
    nand g796(n2182 ,n6536 ,n2149);
    nand g797(n4217 ,n4199 ,n4180);
    or g798(n2350 ,n2288 ,n2293);
    nand g799(n2190 ,n6535 ,n2148);
    not g800(n5613 ,n5612);
    nor g801(n2719 ,n2565 ,n2621);
    xnor g802(n5647 ,n5416 ,n5405);
    not g803(n49 ,n48);
    nand g804(n1358 ,n1112 ,n890);
    xnor g805(n3133 ,n6560 ,n6583);
    nand g806(n3864 ,n3652 ,n3807);
    not g807(n1849 ,n1841);
    xnor g808(n6023 ,n5976 ,n5912);
    nor g809(n2706 ,n2567 ,n2632);
    nand g810(n4868 ,n4462 ,n4620);
    nor g811(n337 ,n269 ,n310);
    nand g812(n1715 ,n1586 ,n1675);
    nand g813(n1319 ,n921 ,n1099);
    not g814(n717 ,n718);
    xnor g815(n3762 ,n3538 ,n3505);
    xnor g816(n6188 ,n6158 ,n6156);
    xnor g817(n85 ,n59 ,n43);
    nand g818(n1349 ,n903 ,n1098);
    or g819(n5243 ,n5121 ,n5120);
    or g820(n5273 ,n5081 ,n5125);
    nand g821(n4274 ,n4243 ,n4260);
    not g822(n663 ,n662);
    nand g823(n867 ,n33[12] ,n712);
    or g824(n726 ,n715 ,n688);
    xor g825(n39[5] ,n6613 ,n38[5]);
    nand g826(n5118 ,n4760 ,n5030);
    nand g827(n6009 ,n5952 ,n5985);
    nand g828(n6327 ,n38[12] ,n6246);
    xnor g829(n5835 ,n5690 ,n5498);
    nand g830(n6430 ,n6243 ,n6261);
    nor g831(n2554 ,n2553 ,n2540);
    nand g832(n5391 ,n5213 ,n5212);
    nand g833(n5504 ,n5268 ,n5368);
    nand g834(n941 ,n28[2] ,n717);
    nand g835(n645 ,n33[9] ,n35[9]);
    nand g836(n1053 ,n2[1] ,n557);
    nor g837(n2764 ,n2642 ,n2726);
    nor g838(n2799 ,n2637 ,n2678);
    nand g839(n1385 ,n628 ,n774);
    dff g840(.RN(n1), .SN(1'b1), .CK(n0), .D(n1409), .Q(n20[7]));
    nand g841(n1074 ,n10[6] ,n555);
    xnor g842(n2373 ,n2310 ,n2268);
    xnor g843(n5309 ,n5121 ,n5120);
    nor g844(n2615 ,n2565 ,n2582);
    nand g845(n6155 ,n6076 ,n6134);
    nand g846(n4668 ,n20[0] ,n4365);
    or g847(n2352 ,n2296 ,n2291);
    nand g848(n5898 ,n5823 ,n5852);
    nand g849(n4642 ,n21[5] ,n4361);
    nand g850(n4254 ,n4203 ,n4233);
    nand g851(n1086 ,n1550 ,n716);
    nand g852(n5021 ,n4503 ,n4862);
    or g853(n4762 ,n4490 ,n4454);
    xnor g854(n1946 ,n1904 ,n1905);
    xnor g855(n2284 ,n2232 ,n2234);
    nand g856(n765 ,n724 ,n694);
    not g857(n4376 ,n4375);
    xnor g858(n2369 ,n2290 ,n2308);
    nor g859(n3393 ,n6557 ,n6542);
    xnor g860(n1548 ,n32[2] ,n134);
    nor g861(n2654 ,n2565 ,n2592);
    nor g862(n2497 ,n2405 ,n2474);
    nor g863(n5662 ,n5577 ,n5538);
    nor g864(n756 ,n591 ,n720);
    dff g865(.RN(n1), .SN(1'b1), .CK(n0), .D(n1321), .Q(n34[13]));
    xnor g866(n5931 ,n5819 ,n5755);
    nor g867(n3943 ,n3791 ,n3840);
    nand g868(n4847 ,n4486 ,n4475);
    xnor g869(n4174 ,n4079 ,n4137);
    nor g870(n613 ,n17[6] ,n17[7]);
    xor g871(n3750 ,n3642 ,n3510);
    nand g872(n4564 ,n21[0] ,n4367);
    nor g873(n2932 ,n2834 ,n2899);
    xnor g874(n3197 ,n3151 ,n6551);
    nor g875(n133 ,n32[1] ,n32[0]);
    nand g876(n3816 ,n3557 ,n3709);
    xnor g877(n4058 ,n3949 ,n3889);
    nand g878(n2504 ,n2430 ,n2477);
    xnor g879(n424 ,n367 ,n342);
    nor g880(n6115 ,n6068 ,n6091);
    nor g881(n2669 ,n2568 ,n2585);
    xnor g882(n5171 ,n4880 ,n4668);
    nand g883(n233 ,n167 ,n150);
    xnor g884(n2954 ,n2859 ,n2902);
    nand g885(n4306 ,n4275 ,n4289);
    nor g886(n5651 ,n5549 ,n5525);
    or g887(n521 ,n513 ,n511);
    nand g888(n1321 ,n878 ,n1077);
    xnor g889(n4063 ,n3950 ,n3879);
    nand g890(n4815 ,n4593 ,n4431);
    nand g891(n4819 ,n4460 ,n4571);
    nand g892(n4513 ,n20[2] ,n4371);
    xnor g893(n2872 ,n2793 ,n2730);
    nor g894(n5323 ,n5082 ,n5189);
    nand g895(n6081 ,n6013 ,n6050);
    xnor g896(n6145 ,n6108 ,n6114);
    not g897(n111 ,n110);
    nand g898(n411 ,n363 ,n361);
    or g899(n788 ,n715 ,n709);
    not g900(n47 ,n46);
    nand g901(n1037 ,n12[0] ,n711);
    nand g902(n78 ,n61 ,n47);
    not g903(n6028 ,n6027);
    nand g904(n4161 ,n3944 ,n4125);
    nand g905(n3798 ,n3574 ,n3696);
    nand g906(n4651 ,n21[7] ,n4374);
    nand g907(n3210 ,n3166 ,n3183);
    nand g908(n5135 ,n4707 ,n5040);
    not g909(n2060 ,n6538);
    nor g910(n571 ,n21[7] ,n30[7]);
    not g911(n4584 ,n4583);
    or g912(n5349 ,n5187 ,n5186);
    nand g913(n1863 ,n1751 ,n1798);
    nand g914(n1487 ,n722 ,n1485);
    nand g915(n4809 ,n4642 ,n4464);
    or g916(n6178 ,n6155 ,n6166);
    nor g917(n2481 ,n2434 ,n2457);
    xnor g918(n3151 ,n6574 ,n3120);
    nand g919(n4304 ,n4296 ,n4287);
    nand g920(n1626 ,n1616 ,n1604);
    nand g921(n1120 ,n31[4] ,n720);
    xnor g922(n5227 ,n4974 ,n4686);
    nand g923(n1686 ,n1577 ,n1655);
    nand g924(n3842 ,n3648 ,n3806);
    not g925(n4408 ,n20[1]);
    not g926(n4685 ,n4684);
    nand g927(n380 ,n288 ,n341);
    xnor g928(n3125 ,n6563 ,n6586);
    or g929(n2445 ,n2377 ,n2422);
    xnor g930(n2124 ,n2110 ,n2063);
    nand g931(n2966 ,n2903 ,n2936);
    not g932(n2624 ,n2625);
    nand g933(n5074 ,n4743 ,n4982);
    xnor g934(n2374 ,n2300 ,n2264);
    nor g935(n2969 ,n2833 ,n2937);
    not g936(n4059 ,n4058);
    nand g937(n6425 ,n6288 ,n6354);
    not g938(n3279 ,n3278);
    xnor g939(n2031 ,n1993 ,n2020);
    or g940(n2036 ,n2018 ,n2024);
    nand g941(n955 ,n35[13] ,n712);
    xnor g942(n4911 ,n4607 ,n4643);
    nand g943(n5589 ,n5344 ,n5480);
    xor g944(n4943 ,n4553 ,n4582);
    nor g945(n3437 ,n3397 ,n3436);
    not g946(n208 ,n207);
    nand g947(n3789 ,n3606 ,n3690);
    xnor g948(n6601 ,n3412 ,n3431);
    nand g949(n3696 ,n3609 ,n3602);
    nand g950(n2112 ,n2086 ,n2104);
    nand g951(n6222 ,n25[2] ,n6225);
    xnor g952(n2867 ,n2758 ,n2663);
    xnor g953(n3748 ,n3541 ,n3545);
    nand g954(n2621 ,n2595 ,n2573);
    xor g955(n1530 ,n423 ,n420);
    nand g956(n1363 ,n1049 ,n913);
    nand g957(n102 ,n81 ,n101);
    xor g958(n3742 ,n3613 ,n3585);
    xnor g959(n1613 ,n19[1] ,n1574);
    nand g960(n3250 ,n3189 ,n3249);
    nand g961(n823 ,n23[0] ,n715);
    nand g962(n919 ,n33[1] ,n712);
    nor g963(n2986 ,n2916 ,n2951);
    xnor g964(n5185 ,n4925 ,n4630);
    xor g965(n4886 ,n4523 ,n4474);
    nand g966(n5659 ,n5526 ,n5535);
    or g967(n6078 ,n5990 ,n6036);
    nand g968(n1919 ,n1859 ,n1895);
    nor g969(n576 ,n26[3] ,n26[4]);
    nand g970(n1760 ,n1669 ,n1717);
    nand g971(n1022 ,n12[6] ,n710);
    xnor g972(n4183 ,n4096 ,n4057);
    nor g973(n6469 ,n6443 ,n6441);
    xnor g974(n2495 ,n2444 ,n2419);
    xnor g975(n5207 ,n4908 ,n4619);
    not g976(n5933 ,n5923);
    nand g977(n3014 ,n2943 ,n2985);
    nor g978(n3840 ,n3792 ,n3787);
    nand g979(n4620 ,n20[5] ,n4367);
    nand g980(n5296 ,n4757 ,n5104);
    nand g981(n354 ,n255 ,n332);
    xnor g982(n6530 ,n3451 ,n3458);
    not g983(n2449 ,n2448);
    nand g984(n1230 ,n1001 ,n886);
    nor g985(n2064 ,n20[1] ,n21[1]);
    dff g986(.RN(n1), .SN(1'b1), .CK(n0), .D(n1290), .Q(n11[12]));
    nand g987(n1719 ,n1577 ,n1675);
    dff g988(.RN(n1), .SN(1'b1), .CK(n0), .D(n1376), .Q(n23[1]));
    nand g989(n1316 ,n1074 ,n889);
    nand g990(n3359 ,n6578 ,n3358);
    xor g991(n6089 ,n6017 ,n6029);
    xnor g992(n2507 ,n2473 ,n2405);
    xnor g993(n5446 ,n5296 ,n5207);
    nand g994(n544 ,n536 ,n543);
    nor g995(n606 ,n23[0] ,n34[0]);
    nand g996(n4622 ,n20[4] ,n4363);
    nor g997(n6480 ,n6389 ,n6476);
    nand g998(n3852 ,n3647 ,n3801);
    or g999(n336 ,n185 ,n311);
    not g1000(n3493 ,n19[7]);
    xnor g1001(n2259 ,n2120 ,n2206);
    nand g1002(n1131 ,n20[6] ,n722);
    nor g1003(n263 ,n188 ,n227);
    nand g1004(n1305 ,n1062 ,n810);
    xnor g1005(n5524 ,n5312 ,n5068);
    xnor g1006(n2109 ,n2075 ,n2072);
    nor g1007(n2773 ,n2651 ,n2689);
    nor g1008(n2017 ,n1973 ,n1992);
    nor g1009(n5246 ,n5079 ,n5119);
    nand g1010(n4351 ,n4350 ,n4335);
    or g1011(n4764 ,n4494 ,n4572);
    xor g1012(n4934 ,n4557 ,n4495);
    dff g1013(.RN(n1), .SN(1'b1), .CK(n0), .D(n1305), .Q(n11[1]));
    not g1014(n4786 ,n4785);
    xnor g1015(n2271 ,n2109 ,n2209);
    not g1016(n2108 ,n2109);
    xnor g1017(n2393 ,n2325 ,n2274);
    nand g1018(n3818 ,n3566 ,n3711);
    nor g1019(n3018 ,n2901 ,n2988);
    nand g1020(n1284 ,n864 ,n1039);
    xor g1021(n6525 ,n6587 ,n6564);
    nor g1022(n3389 ,n6559 ,n6544);
    nor g1023(n6462 ,n6384 ,n6445);
    or g1024(n3225 ,n3178 ,n3197);
    nand g1025(n3809 ,n3621 ,n3714);
    nand g1026(n2463 ,n2280 ,n2432);
    xnor g1027(n4301 ,n4267 ,n4227);
    nand g1028(n2134 ,n6536 ,n2121);
    nand g1029(n3327 ,n6586 ,n41[13]);
    nand g1030(n3530 ,n3468 ,n3485);
    nand g1031(n3700 ,n3575 ,n3580);
    not g1032(n5407 ,n5380);
    dff g1033(.RN(n1), .SN(1'b1), .CK(n0), .D(n1313), .Q(n10[9]));
    nand g1034(n199 ,n165 ,n157);
    xnor g1035(n664 ,n35[15] ,n33[15]);
    nand g1036(n6384 ,n6311 ,n6350);
    nor g1037(n4021 ,n3935 ,n3969);
    not g1038(n313 ,n312);
    nand g1039(n1493 ,n796 ,n1490);
    or g1040(n4759 ,n4623 ,n4592);
    nand g1041(n4638 ,n4384 ,n20[3]);
    dff g1042(.RN(n1), .SN(1'b1), .CK(n0), .D(n1428), .Q(n19[6]));
    nand g1043(n627 ,n23[4] ,n34[4]);
    xor g1044(n4890 ,n4678 ,n4433);
    nand g1045(n5256 ,n5068 ,n5074);
    nand g1046(n4577 ,n21[0] ,n4373);
    nand g1047(n1415 ,n984 ,n1171);
    nand g1048(n5501 ,n5251 ,n5354);
    nand g1049(n4616 ,n4388 ,n20[1]);
    nand g1050(n1241 ,n1102 ,n750);
    nor g1051(n794 ,n17[0] ,n707);
    nand g1052(n1697 ,n1576 ,n1654);
    nor g1053(n5234 ,n5114 ,n5109);
    not g1054(n4521 ,n4520);
    xnor g1055(n2294 ,n2249 ,n2118);
    xor g1056(n4905 ,n4672 ,n4623);
    nand g1057(n6223 ,n25[1] ,n6226);
    xnor g1058(n5442 ,n5299 ,n5122);
    nand g1059(n6183 ,n6142 ,n6170);
    nand g1060(n1656 ,n1586 ,n1652);
    nand g1061(n3154 ,n38[0] ,n3136);
    nand g1062(n1433 ,n1189 ,n888);
    nand g1063(n5511 ,n5205 ,n5458);
    nand g1064(n3869 ,n3676 ,n3816);
    buf g1065(n13[14], n10[14]);
    or g1066(n5332 ,n5167 ,n5184);
    xnor g1067(n1880 ,n1749 ,n1805);
    nand g1068(n5586 ,n5318 ,n5475);
    xnor g1069(n5833 ,n5697 ,n5506);
    nand g1070(n1370 ,n819 ,n1119);
    nand g1071(n1862 ,n1701 ,n1820);
    nand g1072(n4869 ,n4624 ,n4455);
    dff g1073(.RN(n1), .SN(1'b1), .CK(n0), .D(n1259), .Q(n19[2]));
    nand g1074(n5317 ,n4877 ,n5162);
    nor g1075(n266 ,n248 ,n210);
    xnor g1076(n3451 ,n36[3] ,n19[3]);
    nand g1077(n3572 ,n3486 ,n19[7]);
    nand g1078(n3994 ,n3862 ,n3889);
    nand g1079(n1448 ,n1033 ,n1281);
    dff g1080(.RN(n1), .SN(1'b1), .CK(n0), .D(n1265), .Q(n1507));
    xnor g1081(n2414 ,n2378 ,n2262);
    or g1082(n5680 ,n5522 ,n5521);
    xnor g1083(n675 ,n35[7] ,n33[7]);
    nand g1084(n3417 ,n3387 ,n3416);
    nand g1085(n4612 ,n20[4] ,n4374);
    xnor g1086(n2983 ,n2913 ,n2732);
    xnor g1087(n5823 ,n5693 ,n5500);
    nand g1088(n5544 ,n5347 ,n5449);
    nand g1089(n4445 ,n4386 ,n20[5]);
    nor g1090(n2345 ,n2318 ,n2285);
    nand g1091(n3502 ,n3476 ,n19[5]);
    xnor g1092(n6607 ,n3411 ,n3419);
    nor g1093(n695 ,n620 ,n662);
    nor g1094(n3614 ,n3496 ,n3498);
    xnor g1095(n2870 ,n2801 ,n2671);
    xor g1096(n6609 ,n3405 ,n3400);
    nor g1097(n2518 ,n2504 ,n2494);
    xnor g1098(n5174 ,n4930 ,n4457);
    dff g1099(.RN(n1), .SN(1'b1), .CK(n0), .D(n1279), .Q(n1501));
    nand g1100(n1725 ,n1576 ,n1675);
    xnor g1101(n4064 ,n3953 ,n3854);
    xnor g1102(n1539 ,n91 ,n96);
    nand g1103(n181 ,n159 ,n150);
    nand g1104(n2048 ,n2034 ,n2047);
    not g1105(n3338 ,n3337);
    not g1106(n3683 ,n3682);
    or g1107(n4337 ,n4316 ,n4325);
    nor g1108(n121 ,n24[1] ,n24[0]);
    nand g1109(n5540 ,n5326 ,n5467);
    nand g1110(n904 ,n23[12] ,n715);
    nand g1111(n1692 ,n1580 ,n1654);
    nand g1112(n5046 ,n4559 ,n4802);
    not g1113(n4399 ,n4365);
    nand g1114(n6219 ,n6218 ,n6192);
    nand g1115(n6410 ,n6279 ,n6337);
    nand g1116(n1098 ,n1520 ,n716);
    xnor g1117(n5600 ,n5497 ,n5492);
    or g1118(n4719 ,n4641 ,n4600);
    nand g1119(n3080 ,n3062 ,n3079);
    nand g1120(n1016 ,n3[5] ,n713);
    not g1121(n156 ,n37[1]);
    nand g1122(n5951 ,n5737 ,n5888);
    nor g1123(n3178 ,n38[1] ,n3155);
    nor g1124(n2716 ,n2566 ,n2631);
    or g1125(n743 ,n717 ,n672);
    nand g1126(n5108 ,n4712 ,n5017);
    or g1127(n4772 ,n4621 ,n4422);
    xnor g1128(n5519 ,n5301 ,n5220);
    xnor g1129(n466 ,n424 ,n442);
    xnor g1130(n367 ,n307 ,n237);
    or g1131(n4748 ,n4585 ,n4608);
    nand g1132(n1712 ,n1586 ,n1677);
    xnor g1133(n4224 ,n4184 ,n4194);
    nand g1134(n1110 ,n1524 ,n716);
    nand g1135(n471 ,n457 ,n446);
    nand g1136(n4623 ,n21[3] ,n4373);
    nand g1137(n5012 ,n4687 ,n4833);
    nand g1138(n6123 ,n6077 ,n6101);
    nand g1139(n935 ,n28[7] ,n717);
    nand g1140(n1108 ,n1523 ,n716);
    xnor g1141(n5834 ,n5694 ,n5586);
    xnor g1142(n537 ,n522 ,n515);
    nand g1143(n4430 ,n4388 ,n20[4]);
    nor g1144(n2781 ,n2609 ,n2687);
    nor g1145(n770 ,n601 ,n555);
    nand g1146(n1242 ,n1106 ,n752);
    not g1147(n5520 ,n5519);
    xnor g1148(n1870 ,n1800 ,n1819);
    or g1149(n1499 ,n1495 ,n1498);
    dff g1150(.RN(n1), .SN(1'b1), .CK(n0), .D(n1451), .Q(n34[2]));
    nor g1151(n2042 ,n2012 ,n2041);
    nor g1152(n2564 ,n2519 ,n2563);
    nor g1153(n3802 ,n3572 ,n3737);
    xnor g1154(n2296 ,n2226 ,n2120);
    nand g1155(n5255 ,n5110 ,n5135);
    nor g1156(n5447 ,n5226 ,n5346);
    nand g1157(n3416 ,n3400 ,n3406);
    xnor g1158(n4186 ,n4095 ,n4055);
    not g1159(n5800 ,n5799);
    xnor g1160(n690 ,n23[3] ,n34[3]);
    nand g1161(n4294 ,n4245 ,n4270);
    nand g1162(n6352 ,n6588 ,n6247);
    xnor g1163(n2073 ,n21[6] ,n21[5]);
    nand g1164(n5366 ,n5150 ,n5244);
    xnor g1165(n3887 ,n3776 ,n3503);
    nor g1166(n2941 ,n2835 ,n2905);
    nand g1167(n2216 ,n6539 ,n2178);
    buf g1168(n36[4] ,n1512);
    nor g1169(n1556 ,n123 ,n121);
    nand g1170(n2537 ,n2522 ,n2533);
    nor g1171(n580 ,n16[8] ,n23[8]);
    nand g1172(n1743 ,n1661 ,n1708);
    nand g1173(n1359 ,n910 ,n1110);
    nand g1174(n5069 ,n4705 ,n4988);
    nand g1175(n1912 ,n1855 ,n1898);
    not g1176(n3280 ,n36[1]);
    nand g1177(n4435 ,n20[6] ,n4373);
    nand g1178(n5095 ,n4724 ,n5039);
    xnor g1179(n1993 ,n1946 ,n1964);
    nand g1180(n1911 ,n1848 ,n1896);
    nand g1181(n4482 ,n4380 ,n20[5]);
    xor g1182(n40[14] ,n6597 ,n38[15]);
    nand g1183(n4634 ,n20[6] ,n4374);
    nor g1184(n5924 ,n5876 ,n5868);
    xor g1185(n6517 ,n6579 ,n6556);
    dff g1186(.RN(n1), .SN(1'b1), .CK(n0), .D(n1472), .Q(n27[6]));
    dff g1187(.RN(n1), .SN(1'b1), .CK(n0), .D(n1466), .Q(n28[6]));
    xnor g1188(n5771 ,n5648 ,n5576);
    not g1189(n5119 ,n5044);
    nand g1190(n2248 ,n2164 ,n2197);
    not g1191(n2231 ,n2232);
    nand g1192(n972 ,n21[0] ,n714);
    not g1193(n6252 ,n6253);
    nor g1194(n3440 ,n3410 ,n3439);
    nand g1195(n1609 ,n19[4] ,n1595);
    nand g1196(n4702 ,n21[2] ,n4369);
    nand g1197(n6356 ,n6503 ,n6249);
    nand g1198(n1660 ,n1577 ,n1652);
    nand g1199(n5005 ,n4657 ,n4832);
    nand g1200(n3851 ,n3663 ,n3814);
    nand g1201(n5506 ,n5262 ,n5361);
    dff g1202(.RN(n1), .SN(1'b1), .CK(n0), .D(n1471), .Q(n27[8]));
    nand g1203(n5904 ,n5752 ,n5843);
    nand g1204(n1154 ,n23[11] ,n716);
    or g1205(n2944 ,n2827 ,n2926);
    nand g1206(n5017 ,n4693 ,n4836);
    nor g1207(n2063 ,n20[7] ,n21[7]);
    nand g1208(n5107 ,n4716 ,n5024);
    or g1209(n4723 ,n4624 ,n4455);
    not g1210(n3736 ,n3716);
    not g1211(n145 ,n37[6]);
    nand g1212(n1366 ,n817 ,n1051);
    nand g1213(n959 ,n27[12] ,n715);
    nand g1214(n1964 ,n1788 ,n1941);
    xnor g1215(n677 ,n35[0] ,n33[0]);
    nor g1216(n6258 ,n6232 ,n6252);
    xnor g1217(n309 ,n199 ,n197);
    not g1218(n2152 ,n2151);
    not g1219(n3577 ,n3576);
    nor g1220(n2332 ,n2263 ,n2312);
    nand g1221(n2213 ,n6536 ,n2178);
    dff g1222(.RN(n1), .SN(1'b1), .CK(n0), .D(n1393), .Q(n27[14]));
    nand g1223(n1332 ,n896 ,n1086);
    xnor g1224(n3953 ,n3844 ,n3684);
    nand g1225(n1695 ,n1588 ,n1654);
    nand g1226(n3386 ,n3324 ,n3385);
    nor g1227(n582 ,n34[9] ,n34[10]);
    xor g1228(n1796 ,n1757 ,n1701);
    nand g1229(n1413 ,n658 ,n786);
    nand g1230(n4316 ,n4292 ,n4304);
    nand g1231(n4451 ,n4382 ,n20[1]);
    xnor g1232(n5633 ,n5437 ,n5158);
    nand g1233(n1662 ,n1584 ,n1651);
    nand g1234(n6436 ,n6297 ,n6362);
    dff g1235(.RN(n1), .SN(1'b1), .CK(n0), .D(n1424), .Q(n26[3]));
    not g1236(n2917 ,n2916);
    nor g1237(n616 ,n16[4] ,n23[4]);
    or g1238(n3184 ,n3166 ,n3183);
    xnor g1239(n5974 ,n5860 ,n5885);
    not g1240(n2505 ,n2504);
    nor g1241(n2536 ,n2497 ,n2534);
    xnor g1242(n2288 ,n2225 ,n2120);
    xnor g1243(n2953 ,n2866 ,n2898);
    nand g1244(n6361 ,n6586 ,n6247);
    nand g1245(n4808 ,n4437 ,n4596);
    dff g1246(.RN(n1), .SN(1'b1), .CK(n0), .D(n1255), .Q(n25[0]));
    nand g1247(n5035 ,n4522 ,n4856);
    xor g1248(n3955 ,n3843 ,n3874);
    nand g1249(n3583 ,n3462 ,n3480);
    nand g1250(n2239 ,n2130 ,n2215);
    nand g1251(n2962 ,n2914 ,n2922);
    or g1252(n4743 ,n4628 ,n4635);
    nand g1253(n5001 ,n4694 ,n4803);
    nor g1254(n2011 ,n1958 ,n2007);
    nand g1255(n4875 ,n4490 ,n4454);
    nand g1256(n6338 ,n6582 ,n6247);
    xnor g1257(n5968 ,n5863 ,n5830);
    nand g1258(n1747 ,n1671 ,n1736);
    nand g1259(n2129 ,n6533 ,n2121);
    or g1260(n5927 ,n5834 ,n5870);
    xnor g1261(n5179 ,n4886 ,n4622);
    not g1262(n2924 ,n2923);
    nand g1263(n1492 ,n661 ,n1490);
    nand g1264(n1173 ,n29[7] ,n724);
    xor g1265(n6608 ,n3408 ,n3417);
    xnor g1266(n5820 ,n5725 ,n5598);
    not g1267(n3271 ,n3270);
    nor g1268(n2459 ,n2360 ,n2420);
    nand g1269(n4532 ,n20[1] ,n4367);
    xnor g1270(n1968 ,n1929 ,n1867);
    xnor g1271(n4342 ,n4315 ,n4326);
    nor g1272(n5663 ,n5576 ,n5579);
    dff g1273(.RN(n1), .SN(1'b1), .CK(n0), .D(n1458), .Q(n31[0]));
    not g1274(n2483 ,n2482);
    nand g1275(n4568 ,n21[4] ,n4365);
    dff g1276(.RN(n1), .SN(1'b1), .CK(n0), .D(n1312), .Q(n10[10]));
    xnor g1277(n666 ,n19[7] ,n27[7]);
    dff g1278(.RN(n1), .SN(1'b1), .CK(n0), .D(n1419), .Q(n26[6]));
    xnor g1279(n6108 ,n6027 ,n6080);
    nor g1280(n2751 ,n2612 ,n2688);
    xnor g1281(n6546 ,n3333 ,n3380);
    xor g1282(n3743 ,n3639 ,n3518);
    not g1283(n1573 ,n37[1]);
    nand g1284(n3806 ,n3630 ,n3730);
    nand g1285(n3165 ,n3109 ,n3147);
    not g1286(n154 ,n37[3]);
    xnor g1287(n6176 ,n6122 ,n6146);
    xnor g1288(n2866 ,n2706 ,n2753);
    nand g1289(n2845 ,n2781 ,n2755);
    nand g1290(n6444 ,n6244 ,n6262);
    or g1291(n3012 ,n2983 ,n2982);
    nand g1292(n5266 ,n5121 ,n5120);
    xnor g1293(n2869 ,n2745 ,n2660);
    nand g1294(n4656 ,n21[1] ,n4371);
    not g1295(n4559 ,n4558);
    nand g1296(n6011 ,n5931 ,n5971);
    nor g1297(n1533 ,n177 ,n175);
    nand g1298(n3044 ,n3019 ,n3023);
    nand g1299(n6288 ,n6560 ,n6251);
    xnor g1300(n5208 ,n4910 ,n4572);
    nand g1301(n847 ,n19[0] ,n714);
    nor g1302(n6483 ,n6406 ,n6474);
    xnor g1303(n4142 ,n4044 ,n4078);
    nand g1304(n653 ,n23[0] ,n34[0]);
    xnor g1305(n4095 ,n4026 ,n4047);
    not g1306(n3480 ,n3479);
    nor g1307(n2637 ,n2566 ,n2585);
    nand g1308(n548 ,n527 ,n547);
    nand g1309(n1475 ,n927 ,n1214);
    nand g1310(n927 ,n29[7] ,n721);
    not g1311(n5621 ,n5620);
    xnor g1312(n4895 ,n4631 ,n4439);
    nand g1313(n1899 ,n1785 ,n1856);
    nand g1314(n5808 ,n5675 ,n5749);
    nand g1315(n5150 ,n4774 ,n5032);
    xnor g1316(n6095 ,n6024 ,n6002);
    not g1317(n135 ,n134);
    or g1318(n252 ,n186 ,n216);
    xnor g1319(n1637 ,n1613 ,n1601);
    xnor g1320(n2008 ,n1975 ,n1912);
    nand g1321(n457 ,n398 ,n437);
    nand g1322(n635 ,n33[3] ,n35[3]);
    nand g1323(n191 ,n172 ,n146);
    xnor g1324(n538 ,n523 ,n517);
    dff g1325(.RN(n1), .SN(1'b1), .CK(n0), .D(n1371), .Q(n23[3]));
    xnor g1326(n3769 ,n3581 ,n3533);
    xnor g1327(n6547 ,n3340 ,n3382);
    nor g1328(n2068 ,n20[3] ,n21[3]);
    xnor g1329(n1535 ,n85 ,n104);
    xnor g1330(n5640 ,n5436 ,n5114);
    xnor g1331(n2263 ,n2108 ,n2205);
    nor g1332(n4523 ,n4415 ,n4401);
    nand g1333(n1426 ,n991 ,n1181);
    xor g1334(n6512 ,n6551 ,n6574);
    dff g1335(.RN(n1), .SN(1'b1), .CK(n0), .D(n1256), .Q(n16[6]));
    nor g1336(n2679 ,n2565 ,n2627);
    nor g1337(n1959 ,n1908 ,n1931);
    not g1338(n3472 ,n3471);
    nand g1339(n4293 ,n4218 ,n4271);
    nand g1340(n2234 ,n2132 ,n2213);
    not g1341(n53 ,n52);
    nor g1342(n609 ,n21[6] ,n30[6]);
    nand g1343(n1247 ,n1136 ,n781);
    nand g1344(n5109 ,n4750 ,n5015);
    nor g1345(n2885 ,n2771 ,n2820);
    nand g1346(n848 ,n1507 ,n714);
    xnor g1347(n6032 ,n5958 ,n5975);
    xnor g1348(n1653 ,n1617 ,n1637);
    xnor g1349(n5645 ,n5446 ,n5208);
    nand g1350(n2205 ,n2090 ,n2160);
    nand g1351(n3528 ,n3486 ,n19[1]);
    nand g1352(n6336 ,n6574 ,n6247);
    nand g1353(n1941 ,n1787 ,n1918);
    xnor g1354(n3179 ,n38[8] ,n3130);
    xnor g1355(n2038 ,n2024 ,n2018);
    nor g1356(n4135 ,n3959 ,n4075);
    not g1357(n4027 ,n4026);
    nand g1358(n5940 ,n5834 ,n5870);
    xnor g1359(n447 ,n394 ,n368);
    nand g1360(n1041 ,n1541 ,n557);
    buf g1361(n36[1] ,n1509);
    nand g1362(n215 ,n167 ,n152);
    nand g1363(n4133 ,n4048 ,n4053);
    xnor g1364(n4912 ,n4437 ,n4596);
    nand g1365(n3376 ,n3326 ,n3375);
    not g1366(n1589 ,n36[3]);
    or g1367(n2066 ,n20[4] ,n20[3]);
    nand g1368(n4467 ,n21[2] ,n4384);
    or g1369(n3664 ,n3509 ,n3534);
    nor g1370(n3613 ,n3496 ,n3494);
    buf g1371(n36[2] ,n1510);
    nand g1372(n4284 ,n4229 ,n4269);
    not g1373(n6026 ,n6025);
    not g1374(n5907 ,n5906);
    not g1375(n2853 ,n2845);
    xnor g1376(n3915 ,n3779 ,n3682);
    nand g1377(n491 ,n447 ,n463);
    nand g1378(n3596 ,n3480 ,n19[6]);
    xnor g1379(n3051 ,n3022 ,n2996);
    dff g1380(.RN(n1), .SN(1'b1), .CK(n0), .D(n1328), .Q(n34[8]));
    nand g1381(n5151 ,n4758 ,n5038);
    xnor g1382(n5522 ,n5314 ,n5102);
    xnor g1383(n4209 ,n4139 ,n4061);
    nor g1384(n107 ,n24[3] ,n24[2]);
    nand g1385(n3367 ,n41[6] ,n3366);
    xnor g1386(n5599 ,n5494 ,n5499);
    not g1387(n6006 ,n6005);
    xnor g1388(n4963 ,n4555 ,n4539);
    nand g1389(n4686 ,n21[5] ,n4388);
    nand g1390(n5676 ,n5580 ,n5572);
    nand g1391(n3240 ,n3196 ,n3239);
    xor g1392(n4917 ,n4509 ,n4448);
    nand g1393(n976 ,n27[4] ,n715);
    nand g1394(n5014 ,n4529 ,n4835);
    nand g1395(n2281 ,n2120 ,n2241);
    nand g1396(n1722 ,n1622 ,n1683);
    nand g1397(n4655 ,n21[0] ,n4374);
    nand g1398(n5018 ,n4517 ,n4838);
    nor g1399(n619 ,n22[3] ,n26[3]);
    nand g1400(n3538 ,n3462 ,n3476);
    nand g1401(n5064 ,n4789 ,n4958);
    nand g1402(n920 ,n30[4] ,n723);
    nand g1403(n182 ,n167 ,n148);
    nand g1404(n4983 ,n4546 ,n4868);
    nand g1405(n3076 ,n3053 ,n3075);
    nor g1406(n2988 ,n2927 ,n2954);
    nand g1407(n4601 ,n20[5] ,n4369);
    not g1408(n1193 ,n1135);
    xnor g1409(n307 ,n190 ,n181);
    nor g1410(n6251 ,n6227 ,n6228);
    nand g1411(n1661 ,n1580 ,n1652);
    nand g1412(n6107 ,n6039 ,n6074);
    nand g1413(n3251 ,n3208 ,n3250);
    nand g1414(n829 ,n17[1] ,n721);
    nand g1415(n4486 ,n4384 ,n20[5]);
    not g1416(n3489 ,n36[4]);
    dff g1417(.RN(n1), .SN(1'b1), .CK(n0), .D(n1318), .Q(n10[5]));
    nor g1418(n1960 ,n1842 ,n1932);
    nand g1419(n459 ,n414 ,n434);
    or g1420(n772 ,n720 ,n674);
    xnor g1421(n5648 ,n5441 ,n5087);
    xnor g1422(n6551 ,n3681 ,n4017);
    nand g1423(n6218 ,n6190 ,n6217);
    not g1424(n169 ,n168);
    or g1425(n3672 ,n3508 ,n3507);
    xnor g1426(n4050 ,n4001 ,n3892);
    nand g1427(n2172 ,n6541 ,n2122);
    xnor g1428(n2367 ,n2286 ,n2317);
    nand g1429(n2282 ,n2119 ,n2240);
    not g1430(n3780 ,n3779);
    nor g1431(n4202 ,n4196 ,n4183);
    nand g1432(n1156 ,n23[10] ,n716);
    or g1433(n886 ,n710 ,n670);
    nand g1434(n4479 ,n21[4] ,n4373);
    nand g1435(n4018 ,n3902 ,n3974);
    nor g1436(n4976 ,n4612 ,n4786);
    xnor g1437(n1804 ,n1648 ,n1740);
    nand g1438(n1028 ,n3[1] ,n713);
    nor g1439(n344 ,n263 ,n333);
    nand g1440(n5143 ,n4710 ,n5010);
    nand g1441(n4192 ,n4131 ,n4170);
    xnor g1442(n6166 ,n6126 ,n6131);
    nor g1443(n2743 ,n2662 ,n2729);
    xnor g1444(n1634 ,n1591 ,n1607);
    nand g1445(n3998 ,n3877 ,n3918);
    xnor g1446(n2894 ,n2795 ,n2850);
    nand g1447(n923 ,n30[2] ,n723);
    not g1448(n5778 ,n5777);
    nand g1449(n1312 ,n1070 ,n952);
    nor g1450(n4510 ,n4417 ,n4415);
    xnor g1451(n4116 ,n4011 ,n4029);
    nand g1452(n4991 ,n4553 ,n4822);
    nand g1453(n5019 ,n4670 ,n4809);
    not g1454(n4792 ,n4791);
    xnor g1455(n6186 ,n6155 ,n6166);
    xnor g1456(n4222 ,n4197 ,n4154);
    xnor g1457(n485 ,n426 ,n449);
    nor g1458(n3351 ,n3348 ,n3350);
    not g1459(n3484 ,n3483);
    nand g1460(n1453 ,n1104 ,n1351);
    nand g1461(n4040 ,n3853 ,n3962);
    not g1462(n4956 ,n4955);
    not g1463(n2268 ,n2267);
    nand g1464(n5674 ,n5587 ,n5515);
    nor g1465(n589 ,n31[4] ,n35[4]);
    xnor g1466(n687 ,n35[4] ,n33[4]);
    not g1467(n205 ,n204);
    not g1468(n3356 ,n3355);
    or g1469(n5451 ,n5191 ,n5350);
    xnor g1470(n6491 ,n3214 ,n3239);
    not g1471(n4407 ,n20[0]);
    or g1472(n5467 ,n5228 ,n5409);
    not g1473(n4677 ,n4676);
    nor g1474(n1839 ,n1780 ,n1825);
    nand g1475(n6303 ,n40[0] ,n6250);
    nand g1476(n3238 ,n3184 ,n3237);
    nand g1477(n1140 ,n22[2] ,n720);
    xnor g1478(n6493 ,n3220 ,n3243);
    xnor g1479(n3413 ,n39[5] ,n6554);
    nand g1480(n6351 ,n6492 ,n6253);
    xnor g1481(n2371 ,n2119 ,n2297);
    xnor g1482(n5866 ,n5786 ,n5609);
    nand g1483(n3924 ,n3876 ,n3834);
    nor g1484(n568 ,n26[5] ,n26[6]);
    xnor g1485(n4287 ,n4250 ,n4211);
    nand g1486(n2224 ,n2144 ,n2182);
    xnor g1487(n362 ,n298 ,n182);
    nand g1488(n1627 ,n1607 ,n1603);
    not g1489(n3341 ,n3340);
    nand g1490(n1737 ,n1588 ,n1677);
    xnor g1491(n393 ,n308 ,n345);
    xnor g1492(n4016 ,n3895 ,n3896);
    nand g1493(n4480 ,n4382 ,n20[0]);
    nand g1494(n6280 ,n6559 ,n6251);
    nand g1495(n2740 ,n6527 ,n2618);
    nand g1496(n2050 ,n2037 ,n2049);
    nand g1497(n1696 ,n1588 ,n1652);
    nand g1498(n5893 ,n5781 ,n5835);
    nand g1499(n6182 ,n6155 ,n6166);
    nand g1500(n1841 ,n1645 ,n1817);
    nand g1501(n940 ,n28[3] ,n717);
    nand g1502(n2186 ,n6535 ,n2150);
    nand g1503(n1202 ,n828 ,n792);
    nand g1504(n6329 ,n38[0] ,n6246);
    nand g1505(n1049 ,n31[7] ,n720);
    xnor g1506(n3781 ,n3622 ,n3610);
    nor g1507(n3388 ,n6556 ,n39[7]);
    nand g1508(n1043 ,n2[4] ,n713);
    xnor g1509(n676 ,n23[7] ,n16[7]);
    xnor g1510(n5183 ,n4890 ,n4565);
    xnor g1511(n5224 ,n4891 ,n4549);
    nor g1512(n3794 ,n3526 ,n3681);
    nand g1513(n188 ,n167 ,n155);
    nand g1514(n6075 ,n5990 ,n6036);
    xnor g1515(n2078 ,n21[2] ,n20[2]);
    nand g1516(n1170 ,n5[4] ,n557);
    xnor g1517(n5879 ,n5763 ,n5612);
    nand g1518(n5088 ,n4776 ,n5012);
    dff g1519(.RN(n1), .SN(1'b1), .CK(n0), .D(n1250), .Q(n22[2]));
    xor g1520(n4950 ,n4659 ,n4563);
    nor g1521(n3436 ,n3402 ,n3435);
    nand g1522(n5084 ,n4714 ,n5007);
    nand g1523(n840 ,n19[4] ,n556);
    nand g1524(n35[11] ,n6462 ,n6468);
    nand g1525(n2220 ,n6540 ,n2149);
    nor g1526(n1840 ,n1645 ,n1817);
    dff g1527(.RN(n1), .SN(1'b1), .CK(n0), .D(n1331), .Q(n10[0]));
    xnor g1528(n4229 ,n4175 ,n4116);
    nor g1529(n5706 ,n5638 ,n5649);
    not g1530(n123 ,n122);
    not g1531(n3459 ,n37[7]);
    nand g1532(n1665 ,n1584 ,n1649);
    nand g1533(n2936 ,n2849 ,n2906);
    xnor g1534(n519 ,n506 ,n466);
    nor g1535(n6236 ,n41[6] ,n6594);
    nor g1536(n2007 ,n1962 ,n1983);
    xnor g1537(n5767 ,n5627 ,n5574);
    nand g1538(n6427 ,n6360 ,n6359);
    not g1539(n1618 ,n19[0]);
    nand g1540(n1856 ,n1802 ,n1801);
    nor g1541(n2402 ,n2345 ,n2383);
    not g1542(n4372 ,n37[3]);
    nor g1543(n4512 ,n4406 ,n4402);
    nor g1544(n2898 ,n2814 ,n2885);
    nand g1545(n926 ,n30[0] ,n723);
    nor g1546(n2635 ,n2566 ,n2594);
    or g1547(n3103 ,n38[11] ,n6584);
    nand g1548(n2253 ,n2170 ,n2194);
    not g1549(n315 ,n314);
    nand g1550(n705 ,n596 ,n599);
    nand g1551(n3715 ,n3587 ,n3592);
    not g1552(n3574 ,n3573);
    nand g1553(n4988 ,n4703 ,n4811);
    nand g1554(n2196 ,n6539 ,n2148);
    xnor g1555(n1877 ,n1776 ,n1821);
    nor g1556(n2768 ,n2615 ,n2717);
    not g1557(n176 ,n148);
    nand g1558(n4500 ,n4389 ,n20[7]);
    nor g1559(n2357 ,n2236 ,n2315);
    nand g1560(n3527 ,n3476 ,n19[3]);
    xnor g1561(n464 ,n422 ,n431);
    nand g1562(n873 ,n1510 ,n714);
    xnor g1563(n5970 ,n5859 ,n5812);
    buf g1564(n14[11], n11[11]);
    not g1565(n1195 ,n1166);
    nand g1566(n2257 ,n2174 ,n2196);
    nand g1567(n1425 ,n801 ,n1182);
    xnor g1568(n2632 ,n40[13] ,n6524);
    nand g1569(n5792 ,n5754 ,n5719);
    xnor g1570(n5314 ,n5108 ,n5085);
    or g1571(n4704 ,n4442 ,n4459);
    dff g1572(.RN(n1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n33[8]));
    nand g1573(n1017 ,n12[8] ,n555);
    nand g1574(n865 ,n33[14] ,n554);
    or g1575(n5336 ,n5221 ,n5246);
    or g1576(n5749 ,n5585 ,n5662);
    nand g1577(n2157 ,n6539 ,n2127);
    nand g1578(n2093 ,n6535 ,n2085);
    nor g1579(n4099 ,n4046 ,n4077);
    nor g1580(n597 ,n22[0] ,n26[0]);
    xnor g1581(n5688 ,n5445 ,n5165);
    nand g1582(n2169 ,n6536 ,n2126);
    or g1583(n2056 ,n2055 ,n1998);
    nand g1584(n6314 ,n6549 ,n6248);
    nand g1585(n3723 ,n3584 ,n3547);
    nand g1586(n2429 ,n2391 ,n2396);
    nand g1587(n4159 ,n4088 ,n4127);
    not g1588(n369 ,n368);
    xnor g1589(n3946 ,n3847 ,n3853);
    nand g1590(n5149 ,n4765 ,n5041);
    or g1591(n4236 ,n4192 ,n4206);
    nor g1592(n4648 ,n4393 ,n4416);
    nand g1593(n3531 ,n3484 ,n19[2]);
    nand g1594(n1292 ,n869 ,n1045);
    xnor g1595(n4062 ,n3954 ,n3849);
    nand g1596(n1897 ,n1791 ,n1846);
    not g1597(n3454 ,n3453);
    xnor g1598(n672 ,n19[0] ,n27[0]);
    nor g1599(n5324 ,n5193 ,n5192);
    nor g1600(n1823 ,n1783 ,n1795);
    xnor g1601(n303 ,n180 ,n222);
    nand g1602(n907 ,n1544 ,n712);
    nor g1603(n5841 ,n5617 ,n5801);
    nand g1604(n808 ,n35[3] ,n712);
    not g1605(n558 ,n18[0]);
    or g1606(n4734 ,n4498 ,n4500);
    xnor g1607(n5160 ,n4934 ,n4639);
    nand g1608(n6044 ,n5950 ,n6005);
    not g1609(n5403 ,n5402);
    xnor g1610(n4961 ,n4526 ,n4666);
    xor g1611(n2116 ,n2098 ,n2087);
    nor g1612(n5656 ,n5550 ,n5537);
    xnor g1613(n6573 ,n1636 ,n1653);
    not g1614(n5123 ,n5122);
    dff g1615(.RN(n1), .SN(1'b1), .CK(n0), .D(n1432), .Q(n25[1]));
    nand g1616(n4340 ,n4319 ,n4324);
    xnor g1617(n403 ,n303 ,n354);
    nor g1618(n260 ,n232 ,n187);
    nand g1619(n2147 ,n6536 ,n2123);
    xnor g1620(n427 ,n386 ,n371);
    nand g1621(n348 ,n272 ,n315);
    nor g1622(n2729 ,n2567 ,n2633);
    nand g1623(n1132 ,n22[6] ,n720);
    dff g1624(.RN(n1), .SN(1'b1), .CK(n0), .D(n1436), .Q(n29[4]));
    nand g1625(n917 ,n17[7] ,n721);
    xnor g1626(n41[12] ,n6204 ,n6215);
    nand g1627(n3326 ,n6582 ,n6570);
    nand g1628(n2228 ,n2142 ,n2179);
    nor g1629(n2817 ,n2664 ,n2758);
    nand g1630(n1221 ,n940 ,n747);
    nand g1631(n4626 ,n4376 ,n20[1]);
    nor g1632(n2381 ,n2297 ,n2341);
    xnor g1633(n3760 ,n3584 ,n3547);
    nand g1634(n3612 ,n3474 ,n3478);
    not g1635(n6096 ,n6095);
    nand g1636(n809 ,n35[2] ,n712);
    nand g1637(n5050 ,n4671 ,n4844);
    nand g1638(n5111 ,n4736 ,n5018);
    not g1639(n3621 ,n3620);
    nor g1640(n1889 ,n1835 ,n1807);
    nor g1641(n2711 ,n2568 ,n2630);
    nand g1642(n3797 ,n3617 ,n3720);
    xnor g1643(n3216 ,n3165 ,n3180);
    dff g1644(.RN(n1), .SN(1'b1), .CK(n0), .D(n1232), .Q(n12[7]));
    nand g1645(n3847 ,n3654 ,n3796);
    nand g1646(n1726 ,n1576 ,n1676);
    nand g1647(n4442 ,n4376 ,n20[7]);
    nand g1648(n183 ,n165 ,n155);
    nor g1649(n2541 ,n2513 ,n2529);
    or g1650(n2577 ,n40[2] ,n6513);
    nor g1651(n2738 ,n2567 ,n2617);
    nand g1652(n5944 ,n5753 ,n5895);
    dff g1653(.RN(n1), .SN(1'b1), .CK(n0), .D(n1378), .Q(n23[0]));
    nand g1654(n5572 ,n5332 ,n5470);
    not g1655(n4395 ,n21[4]);
    dff g1656(.RN(n1), .SN(1'b1), .CK(n0), .D(n1268), .Q(n1506));
    xnor g1657(n4115 ,n4015 ,n3912);
    nand g1658(n1357 ,n1111 ,n909);
    nand g1659(n5395 ,n5182 ,n5179);
    xnor g1660(n5960 ,n5875 ,n5802);
    xnor g1661(n5201 ,n4972 ,n4431);
    nand g1662(n1186 ,n8[2] ,n713);
    nand g1663(n1412 ,n978 ,n1169);
    nand g1664(n1480 ,n830 ,n1246);
    not g1665(n5525 ,n5524);
    nand g1666(n3140 ,n6558 ,n3093);
    or g1667(n4765 ,n4423 ,n4458);
    nand g1668(n6202 ,n6188 ,n6194);
    nand g1669(n6192 ,n6165 ,n6183);
    nor g1670(n2715 ,n2565 ,n2631);
    nand g1671(n6284 ,n40[9] ,n6250);
    nand g1672(n6271 ,n41[7] ,n6254);
    nor g1673(n5721 ,n5608 ,n5634);
    nand g1674(n3721 ,n3541 ,n3545);
    nand g1675(n5526 ,n5329 ,n5469);
    nor g1676(n1983 ,n1961 ,n1963);
    xnor g1677(n4226 ,n4173 ,n4201);
    xnor g1678(n1531 ,n358 ,n266);
    nand g1679(n4617 ,n20[4] ,n4371);
    or g1680(n3188 ,n3162 ,n3175);
    nand g1681(n214 ,n169 ,n148);
    not g1682(n5164 ,n5163);
    nand g1683(n862 ,n33[15] ,n712);
    xnor g1684(n359 ,n297 ,n316);
    nand g1685(n452 ,n409 ,n443);
    nand g1686(n286 ,n220 ,n221);
    xnor g1687(n6542 ,n6569 ,n3372);
    nand g1688(n5049 ,n4512 ,n4874);
    xor g1689(n2121 ,n2107 ,n2111);
    nand g1690(n236 ,n169 ,n153);
    nand g1691(n515 ,n488 ,n503);
    xnor g1692(n1872 ,n1804 ,n1803);
    nand g1693(n5742 ,n5584 ,n5652);
    nand g1694(n3456 ,n3448 ,n3455);
    nor g1695(n4554 ,n4408 ,n4413);
    nand g1696(n1745 ,n1663 ,n1711);
    nand g1697(n1482 ,n968 ,n1208);
    nand g1698(n3145 ,n6562 ,n3092);
    nor g1699(n2958 ,n2810 ,n2931);
    nand g1700(n6390 ,n6302 ,n6352);
    nand g1701(n5298 ,n4771 ,n5103);
    nand g1702(n504 ,n490 ,n494);
    nand g1703(n1622 ,n1580 ,n1612);
    not g1704(n365 ,n364);
    xnor g1705(n5176 ,n4894 ,n4644);
    or g1706(n3307 ,n3302 ,n3306);
    nor g1707(n5450 ,n5217 ,n5323);
    not g1708(n3295 ,n3294);
    xnor g1709(n6165 ,n6125 ,n6123);
    xnor g1710(n3782 ,n3570 ,n3643);
    nand g1711(n1368 ,n634 ,n756);
    xnor g1712(n5766 ,n5633 ,n5534);
    nand g1713(n3928 ,n3842 ,n3859);
    nand g1714(n4979 ,n4583 ,n4783);
    nand g1715(n1174 ,n5[1] ,n713);
    nor g1716(n1939 ,n1847 ,n1906);
    not g1717(n2752 ,n2751);
    xor g1718(n40[7] ,n6604 ,n38[8]);
    not g1719(n167 ,n166);
    nor g1720(n4508 ,n4404 ,n4396);
    not g1721(n4613 ,n4612);
    nand g1722(n5897 ,n5824 ,n5829);
    nand g1723(n1162 ,n6[1] ,n713);
    dff g1724(.RN(n1), .SN(1'b1), .CK(n0), .D(n1457), .Q(n31[1]));
    xnor g1725(n363 ,n319 ,n228);
    not g1726(n147 ,n37[4]);
    nand g1727(n4493 ,n21[5] ,n4373);
    dff g1728(.RN(n1), .SN(1'b1), .CK(n0), .D(n1360), .Q(n32[2]));
    xnor g1729(n698 ,n26[2] ,n22[2]);
    nor g1730(n4101 ,n3970 ,n4065);
    xnor g1731(n5217 ,n4882 ,n4499);
    nand g1732(n4641 ,n21[0] ,n4376);
    nand g1733(n1472 ,n971 ,n1407);
    nand g1734(n5895 ,n5779 ,n5830);
    nand g1735(n1339 ,n962 ,n1160);
    nand g1736(n2412 ,n2358 ,n2386);
    nand g1737(n501 ,n475 ,n479);
    nand g1738(n5295 ,n4742 ,n5105);
    nor g1739(n3420 ,n3411 ,n3419);
    nand g1740(n4081 ,n3963 ,n4041);
    xnor g1741(n3071 ,n3037 ,n3032);
    xnor g1742(n1197 ,n710 ,n32[0]);
    xnor g1743(n6005 ,n5913 ,n5826);
    nand g1744(n4123 ,n4082 ,n4058);
    nand g1745(n5584 ,n5327 ,n5489);
    nand g1746(n3593 ,n3464 ,n3482);
    nand g1747(n807 ,n35[4] ,n712);
    nor g1748(n5297 ,n4976 ,n5058);
    nor g1749(n602 ,n22[6] ,n26[6]);
    nand g1750(n1730 ,n1629 ,n1684);
    xor g1751(n3746 ,n3553 ,n3603);
    or g1752(n5337 ,n5198 ,n5156);
    nand g1753(n229 ,n170 ,n155);
    not g1754(n2828 ,n2823);
    xnor g1755(n4009 ,n3937 ,n3938);
    nor g1756(n1948 ,n1885 ,n1926);
    nor g1757(n2704 ,n2567 ,n2630);
    nand g1758(n4851 ,n4577 ,n4449);
    xnor g1759(n371 ,n300 ,n244);
    nand g1760(n247 ,n167 ,n157);
    nor g1761(n1906 ,n1866 ,n1891);
    not g1762(n2342 ,n2336);
    nand g1763(n6441 ,n6305 ,n6375);
    nor g1764(n1910 ,n1837 ,n1889);
    xnor g1765(n2300 ,n2118 ,n2238);
    nand g1766(n528 ,n513 ,n511);
    nor g1767(n736 ,n702 ,n701);
    nand g1768(n5753 ,n5565 ,n5665);
    nand g1769(n3510 ,n3481 ,n19[2]);
    xnor g1770(n4955 ,n4556 ,n4545);
    nand g1771(n6369 ,n38[4] ,n6246);
    xnor g1772(n1879 ,n1780 ,n1810);
    not g1773(n3481 ,n3489);
    nor g1774(n2665 ,n2568 ,n2586);
    xnor g1775(n5417 ,n5184 ,n5167);
    nand g1776(n5978 ,n5910 ,n5920);
    xnor g1777(n5956 ,n5877 ,n5831);
    nand g1778(n4565 ,n20[6] ,n4363);
    nand g1779(n4169 ,n4045 ,n4124);
    buf g1780(n13[8], n10[8]);
    xnor g1781(n5444 ,n5293 ,n5138);
    nand g1782(n3537 ,n3485 ,n19[2]);
    xor g1783(n4906 ,n4674 ,n4456);
    xnor g1784(n2863 ,n2782 ,n2667);
    nand g1785(n2331 ,n2317 ,n2286);
    xnor g1786(n2365 ,n2298 ,n2318);
    nand g1787(n1253 ,n28[0] ,n1195);
    xnor g1788(n4323 ,n4272 ,n4303);
    nand g1789(n4346 ,n4345 ,n4330);
    not g1790(n3884 ,n3883);
    nand g1791(n1761 ,n1658 ,n1702);
    nand g1792(n6105 ,n6047 ,n6072);
    nor g1793(n1597 ,n1568 ,n19[5]);
    nor g1794(n5546 ,n5363 ,n5452);
    nor g1795(n2765 ,n2638 ,n2693);
    nand g1796(n1239 ,n1097 ,n737);
    nand g1797(n4990 ,n4518 ,n4814);
    nor g1798(n725 ,n610 ,n710);
    nor g1799(n2460 ,n2361 ,n2421);
    xnor g1800(n3786 ,n3559 ,n3560);
    nand g1801(n6305 ,n6555 ,n6251);
    nor g1802(n2339 ,n2267 ,n2310);
    nor g1803(n2787 ,n2650 ,n2725);
    or g1804(n3286 ,n3281 ,n3269);
    not g1805(n5458 ,n5457);
    nand g1806(n2346 ,n2309 ,n2295);
    not g1807(n1579 ,n1578);
    xnor g1808(n2876 ,n2747 ,n2658);
    xnor g1809(n2287 ,n2227 ,n2118);
    xnor g1810(n6594 ,n3216 ,n3235);
    dff g1811(.RN(n1), .SN(1'b1), .CK(n0), .D(n1350), .Q(n23[12]));
    dff g1812(.RN(n1), .SN(1'b1), .CK(n0), .D(n1392), .Q(n21[7]));
    nand g1813(n5100 ,n4754 ,n5034);
    xnor g1814(n2895 ,n2778 ,n2852);
    or g1815(n6060 ,n5882 ,n6037);
    not g1816(n2915 ,n2914);
    nand g1817(n5394 ,n5173 ,n5176);
    nor g1818(n3017 ,n2969 ,n2992);
    nand g1819(n4800 ,n4585 ,n4608);
    not g1820(n723 ,n724);
    xor g1821(n5864 ,n5781 ,n5814);
    nand g1822(n4853 ,n4609 ,n4630);
    xnor g1823(n3411 ,n39[4] ,n6553);
    nand g1824(n445 ,n355 ,n432);
    xnor g1825(n404 ,n304 ,n352);
    nand g1826(n3312 ,n3290 ,n3311);
    xnor g1827(n6581 ,n2021 ,n2042);
    nand g1828(n1115 ,n32[1] ,n555);
    nor g1829(n436 ,n353 ,n415);
    nand g1830(n850 ,n1505 ,n714);
    nand g1831(n1204 ,n812 ,n739);
    xnor g1832(n6159 ,n6079 ,n6128);
    nand g1833(n434 ,n356 ,n410);
    xnor g1834(n6560 ,n4343 ,n4348);
    not g1835(n3544 ,n3543);
    nor g1836(n5369 ,n5132 ,n5163);
    nand g1837(n4660 ,n21[3] ,n4371);
    nand g1838(n3239 ,n3210 ,n3238);
    nand g1839(n2356 ,n2233 ,n2292);
    not g1840(n5413 ,n5396);
    xnor g1841(n4210 ,n4140 ,n4065);
    nand g1842(n2560 ,n2532 ,n2559);
    nand g1843(n5025 ,n4544 ,n4826);
    nand g1844(n4125 ,n4025 ,n4057);
    dff g1845(.RN(n1), .SN(1'b1), .CK(n0), .D(n1397), .Q(n27[12]));
    nor g1846(n2760 ,n2653 ,n2691);
    xnor g1847(n6603 ,n3404 ,n3427);
    xnor g1848(n5191 ,n4929 ,n4487);
    xnor g1849(n1536 ,n102 ,n84);
    or g1850(n749 ,n555 ,n683);
    buf g1851(n13[2], n10[2]);
    not g1852(n3691 ,n3690);
    dff g1853(.RN(n1), .SN(1'b1), .CK(n0), .D(n1412), .Q(n20[5]));
    nand g1854(n2583 ,n40[14] ,n6525);
    xnor g1855(n392 ,n218 ,n343);
    xnor g1856(n6553 ,n4177 ,n4155);
    xnor g1857(n3172 ,n3123 ,n38[3]);
    nand g1858(n1268 ,n849 ,n1014);
    nand g1859(n2251 ,n2166 ,n2192);
    nand g1860(n5487 ,n5405 ,n5398);
    xnor g1861(n2927 ,n2867 ,n2766);
    nor g1862(n333 ,n241 ,n293);
    xor g1863(n295 ,n198 ,n229);
    nand g1864(n5502 ,n5266 ,n5374);
    nand g1865(n2246 ,n2143 ,n2199);
    nand g1866(n4307 ,n4219 ,n4281);
    nand g1867(n1703 ,n1577 ,n1677);
    xnor g1868(n4266 ,n4195 ,n4228);
    nand g1869(n6294 ,n40[4] ,n6250);
    nand g1870(n2083 ,n21[2] ,n2065);
    nand g1871(n5741 ,n5504 ,n5661);
    xnor g1872(n6127 ,n6087 ,n6082);
    or g1873(n2279 ,n2234 ,n2232);
    nand g1874(n903 ,n23[13] ,n715);
    nand g1875(n1272 ,n852 ,n1021);
    nand g1876(n2094 ,n6534 ,n2085);
    not g1877(n2736 ,n2735);
    nor g1878(n3430 ,n3409 ,n3429);
    nand g1879(n3923 ,n3869 ,n3837);
    nand g1880(n6387 ,n6245 ,n6256);
    nor g1881(n6262 ,n6236 ,n6252);
    nand g1882(n1391 ,n946 ,n1147);
    nor g1883(n3438 ,n3407 ,n3437);
    nand g1884(n1178 ,n5[0] ,n557);
    nand g1885(n6317 ,n6502 ,n6249);
    nand g1886(n5845 ,n5617 ,n5801);
    nand g1887(n535 ,n499 ,n526);
    xnor g1888(n2422 ,n2366 ,n2392);
    nand g1889(n6281 ,n40[1] ,n6250);
    nor g1890(n6459 ,n6417 ,n6416);
    xnor g1891(n4332 ,n4310 ,n4318);
    nor g1892(n2382 ,n2301 ,n2343);
    xnor g1893(n2543 ,n2528 ,n2513);
    nand g1894(n283 ,n192 ,n226);
    or g1895(n4769 ,n4629 ,n4424);
    not g1896(n3268 ,n37[1]);
    nor g1897(n2886 ,n2767 ,n2816);
    or g1898(n2934 ,n2853 ,n2897);
    nand g1899(n6306 ,n41[15] ,n6254);
    nor g1900(n4693 ,n4395 ,n4406);
    nand g1901(n4812 ,n4574 ,n4468);
    nand g1902(n3820 ,n3553 ,n3706);
    nand g1903(n1731 ,n1579 ,n1700);
    nand g1904(n6309 ,n40[6] ,n6250);
    nor g1905(n2696 ,n2566 ,n2623);
    nor g1906(n6259 ,n6230 ,n6252);
    xor g1907(n4947 ,n4538 ,n4484);
    nor g1908(n2127 ,n2085 ,n2113);
    nand g1909(n3828 ,n3626 ,n3698);
    xnor g1910(n4113 ,n4012 ,n3906);
    xnor g1911(n3951 ,n3842 ,n3859);
    or g1912(n5739 ,n5571 ,n5688);
    not g1913(n5530 ,n5529);
    nand g1914(n4454 ,n21[4] ,n4389);
    or g1915(n5335 ,n5286 ,n5159);
    not g1916(n3254 ,n37[7]);
    dff g1917(.RN(n1), .SN(1'b1), .CK(n0), .D(n1427), .Q(n26[1]));
    dff g1918(.RN(n1), .SN(1'b1), .CK(n0), .D(n1403), .Q(n33[15]));
    nand g1919(n3363 ,n3359 ,n3362);
    nor g1920(n1917 ,n1853 ,n1892);
    nand g1921(n138 ,n32[3] ,n137);
    nand g1922(n986 ,n20[2] ,n714);
    not g1923(n2561 ,n2560);
    nand g1924(n3313 ,n3301 ,n3312);
    nor g1925(n3793 ,n3544 ,n3689);
    not g1926(n3487 ,n36[6]);
    or g1927(n2569 ,n40[11] ,n6522);
    nand g1928(n878 ,n34[13] ,n717);
    not g1929(n3473 ,n37[1]);
    nand g1930(n1387 ,n641 ,n777);
    nor g1931(n4531 ,n4406 ,n4405);
    xnor g1932(n2375 ,n2270 ,n2296);
    not g1933(n5783 ,n5782);
    nand g1934(n1445 ,n1017 ,n1269);
    nand g1935(n997 ,n4[4] ,n713);
    nand g1936(n819 ,n23[4] ,n715);
    nand g1937(n287 ,n183 ,n212);
    nand g1938(n3874 ,n3650 ,n3798);
    not g1939(n55 ,n54);
    xnor g1940(n319 ,n233 ,n179);
    nor g1941(n2809 ,n2704 ,n2757);
    nand g1942(n5756 ,n5560 ,n5678);
    nand g1943(n276 ,n213 ,n214);
    nand g1944(n3518 ,n3468 ,n3484);
    not g1945(n2416 ,n2415);
    nand g1946(n1599 ,n1564 ,n1572);
    nand g1947(n3962 ,n3848 ,n3890);
    nor g1948(n6231 ,n41[12] ,n6592);
    nand g1949(n2970 ,n2812 ,n2934);
    xnor g1950(n5932 ,n5817 ,n5776);
    nand g1951(n4048 ,n3928 ,n3966);
    not g1952(n5189 ,n5188);
    nand g1953(n6328 ,n6542 ,n6248);
    not g1954(n4006 ,n3990);
    nand g1955(n1690 ,n1582 ,n1654);
    nand g1956(n937 ,n28[6] ,n717);
    xnor g1957(n6599 ,n3402 ,n3435);
    nand g1958(n6100 ,n6040 ,n6081);
    nand g1959(n3120 ,n6573 ,n6550);
    nor g1960(n4524 ,n4402 ,n4418);
    nor g1961(n2552 ,n2515 ,n2551);
    nand g1962(n5682 ,n5495 ,n5528);
    nand g1963(n6296 ,n6554 ,n6251);
    not g1964(n3447 ,n3446);
    nor g1965(n581 ,n34[8] ,n34[15]);
    not g1966(n59 ,n58);
    dff g1967(.RN(n1), .SN(1'b1), .CK(n0), .D(n1336), .Q(n24[5]));
    not g1968(n2565 ,n6528);
    nor g1969(n3427 ,n3388 ,n3426);
    nand g1970(n5121 ,n4769 ,n5046);
    nand g1971(n1965 ,n1861 ,n1943);
    xnor g1972(n1883 ,n1830 ,n1811);
    nand g1973(n6416 ,n6283 ,n6331);
    nand g1974(n817 ,n23[6] ,n715);
    nor g1975(n2403 ,n2338 ,n2382);
    nand g1976(n4000 ,n3838 ,n3933);
    xnor g1977(n3971 ,n3831 ,n3855);
    or g1978(n4074 ,n4043 ,n3972);
    xnor g1979(n1605 ,n1560 ,n19[7]);
    nor g1980(n4789 ,n4555 ,n4539);
    nand g1981(n2978 ,n2957 ,n2946);
    nand g1982(n5985 ,n5907 ,n5929);
    not g1983(n1907 ,n1906);
    xor g1984(n4923 ,n4508 ,n4475);
    nand g1985(n866 ,n33[13] ,n712);
    nor g1986(n1835 ,n1637 ,n1827);
    nand g1987(n1377 ,n624 ,n762);
    nor g1988(n837 ,n567 ,n721);
    nand g1989(n768 ,n724 ,n691);
    nor g1990(n2717 ,n2566 ,n2629);
    nand g1991(n35[7] ,n6449 ,n6481);
    xnor g1992(n6084 ,n6037 ,n5882);
    nand g1993(n1066 ,n10[14] ,n711);
    nor g1994(n2808 ,n2670 ,n2762);
    nand g1995(n1295 ,n1050 ,n872);
    nor g1996(n5552 ,n5372 ,n5450);
    nor g1997(n6486 ,n6394 ,n6472);
    nand g1998(n2843 ,n2734 ,n2778);
    not g1999(n4386 ,n4385);
    xnor g2000(n6031 ,n5956 ,n5883);
    xor g2001(n6524 ,n6586 ,n6563);
    not g2002(n3460 ,n3459);
    nor g2003(n833 ,n561 ,n721);
    nand g2004(n4639 ,n4382 ,n20[3]);
    nand g2005(n892 ,n33[4] ,n712);
    nand g2006(n4691 ,n20[1] ,n4373);
    nand g2007(n1060 ,n11[3] ,n711);
    nand g2008(n804 ,n35[7] ,n712);
    nor g2009(n2436 ,n2409 ,n2394);
    nand g2010(n805 ,n35[6] ,n712);
    nand g2011(n1166 ,n20[0] ,n722);
    nand g2012(n4087 ,n3978 ,n4038);
    xnor g2013(n1774 ,n1721 ,n1637);
    nand g2014(n1630 ,n1599 ,n1609);
    xnor g2015(n2442 ,n2391 ,n2412);
    nand g2016(n4583 ,n20[5] ,n4363);
    xnor g2017(n6555 ,n4264 ,n4277);
    or g2018(n5514 ,n5277 ,n5460);
    xnor g2019(n3902 ,n3747 ,n3512);
    nand g2020(n854 ,n1502 ,n714);
    nand g2021(n6368 ,n6493 ,n6253);
    xnor g2022(n1785 ,n1724 ,n1645);
    nand g2023(n3139 ,n6561 ,n3103);
    nand g2024(n4425 ,n21[2] ,n4365);
    nand g2025(n1689 ,n1577 ,n1654);
    nand g2026(n6376 ,n38[5] ,n6246);
    nand g2027(n911 ,n1548 ,n554);
    nand g2028(n5365 ,n5145 ,n5238);
    nand g2029(n1113 ,n32[2] ,n710);
    nand g2030(n2164 ,n6540 ,n2122);
    nand g2031(n3872 ,n3649 ,n3823);
    nand g2032(n4664 ,n21[0] ,n4371);
    dff g2033(.RN(n1), .SN(1'b1), .CK(n0), .D(n1286), .Q(n16[0]));
    buf g2034(n13[12], n10[12]);
    nor g2035(n6465 ,n6434 ,n6432);
    nand g2036(n4162 ,n4047 ,n4098);
    nor g2037(n4530 ,n4411 ,n4413);
    nand g2038(n4030 ,n3870 ,n3994);
    nand g2039(n5981 ,n5908 ,n5932);
    xnor g2040(n3337 ,n6570 ,n6582);
    xnor g2041(n4957 ,n4652 ,n4700);
    nand g2042(n3450 ,n3447 ,n19[2]);
    not g2043(n1997 ,n1996);
    nand g2044(n3631 ,n3478 ,n19[5]);
    nand g2045(n6415 ,n6282 ,n6339);
    dff g2046(.RN(n1), .SN(1'b1), .CK(n0), .D(n1311), .Q(n10[11]));
    nand g2047(n437 ,n420 ,n402);
    or g2048(n2576 ,n40[0] ,n6511);
    not g2049(n4382 ,n4381);
    nand g2050(n5028 ,n4654 ,n4839);
    xnor g2051(n5643 ,n5423 ,n5295);
    xnor g2052(n6054 ,n5991 ,n6003);
    nand g2053(n6272 ,n6564 ,n6251);
    nand g2054(n1767 ,n1689 ,n1705);
    nand g2055(n1421 ,n988 ,n1174);
    nand g2056(n1003 ,n12[13] ,n710);
    nand g2057(n1189 ,n10[7] ,n555);
    not g2058(n3485 ,n3490);
    nor g2059(n2458 ,n2335 ,n2426);
    dff g2060(.RN(n1), .SN(1'b1), .CK(n0), .D(n1359), .Q(n23[9]));
    nand g2061(n4598 ,n21[1] ,n4384);
    xnor g2062(n5311 ,n5067 ,n4793);
    xnor g2063(n498 ,n465 ,n450);
    buf g2064(n15[2], n15[6]);
    nand g2065(n4443 ,n21[6] ,n4386);
    xnor g2066(n5636 ,n5421 ,n5229);
    dff g2067(.RN(n1), .SN(1'b1), .CK(n0), .D(n1405), .Q(n21[2]));
    nor g2068(n2722 ,n2565 ,n2617);
    nand g2069(n5945 ,n5854 ,n5892);
    xnor g2070(n6556 ,n4301 ,n4311);
    nor g2071(n3395 ,n6555 ,n39[6]);
    nand g2072(n3611 ,n3485 ,n19[5]);
    nand g2073(n5554 ,n5209 ,n5454);
    or g2074(n396 ,n363 ,n361);
    nand g2075(n5757 ,n5567 ,n5674);
    xnor g2076(n3755 ,n3504 ,n3608);
    nand g2077(n4832 ,n4641 ,n4600);
    nor g2078(n5591 ,n5324 ,n5466);
    nand g2079(n1203 ,n829 ,n793);
    nand g2080(n4836 ,n4588 ,n4626);
    not g2081(n1647 ,n1648);
    nand g2082(n2904 ,n2839 ,n2890);
    nor g2083(n250 ,n179 ,n228);
    xnor g2084(n4061 ,n3952 ,n3941);
    nor g2085(n4784 ,n4679 ,n4675);
    nand g2086(n1326 ,n925 ,n1081);
    not g2087(n4669 ,n4668);
    xnor g2088(n4937 ,n4567 ,n4590);
    not g2089(n3336 ,n3335);
    nand g2090(n4431 ,n20[4] ,n4361);
    or g2091(n5242 ,n5113 ,n5086);
    xnor g2092(n3173 ,n3129 ,n6552);
    nand g2093(n863 ,n1514 ,n714);
    nand g2094(n1419 ,n797 ,n1173);
    xnor g2095(n6204 ,n6188 ,n6194);
    nand g2096(n6053 ,n5984 ,n6009);
    nand g2097(n3605 ,n3478 ,n19[7]);
    nor g2098(n5363 ,n5112 ,n5202);
    nand g2099(n1143 ,n22[1] ,n720);
    not g2100(n4388 ,n4387);
    or g2101(n4738 ,n4489 ,n4633);
    nand g2102(n3358 ,n3354 ,n3357);
    dff g2103(.RN(n1), .SN(1'b1), .CK(n0), .D(n1276), .Q(n1502));
    nand g2104(n5496 ,n5260 ,n5355);
    nand g2105(n4539 ,n21[7] ,n4369);
    nand g2106(n5570 ,n5359 ,n5479);
    nor g2107(n5448 ,n5299 ,n5373);
    xor g2108(n40[11] ,n6600 ,n38[12]);
    nand g2109(n4201 ,n4132 ,n4164);
    nor g2110(n6232 ,n41[13] ,n6591);
    xnor g2111(n314 ,n203 ,n201);
    or g2112(n748 ,n555 ,n686);
    nand g2113(n5658 ,n5527 ,n5536);
    or g2114(n4283 ,n4209 ,n4268);
    not g2115(n3266 ,n37[3]);
    xor g2116(n40[3] ,n38[4] ,n6608);
    not g2117(n4646 ,n4645);
    nand g2118(n5810 ,n5562 ,n5732);
    not g2119(n2750 ,n2749);
    nand g2120(n2155 ,n6533 ,n2126);
    nor g2121(n2478 ,n2423 ,n2447);
    nand g2122(n6337 ,n38[1] ,n6246);
    nand g2123(n3969 ,n3836 ,n3923);
    nand g2124(n179 ,n163 ,n148);
    xnor g2125(n5593 ,n5172 ,n5502);
    xnor g2126(n4026 ,n3881 ,n3689);
    nand g2127(n6019 ,n5925 ,n5988);
    nand g2128(n5730 ,n5575 ,n5627);
    or g2129(n486 ,n451 ,n461);
    nand g2130(n2594 ,n40[4] ,n6515);
    nand g2131(n4602 ,n21[2] ,n4386);
    nand g2132(n1435 ,n929 ,n1209);
    xnor g2133(n1633 ,n1597 ,n1608);
    nand g2134(n6445 ,n6308 ,n6377);
    nand g2135(n3314 ,n3293 ,n3313);
    nor g2136(n2976 ,n2928 ,n2947);
    nand g2137(n178 ,n172 ,n155);
    dff g2138(.RN(n1), .SN(1'b1), .CK(n0), .D(n1346), .Q(n23[15]));
    nand g2139(n945 ,n21[7] ,n714);
    xnor g2140(n6509 ,n3072 ,n3089);
    xnor g2141(n2447 ,n2303 ,n2402);
    nand g2142(n6215 ,n6206 ,n6214);
    nand g2143(n6117 ,n6041 ,n6100);
    nand g2144(n5733 ,n5605 ,n5606);
    nand g2145(n6224 ,n25[2] ,n25[1]);
    xnor g2146(n3213 ,n3157 ,n3172);
    xnor g2147(n5641 ,n5418 ,n5098);
    or g2148(n4708 ,n4598 ,n4610);
    xnor g2149(n6583 ,n2039 ,n2046);
    nor g2150(n585 ,n34[1] ,n34[7]);
    not g2151(n4379 ,n36[6]);
    xnor g2152(n4891 ,n4616 ,n4472);
    nor g2153(n106 ,n24[1] ,n24[0]);
    not g2154(n3483 ,n36[0]);
    nand g2155(n5849 ,n5815 ,n5730);
    nand g2156(n5059 ,n4778 ,n4954);
    xnor g2157(n3775 ,n3591 ,n3501);
    xor g2158(n3948 ,n3858 ,n3871);
    nand g2159(n970 ,n27[7] ,n715);
    xnor g2160(n680 ,n35[5] ,n31[5]);
    not g2161(n2673 ,n2672);
    nand g2162(n180 ,n165 ,n144);
    not g2163(n2529 ,n2528);
    nand g2164(n820 ,n23[3] ,n715);
    nand g2165(n2000 ,n1955 ,n1984);
    nand g2166(n5993 ,n5889 ,n5947);
    or g2167(n3648 ,n3586 ,n3595);
    nor g2168(n575 ,n34[2] ,n34[3]);
    nor g2169(n2774 ,n2671 ,n2739);
    or g2170(n3968 ,n3907 ,n3940);
    xnor g2171(n5825 ,n5696 ,n5724);
    nand g2172(n4570 ,n21[7] ,n4384);
    nor g2173(n2778 ,n2608 ,n2712);
    xnor g2174(n2523 ,n2500 ,n2492);
    nor g2175(n6180 ,n6161 ,n6148);
    or g2176(n4740 ,n4631 ,n4439);
    xnor g2177(n3049 ,n3008 ,n3024);
    xnor g2178(n5167 ,n4898 ,n4640);
    not g2179(n2796 ,n2795);
    nor g2180(n572 ,n33[5] ,n35[5]);
    xnor g2181(n3773 ,n3587 ,n3592);
    nand g2182(n433 ,n366 ,n404);
    xnor g2183(n5202 ,n4905 ,n4592);
    nand g2184(n1056 ,n11[6] ,n711);
    nand g2185(n1460 ,n920 ,n1379);
    nand g2186(n35[5] ,n6469 ,n6482);
    xnor g2187(n1848 ,n1754 ,n1793);
    or g2188(n3649 ,n3516 ,n3548);
    dff g2189(.RN(n1), .SN(1'b1), .CK(n0), .D(n1306), .Q(n11[0]));
    nand g2190(n3319 ,n6580 ,n41[7]);
    nand g2191(n5087 ,n4732 ,n5042);
    nand g2192(n6340 ,n6496 ,n6249);
    nand g2193(n3177 ,n38[1] ,n3155);
    nor g2194(n2655 ,n2565 ,n2593);
    or g2195(n4730 ,n4562 ,n4591);
    not g2196(n2998 ,n2990);
    nor g2197(n397 ,n338 ,n375);
    dff g2198(.RN(n1), .SN(1'b1), .CK(n0), .D(n1297), .Q(n11[8]));
    not g2199(n3526 ,n3525);
    nor g2200(n4698 ,n4411 ,n4396);
    nand g2201(n4998 ,n4677 ,n4817);
    nand g2202(n1078 ,n27[12] ,n718);
    nand g2203(n4684 ,n21[0] ,n4369);
    nand g2204(n2037 ,n2018 ,n2024);
    not g2205(n5626 ,n5625);
    nand g2206(n1744 ,n1674 ,n1710);
    xor g2207(n4904 ,n4673 ,n4500);
    xnor g2208(n1526 ,n531 ,n535);
    xnor g2209(n4109 ,n4013 ,n4028);
    xnor g2210(n308 ,n243 ,n206);
    nand g2211(n3724 ,n3538 ,n3505);
    nor g2212(n2682 ,n2565 ,n2628);
    not g2213(n6033 ,n6032);
    xnor g2214(n1991 ,n1945 ,n1926);
    nand g2215(n1217 ,n924 ,n768);
    not g2216(n1566 ,n1565);
    nor g2217(n2801 ,n2646 ,n2723);
    or g2218(n3668 ,n3514 ,n3510);
    nor g2219(n3817 ,n3611 ,n3736);
    or g2220(n2065 ,n20[2] ,n20[1]);
    xnor g2221(n1881 ,n1831 ,n1794);
    nand g2222(n3048 ,n3013 ,n3021);
    xnor g2223(n1798 ,n1759 ,n1646);
    nand g2224(n6174 ,n6152 ,n6137);
    nand g2225(n1459 ,n901 ,n1377);
    nand g2226(n6339 ,n38[9] ,n6246);
    nor g2227(n4665 ,n4412 ,n4410);
    nand g2228(n813 ,n34[6] ,n717);
    not g2229(n2451 ,n2450);
    nand g2230(n6405 ,n6264 ,n6330);
    nand g2231(n1399 ,n964 ,n1155);
    xnor g2232(n5963 ,n5777 ,n5872);
    or g2233(n2806 ,n2774 ,n2801);
    or g2234(n1787 ,n1750 ,n1747);
    xnor g2235(n1926 ,n1872 ,n1829);
    xnor g2236(n4300 ,n4245 ,n4270);
    not g2237(n5130 ,n5129);
    nand g2238(n1001 ,n12[14] ,n711);
    nor g2239(n340 ,n268 ,n312);
    nand g2240(n1090 ,n33[14] ,n710);
    not g2241(n2465 ,n2456);
    nand g2242(n3850 ,n3670 ,n3803);
    nor g2243(n777 ,n600 ,n720);
    xnor g2244(n3176 ,n3125 ,n38[13]);
    or g2245(n737 ,n555 ,n680);
    nand g2246(n3540 ,n3478 ,n19[1]);
    nand g2247(n4590 ,n20[1] ,n4371);
    xnor g2248(n2804 ,n2709 ,n2634);
    xnor g2249(n2315 ,n2257 ,n2119);
    nand g2250(n1068 ,n10[12] ,n711);
    xnor g2251(n3066 ,n3033 ,n3026);
    not g2252(n317 ,n316);
    xnor g2253(n2087 ,n20[3] ,n21[3]);
    nand g2254(n4573 ,n4380 ,n20[2]);
    nand g2255(n2344 ,n2318 ,n2285);
    nand g2256(n5903 ,n5804 ,n5826);
    nand g2257(n5988 ,n5856 ,n5938);
    or g2258(n714 ,n18[2] ,n579);
    dff g2259(.RN(n1), .SN(1'b1), .CK(n0), .D(n1240), .Q(n33[3]));
    nand g2260(n5477 ,n5151 ,n5334);
    nand g2261(n6333 ,n6495 ,n6249);
    nand g2262(n5053 ,n4692 ,n4813);
    nand g2263(n4603 ,n20[7] ,n4373);
    not g2264(n2361 ,n2360);
    or g2265(n3677 ,n3603 ,n3513);
    nor g2266(n3433 ,n3389 ,n3432);
    nand g2267(n5392 ,n5167 ,n5184);
    nand g2268(n1788 ,n1750 ,n1747);
    xnor g2269(n5877 ,n5765 ,n5527);
    or g2270(n74 ,n69 ,n57);
    xnor g2271(n3365 ,n3363 ,n6579);
    not g2272(n4069 ,n4068);
    nand g2273(n5020 ,n4683 ,n4815);
    xnor g2274(n3893 ,n3749 ,n3549);
    nand g2275(n35[8] ,n6453 ,n6451);
    nand g2276(n1071 ,n10[9] ,n710);
    xnor g2277(n38[4] ,n2467 ,n2462);
    nor g2278(n2639 ,n2566 ,n2590);
    nand g2279(n2162 ,n6535 ,n2127);
    nor g2280(n5788 ,n5591 ,n5713);
    nor g2281(n4671 ,n4409 ,n4415);
    xnor g2282(n6203 ,n6187 ,n6180);
    or g2283(n4072 ,n3988 ,n4029);
    nand g2284(n545 ,n533 ,n544);
    xnor g2285(n3407 ,n6562 ,n6547);
    not g2286(n148 ,n147);
    or g2287(n2067 ,n20[6] ,n20[5]);
    nand g2288(n5857 ,n5731 ,n5787);
    nand g2289(n1669 ,n1580 ,n1651);
    or g2290(n6073 ,n5992 ,n6030);
    nand g2291(n3857 ,n3725 ,n3785);
    nand g2292(n1681 ,n1576 ,n1652);
    nand g2293(n6372 ,n6500 ,n6249);
    nand g2294(n5989 ,n5901 ,n5944);
    or g2295(n4131 ,n3892 ,n4056);
    xnor g2296(n478 ,n417 ,n448);
    nand g2297(n4822 ,n4582 ,n4637);
    nand g2298(n832 ,n34[3] ,n717);
    nor g2299(n5452 ,n5218 ,n5362);
    or g2300(n259 ,n192 ,n226);
    not g2301(n4418 ,n4369);
    nand g2302(n2630 ,n2591 ,n2571);
    or g2303(n6010 ,n5873 ,n5973);
    xor g2304(n2122 ,n2106 ,n2112);
    xnor g2305(n5961 ,n5878 ,n5785);
    not g2306(n3278 ,n36[5]);
    nand g2307(n4449 ,n21[1] ,n4369);
    xnor g2308(n6537 ,n3310 ,n3294);
    not g2309(n5608 ,n5607);
    or g2310(n1936 ,n1883 ,n1903);
    or g2311(n4252 ,n4195 ,n4228);
    nand g2312(n5854 ,n5708 ,n5792);
    nand g2313(n625 ,n17[2] ,n26[2]);
    nand g2314(n1727 ,n1621 ,n1682);
    nor g2315(n2054 ,n2015 ,n2053);
    or g2316(n4296 ,n4226 ,n4273);
    nand g2317(n4068 ,n3968 ,n4035);
    not g2318(n5723 ,n5722);
    nor g2319(n5559 ,n5494 ,n5499);
    nand g2320(n1345 ,n1138 ,n950);
    nand g2321(n3228 ,n3185 ,n3227);
    nand g2322(n3143 ,n6559 ,n3095);
    nand g2323(n4624 ,n21[1] ,n4374);
    nand g2324(n3339 ,n6574 ,n3323);
    not g2325(n4954 ,n4953);
    not g2326(n2006 ,n2005);
    nand g2327(n2822 ,n2728 ,n2749);
    nand g2328(n2092 ,n6539 ,n2085);
    nand g2329(n1610 ,n19[2] ,n1596);
    nand g2330(n1980 ,n1956 ,n1923);
    nand g2331(n109 ,n107 ,n106);
    nand g2332(n1249 ,n1137 ,n772);
    nor g2333(n3315 ,n3296 ,n3314);
    nand g2334(n4419 ,n20[7] ,n4361);
    nor g2335(n760 ,n604 ,n720);
    not g2336(n3688 ,n3687);
    nand g2337(n5122 ,n4764 ,n5047);
    nand g2338(n3927 ,n3523 ,n3845);
    xnor g2339(n6590 ,n3224 ,n3251);
    nor g2340(n740 ,n700 ,n708);
    nor g2341(n3553 ,n3487 ,n3498);
    xnor g2342(n5692 ,n5528 ,n5495);
    or g2343(n880 ,n715 ,n697);
    xnor g2344(n5178 ,n4887 ,n4635);
    not g2345(n3739 ,n3723);
    nand g2346(n2088 ,n6533 ,n2085);
    nand g2347(n869 ,n1511 ,n714);
    not g2348(n3496 ,n3478);
    nand g2349(n2091 ,n6536 ,n2085);
    xnor g2350(n3035 ,n3000 ,n2950);
    nand g2351(n3032 ,n2993 ,n3014);
    xnor g2352(n673 ,n35[13] ,n33[13]);
    nor g2353(n5372 ,n5083 ,n5188);
    nand g2354(n3985 ,n3938 ,n3937);
    nand g2355(n632 ,n22[3] ,n26[3]);
    xnor g2356(n2081 ,n21[2] ,n21[1]);
    xnor g2357(n678 ,n35[2] ,n33[2]);
    nor g2358(n3695 ,n3541 ,n3545);
    xnor g2359(n463 ,n427 ,n443);
    nand g2360(n1073 ,n1536 ,n713);
    nor g2361(n2556 ,n2555 ,n2541);
    nand g2362(n2029 ,n2006 ,n2013);
    nor g2363(n342 ,n260 ,n329);
    nand g2364(n4848 ,n4631 ,n4439);
    xnor g2365(n2120 ,n2103 ,n2077);
    nand g2366(n1210 ,n34[4] ,n834);
    xnor g2367(n2318 ,n2258 ,n2119);
    xnor g2368(n5693 ,n5539 ,n5504);
    nand g2369(n1458 ,n1125 ,n1374);
    nand g2370(n2171 ,n6541 ,n2121);
    nor g2371(n5707 ,n5530 ,n5618);
    or g2372(n4713 ,n4461 ,n4594);
    nor g2373(n1853 ,n1819 ,n1800);
    nand g2374(n3119 ,n6579 ,n6556);
    nor g2375(n288 ,n199 ,n197);
    nor g2376(n2909 ,n2841 ,n2883);
    nand g2377(n3149 ,n6563 ,n3096);
    nand g2378(n924 ,n30[1] ,n723);
    xnor g2379(n5631 ,n5424 ,n5227);
    not g2380(n1868 ,n1867);
    or g2381(n378 ,n288 ,n341);
    nand g2382(n1304 ,n1061 ,n809);
    nand g2383(n1096 ,n1519 ,n716);
    dff g2384(.RN(n1), .SN(1'b1), .CK(n0), .D(n1479), .Q(n17[5]));
    not g2385(n144 ,n174);
    dff g2386(.RN(n1), .SN(1'b1), .CK(n0), .D(n1418), .Q(n16[7]));
    xnor g2387(n2493 ,n2397 ,n2442);
    nor g2388(n2015 ,n2003 ,n1995);
    nand g2389(n239 ,n172 ,n144);
    xnor g2390(n1648 ,n1630 ,n1606);
    xnor g2391(n5421 ,n5179 ,n5182);
    xor g2392(n6516 ,n6578 ,n6555);
    nand g2393(n1287 ,n1040 ,n865);
    xnor g2394(n3880 ,n3781 ,n3531);
    xnor g2395(n5786 ,n5596 ,n5642);
    nor g2396(n764 ,n573 ,n723);
    nand g2397(n909 ,n1546 ,n712);
    not g2398(n3273 ,n3272);
    nor g2399(n2395 ,n2261 ,n2378);
    nand g2400(n5114 ,n4775 ,n5020);
    xnor g2401(n6558 ,n4333 ,n4344);
    xnor g2402(n2972 ,n2942 ,n2938);
    nor g2403(n2850 ,n2769 ,n2764);
    nand g2404(n1082 ,n32[6] ,n555);
    nand g2405(n1136 ,n22[4] ,n720);
    xnor g2406(n1930 ,n1873 ,n1558);
    not g2407(n3637 ,n3636);
    xnor g2408(n5306 ,n4419 ,n5096);
    nor g2409(n5728 ,n5578 ,n5613);
    nand g2410(n1151 ,n23[13] ,n716);
    nor g2411(n4547 ,n4401 ,n4403);
    dff g2412(.RN(n1), .SN(1'b1), .CK(n0), .D(n1422), .Q(n26[4]));
    nand g2413(n2250 ,n2172 ,n2218);
    nand g2414(n5343 ,n5116 ,n5174);
    xor g2415(n5294 ,n4952 ,n4471);
    nand g2416(n345 ,n262 ,n328);
    nand g2417(n4459 ,n21[7] ,n4361);
    nand g2418(n5129 ,n4767 ,n5026);
    nand g2419(n3086 ,n3064 ,n3085);
    xnor g2420(n6113 ,n6054 ,n6081);
    xnor g2421(n4221 ,n4183 ,n4196);
    xor g2422(n40[12] ,n6599 ,n38[13]);
    or g2423(n3670 ,n3524 ,n3542);
    nand g2424(n6285 ,n6565 ,n6254);
    not g2425(n3284 ,n36[2]);
    nand g2426(n1360 ,n1113 ,n911);
    or g2427(n5316 ,n5173 ,n5176);
    not g2428(n1574 ,n1573);
    nand g2429(n517 ,n482 ,n502);
    nand g2430(n1620 ,n1577 ,n1612);
    not g2431(n268 ,n267);
    nand g2432(n1764 ,n1673 ,n1715);
    or g2433(n4706 ,n4473 ,n4604);
    nand g2434(n4150 ,n4066 ,n4108);
    xnor g2435(n4959 ,n4655 ,n4656);
    xnor g2436(n2444 ,n2398 ,n2403);
    nand g2437(n1348 ,n643 ,n735);
    or g2438(n3034 ,n3008 ,n3024);
    nand g2439(n5949 ,n5793 ,n5867);
    nand g2440(n5115 ,n4735 ,n4997);
    nand g2441(n6240 ,n41[15] ,n6589);
    not g2442(n5181 ,n5180);
    xnor g2443(n5594 ,n5460 ,n5277);
    xnor g2444(n6561 ,n4341 ,n4350);
    nand g2445(n1464 ,n1134 ,n1383);
    xnor g2446(n5528 ,n5311 ,n5093);
    or g2447(n6205 ,n6195 ,n6184);
    dff g2448(.RN(n1), .SN(1'b1), .CK(n0), .D(n1324), .Q(n10[1]));
    dff g2449(.RN(n1), .SN(1'b1), .CK(n0), .D(n1416), .Q(n16[8]));
    nand g2450(n5106 ,n4857 ,n4967);
    nand g2451(n1918 ,n1857 ,n1899);
    not g2452(n2425 ,n2424);
    nor g2453(n2937 ,n2829 ,n2898);
    nand g2454(n6344 ,n6508 ,n6249);
    nor g2455(n2844 ,n2731 ,n2793);
    or g2456(n3098 ,n6580 ,n6557);
    nor g2457(n6250 ,n6227 ,n6222);
    dff g2458(.RN(n1), .SN(1'b1), .CK(n0), .D(n1450), .Q(n34[3]));
    nand g2459(n1248 ,n28[5] ,n1193);
    xnor g2460(n5784 ,n5599 ,n5588);
    or g2461(n5797 ,n5632 ,n5751);
    nand g2462(n5678 ,n5507 ,n5564);
    nor g2463(n6256 ,n6229 ,n6252);
    not g2464(n1748 ,n1749);
    nand g2465(n4218 ,n4148 ,n4189);
    or g2466(n2574 ,n40[1] ,n6512);
    nor g2467(n3687 ,n3638 ,n3625);
    nand g2468(n3517 ,n3468 ,n3481);
    nand g2469(n1379 ,n626 ,n764);
    nor g2470(n5464 ,n5229 ,n5412);
    xnor g2471(n4921 ,n4430 ,n4617);
    nand g2472(n3819 ,n3642 ,n3728);
    nand g2473(n4700 ,n21[7] ,n4373);
    nand g2474(n4038 ,n3875 ,n3967);
    nand g2475(n989 ,n20[0] ,n714);
    nand g2476(n3109 ,n6578 ,n6555);
    nor g2477(n4653 ,n4393 ,n4414);
    nand g2478(n6304 ,n6572 ,n6254);
    nor g2479(n2784 ,n2601 ,n2686);
    nor g2480(n4690 ,n4410 ,n4402);
    nor g2481(n2043 ,n2010 ,n2042);
    xnor g2482(n1808 ,n1742 ,n1646);
    nand g2483(n502 ,n458 ,n491);
    nand g2484(n1717 ,n1588 ,n1676);
    nand g2485(n1172 ,n5[2] ,n713);
    nand g2486(n1356 ,n1109 ,n908);
    nand g2487(n435 ,n345 ,n408);
    nor g2488(n3681 ,n3645 ,n3646);
    xnor g2489(n6531 ,n3441 ,n3401);
    nand g2490(n2456 ,n2398 ,n2419);
    nand g2491(n1327 ,n1079 ,n960);
    xnor g2492(n679 ,n23[2] ,n34[2]);
    not g2493(n4406 ,n4378);
    xnor g2494(n3360 ,n3358 ,n6578);
    nor g2495(n2512 ,n2472 ,n2488);
    nand g2496(n2991 ,n2918 ,n2950);
    xnor g2497(n5959 ,n5869 ,n5834);
    nand g2498(n2139 ,n6535 ,n2123);
    or g2499(n5748 ,n5605 ,n5606);
    nor g2500(n2840 ,n2667 ,n2783);
    not g2501(n4152 ,n4151);
    xnor g2502(n364 ,n306 ,n215);
    nand g2503(n1417 ,n986 ,n1172);
    nand g2504(n4619 ,n21[3] ,n4380);
    nand g2505(n1279 ,n856 ,n1028);
    xnor g2506(n3409 ,n6558 ,n6543);
    nand g2507(n1099 ,n27[14] ,n718);
    nand g2508(n5670 ,n5352 ,n5519);
    nand g2509(n4562 ,n4378 ,n20[4]);
    not g2510(n5536 ,n5535);
    nand g2511(n2046 ,n2029 ,n2045);
    or g2512(n4776 ,n4632 ,n4480);
    nand g2513(n5939 ,n5800 ,n5871);
    not g2514(n3479 ,n36[1]);
    not g2515(n2668 ,n2667);
    nand g2516(n1250 ,n1140 ,n775);
    nand g2517(n3853 ,n3675 ,n3800);
    xnor g2518(n6587 ,n2055 ,n2009);
    nor g2519(n4080 ,n3976 ,n4020);
    or g2520(n4240 ,n4171 ,n4205);
    nand g2521(n5047 ,n4665 ,n4865);
    nand g2522(n6156 ,n6099 ,n6133);
    not g2523(n3264 ,n37[0]);
    not g2524(n152 ,n151);
    or g2525(n432 ,n366 ,n404);
    not g2526(n4380 ,n4379);
    xnor g2527(n6021 ,n5951 ,n5989);
    nand g2528(n5743 ,n5583 ,n5664);
    nand g2529(n6169 ,n6154 ,n6113);
    not g2530(n4106 ,n4105);
    nand g2531(n186 ,n167 ,n144);
    nor g2532(n329 ,n196 ,n292);
    or g2533(n2547 ,n2510 ,n2546);
    xnor g2534(n2261 ,n2108 ,n2207);
    xor g2535(n4889 ,n4506 ,n4444);
    not g2536(n4090 ,n4089);
    nand g2537(n5785 ,n5667 ,n5726);
    nand g2538(n6154 ,n6136 ,n6119);
    nand g2539(n5846 ,n5755 ,n5789);
    nor g2540(n1985 ,n1850 ,n1960);
    nor g2541(n3317 ,n3297 ,n3316);
    or g2542(n4725 ,n4615 ,n4471);
    or g2543(n3666 ,n3585 ,n3607);
    nand g2544(n5334 ,n4878 ,n5161);
    or g2545(n3457 ,n3452 ,n3456);
    nand g2546(n1658 ,n1582 ,n1651);
    xnor g2547(n685 ,n35[7] ,n31[7]);
    nand g2548(n1691 ,n1576 ,n1649);
    nand g2549(n3925 ,n3830 ,n3867);
    not g2550(n1992 ,n1991);
    nand g2551(n5262 ,n5117 ,n5076);
    nand g2552(n5542 ,n5322 ,n5474);
    nand g2553(n1477 ,n826 ,n1251);
    xnor g2554(n5883 ,n5766 ,n5647);
    nand g2555(n830 ,n17[6] ,n721);
    xnor g2556(n5782 ,n5600 ,n5639);
    nand g2557(n3519 ,n3476 ,n19[1]);
    dff g2558(.RN(n1), .SN(1'b1), .CK(n0), .D(n1221), .Q(n28[3]));
    or g2559(n3096 ,n38[13] ,n6586);
    nand g2560(n2102 ,n2070 ,n2083);
    xnor g2561(n1820 ,n1769 ,n1645);
    nor g2562(n2713 ,n2568 ,n2621);
    xnor g2563(n5531 ,n5300 ,n5095);
    not g2564(n3846 ,n3845);
    dff g2565(.RN(n1), .SN(1'b1), .CK(n0), .D(n1247), .Q(n22[4]));
    nand g2566(n5144 ,n4797 ,n5022);
    xnor g2567(n6128 ,n6085 ,n6067);
    nor g2568(n5821 ,n5811 ,n5720);
    nand g2569(n4277 ,n4237 ,n4261);
    nand g2570(n1347 ,n902 ,n1096);
    nand g2571(n979 ,n27[3] ,n715);
    not g2572(n5203 ,n5202);
    nand g2573(n966 ,n21[3] ,n714);
    nor g2574(n103 ,n84 ,n102);
    nor g2575(n601 ,n33[11] ,n35[11]);
    nand g2576(n5952 ,n5848 ,n5905);
    not g2577(n5291 ,n5290);
    nor g2578(n2701 ,n2565 ,n2622);
    or g2579(n2580 ,n40[10] ,n6521);
    nand g2580(n4643 ,n21[2] ,n4389);
    xor g2581(n4903 ,n4701 ,n4490);
    buf g2582(n13[15], n10[15]);
    not g2583(n3467 ,n37[2]);
    nor g2584(n5718 ,n5609 ,n5689);
    nand g2585(n1373 ,n824 ,n1019);
    nand g2586(n3967 ,n3841 ,n3897);
    nand g2587(n5125 ,n4749 ,n4995);
    nand g2588(n4975 ,n4663 ,n4795);
    xor g2589(n1558 ,n1795 ,n1783);
    nor g2590(n1902 ,n1777 ,n1881);
    nand g2591(n4805 ,n4622 ,n4474);
    nor g2592(n2692 ,n2566 ,n2625);
    xnor g2593(n1809 ,n1646 ,n1752);
    nor g2594(n3318 ,n6576 ,n6568);
    or g2595(n3653 ,n3532 ,n3529);
    nand g2596(n5482 ,n5148 ,n5379);
    xnor g2597(n5193 ,n4973 ,n4445);
    xnor g2598(n2420 ,n2374 ,n2312);
    nor g2599(n761 ,n597 ,n720);
    nand g2600(n1914 ,n1864 ,n1893);
    nor g2601(n2697 ,n2566 ,n2619);
    not g2602(n3606 ,n3605);
    or g2603(n5716 ,n5534 ,n5633);
    xnor g2604(n1555 ,n24[2] ,n122);
    xnor g2605(n2857 ,n2755 ,n2781);
    xnor g2606(n3298 ,n3281 ,n3269);
    nand g2607(n417 ,n252 ,n383);
    not g2608(n4394 ,n21[5]);
    nand g2609(n1471 ,n967 ,n1404);
    xnor g2610(n5159 ,n4892 ,n4680);
    xnor g2611(n6606 ,n3413 ,n3421);
    nand g2612(n5471 ,n5403 ,n5288);
    dff g2613(.RN(n1), .SN(1'b1), .CK(n0), .D(n1444), .Q(n12[9]));
    nand g2614(n939 ,n28[4] ,n717);
    nand g2615(n3804 ,n3635 ,n3707);
    nor g2616(n570 ,n33[10] ,n35[10]);
    not g2617(n2731 ,n2730);
    nand g2618(n1112 ,n32[3] ,n710);
    not g2619(n2343 ,n2337);
    nor g2620(n2766 ,n2652 ,n2692);
    dff g2621(.RN(n1), .SN(1'b1), .CK(n0), .D(n1266), .Q(n16[4]));
    xnor g2622(n5281 ,n4921 ,n4536);
    nand g2623(n938 ,n28[5] ,n717);
    nand g2624(n6265 ,n41[6] ,n6254);
    nand g2625(n350 ,n256 ,n324);
    xnor g2626(n5187 ,n4883 ,n4483);
    nand g2627(n4181 ,n4106 ,n4151);
    nand g2628(n1720 ,n1579 ,n1677);
    nand g2629(n1244 ,n1007 ,n759);
    or g2630(n5319 ,n5171 ,n5170);
    nand g2631(n1331 ,n1013 ,n895);
    not g2632(n160 ,n36[0]);
    nand g2633(n4345 ,n4329 ,n4344);
    or g2634(n5839 ,n5631 ,n5776);
    nand g2635(n4627 ,n4386 ,n20[6]);
    nand g2636(n6326 ,n6573 ,n6247);
    nor g2637(n2660 ,n2568 ,n2587);
    nand g2638(n5468 ,n5214 ,n5390);
    xnor g2639(n2372 ,n2293 ,n2288);
    dff g2640(.RN(n1), .SN(1'b1), .CK(n0), .D(n1438), .Q(n29[2]));
    nor g2641(n4657 ,n4394 ,n4391);
    xnor g2642(n5777 ,n5593 ,n5459);
    nor g2643(n3627 ,n3488 ,n3494);
    xnor g2644(n3950 ,n3522 ,n3845);
    nand g2645(n3991 ,n3907 ,n3940);
    nand g2646(n1212 ,n34[2] ,n835);
    not g2647(n565 ,n17[6]);
    nand g2648(n1045 ,n2[3] ,n557);
    nand g2649(n2587 ,n40[3] ,n6514);
    xnor g2650(n2297 ,n2243 ,n2120);
    nand g2651(n331 ,n208 ,n278);
    xnor g2652(n4271 ,n4222 ,n4207);
    nand g2653(n4593 ,n21[4] ,n4361);
    nor g2654(n2648 ,n2565 ,n2589);
    nand g2655(n1276 ,n854 ,n1026);
    not g2656(n1827 ,n1826);
    nand g2657(n1396 ,n887 ,n1151);
    not g2658(n2618 ,n2619);
    nand g2659(n5009 ,n4530 ,n4812);
    nand g2660(n3987 ,n3906 ,n3905);
    nor g2661(n2852 ,n2676 ,n2799);
    not g2662(n4401 ,n20[3]);
    nand g2663(n3861 ,n3655 ,n3810);
    nand g2664(n3979 ,n3860 ,n3941);
    or g2665(n4797 ,n4486 ,n4475);
    nand g2666(n1243 ,n1035 ,n755);
    xnor g2667(n3129 ,n38[2] ,n6575);
    nand g2668(n2979 ,n2970 ,n2963);
    xnor g2669(n2391 ,n2323 ,n2299);
    xnor g2670(n508 ,n473 ,n485);
    nor g2671(n2539 ,n2503 ,n2527);
    xor g2672(n6522 ,n6584 ,n6561);
    nand g2673(n1638 ,n1615 ,n1631);
    or g2674(n5333 ,n5210 ,n5283);
    nand g2675(n514 ,n466 ,n506);
    or g2676(n5937 ,n5785 ,n5878);
    nand g2677(n806 ,n35[5] ,n554);
    nor g2678(n3010 ,n2968 ,n2995);
    nand g2679(n890 ,n1547 ,n712);
    or g2680(n3647 ,n3533 ,n3581);
    not g2681(n4114 ,n4113);
    or g2682(n3958 ,n3906 ,n3905);
    nor g2683(n6457 ,n6415 ,n6411);
    nor g2684(n2347 ,n2309 ,n2295);
    nand g2685(n1759 ,n1668 ,n1713);
    or g2686(n4796 ,n4607 ,n4643);
    nand g2687(n6283 ,n6552 ,n6251);
    buf g2688(n13[4], n11[4]);
    nand g2689(n5484 ,n5098 ,n5384);
    not g2690(n1576 ,n1575);
    nand g2691(n6198 ,n6180 ,n6187);
    xnor g2692(n6563 ,n4322 ,n4354);
    nand g2693(n503 ,n459 ,n486);
    xnor g2694(n5418 ,n5186 ,n5187);
    xnor g2695(n1873 ,n1806 ,n1828);
    nand g2696(n1443 ,n1012 ,n1264);
    nor g2697(n5704 ,n5529 ,n5619);
    nand g2698(n2230 ,n2139 ,n2212);
    or g2699(n114 ,n32[4] ,n32[3]);
    nor g2700(n2153 ,n2109 ,n2125);
    xnor g2701(n2919 ,n2861 ,n2891);
    nor g2702(n6455 ,n6410 ,n6409);
    nand g2703(n3863 ,n3664 ,n3811);
    nand g2704(n5480 ,n5087 ,n5367);
    not g2705(n4391 ,n36[2]);
    xnor g2706(n5301 ,n5069 ,n5075);
    nor g2707(n2394 ,n2262 ,n2379);
    xnor g2708(n2913 ,n2890 ,n2792);
    buf g2709(n36[0] ,n1508);
    xor g2710(n2115 ,n2099 ,n2077);
    xnor g2711(n668 ,n19[1] ,n27[1]);
    nor g2712(n2849 ,n2740 ,n2803);
    nor g2713(n618 ,n19[3] ,n27[3]);
    nand g2714(n3629 ,n3476 ,n19[0]);
    xnor g2715(n2524 ,n2495 ,n2481);
    nand g2716(n1274 ,n855 ,n1025);
    nand g2717(n2101 ,n6541 ,n2085);
    or g2718(n4036 ,n3943 ,n4004);
    nand g2719(n3548 ,n3474 ,n3484);
    nand g2720(n3013 ,n2983 ,n2982);
    or g2721(n5653 ,n5495 ,n5528);
    nand g2722(n1246 ,n28[6] ,n1192);
    xnor g2723(n1602 ,n19[6] ,n19[5]);
    nor g2724(n3391 ,n6558 ,n6543);
    nand g2725(n1054 ,n11[7] ,n711);
    nor g2726(n1938 ,n1557 ,n1907);
    nand g2727(n1318 ,n1075 ,n891);
    xnor g2728(n4154 ,n4051 ,n4002);
    nand g2729(n971 ,n27[6] ,n715);
    nand g2730(n3347 ,n3339 ,n3346);
    nand g2731(n1184 ,n4[6] ,n713);
    nor g2732(n450 ,n406 ,n436);
    nand g2733(n3717 ,n3503 ,n3519);
    nand g2734(n3153 ,n3099 ,n3140);
    nor g2735(n588 ,n34[4] ,n34[11]);
    nand g2736(n1180 ,n1535 ,n713);
    xnor g2737(n496 ,n464 ,n441);
    or g2738(n3448 ,n3443 ,n19[1]);
    or g2739(n4767 ,n4609 ,n4630);
    xnor g2740(n5699 ,n5552 ,n5501);
    nand g2741(n3118 ,n38[9] ,n6582);
    nand g2742(n3730 ,n3586 ,n3595);
    dff g2743(.RN(n1), .SN(1'b1), .CK(n0), .D(n1343), .Q(n24[1]));
    nand g2744(n1104 ,n33[1] ,n710);
    nor g2745(n1483 ,n617 ,n1201);
    not g2746(n225 ,n224);
    or g2747(n3957 ,n3896 ,n3895);
    nand g2748(n4607 ,n21[0] ,n4378);
    nor g2749(n2905 ,n2811 ,n2874);
    nand g2750(n494 ,n453 ,n471);
    nand g2751(n2133 ,n6539 ,n2122);
    or g2752(n2430 ,n2396 ,n2399);
    nand g2753(n6279 ,n6566 ,n6254);
    nand g2754(n5253 ,n4419 ,n5078);
    nand g2755(n1211 ,n34[3] ,n837);
    nand g2756(n1756 ,n1670 ,n1733);
    nand g2757(n6474 ,n6378 ,n6437);
    xnor g2758(n6147 ,n6089 ,n6112);
    nor g2759(n2645 ,n2566 ,n2595);
    or g2760(n5325 ,n5219 ,n5234);
    nor g2761(n786 ,n574 ,n715);
    nand g2762(n1092 ,n1556 ,n716);
    or g2763(n2572 ,n40[7] ,n6518);
    nand g2764(n5079 ,n4747 ,n5048);
    nand g2765(n6437 ,n6240 ,n6257);
    nor g2766(n1892 ,n1808 ,n1869);
    not g2767(n5624 ,n5623);
    nand g2768(n5822 ,n5805 ,n5784);
    xor g2769(n4930 ,n4654 ,n4450);
    nand g2770(n5383 ,n5166 ,n5165);
    not g2771(n69 ,n68);
    xnor g2772(n5761 ,n5646 ,n5547);
    or g2773(n3656 ,n3515 ,n3600);
    nand g2774(n549 ,n509 ,n548);
    nand g2775(n934 ,n34[10] ,n717);
    xnor g2776(n6597 ,n3410 ,n3439);
    xnor g2777(n2376 ,n2304 ,n2315);
    nor g2778(n2770 ,n2648 ,n2695);
    nand g2779(n1290 ,n1044 ,n867);
    or g2780(n3674 ,n3579 ,n3527);
    nor g2781(n4557 ,n4397 ,n4403);
    xnor g2782(n5832 ,n5691 ,n5584);
    nor g2783(n2521 ,n2484 ,n2498);
    xnor g2784(n6544 ,n3342 ,n3376);
    nand g2785(n5270 ,n5113 ,n5086);
    buf g2786(n14[8], n11[8]);
    not g2787(n4969 ,n4968);
    nor g2788(n3684 ,n3570 ,n3643);
    nand g2789(n2207 ,n2091 ,n2162);
    xnor g2790(n2107 ,n2068 ,n2079);
    xnor g2791(n5629 ,n5414 ,n5097);
    xnor g2792(n3168 ,n3121 ,n38[15]);
    xnor g2793(n6086 ,n6032 ,n6052);
    nand g2794(n2145 ,n6534 ,n2123);
    nand g2795(n3581 ,n3482 ,n19[1]);
    not g2796(n5969 ,n5968);
    nand g2797(n1232 ,n1020 ,n727);
    nor g2798(n75 ,n59 ,n43);
    dff g2799(.RN(n1), .SN(1'b1), .CK(n0), .D(n1435), .Q(n29[5]));
    nand g2800(n2168 ,n6537 ,n2126);
    nand g2801(n3532 ,n3468 ,n3480);
    nor g2802(n1667 ,n1590 ,n1650);
    or g2803(n731 ,n555 ,n678);
    nand g2804(n543 ,n532 ,n542);
    xnor g2805(n5182 ,n4888 ,n4452);
    xnor g2806(n6499 ,n3020 ,n3009);
    nand g2807(n5815 ,n5683 ,n5741);
    not g2808(n4049 ,n4037);
    nand g2809(n490 ,n441 ,n464);
    nand g2810(n6239 ,n41[13] ,n6591);
    nor g2811(n3841 ,n3667 ,n3827);
    nand g2812(n5124 ,n4715 ,n5037);
    nand g2813(n1470 ,n894 ,n1389);
    dff g2814(.RN(n1), .SN(1'b1), .CK(n0), .D(n1202), .Q(n17[2]));
    nand g2815(n4845 ,n4501 ,n4573);
    nand g2816(n578 ,n566 ,n561);
    or g2817(n4282 ,n4230 ,n4274);
    not g2818(n3361 ,n3360);
    nor g2819(n2649 ,n2565 ,n2585);
    xnor g2820(n304 ,n186 ,n216);
    not g2821(n1846 ,n1845);
    nand g2822(n5580 ,n5316 ,n5485);
    nand g2823(n5011 ,n4701 ,n4875);
    or g2824(n1214 ,n564 ,n1133);
    nand g2825(n3867 ,n3694 ,n3828);
    not g2826(n3494 ,n19[2]);
    xnor g2827(n3170 ,n3122 ,n38[9]);
    xnor g2828(n3947 ,n3863 ,n3861);
    xnor g2829(n1987 ,n1952 ,n1924);
    nand g2830(n6438 ,n6242 ,n6260);
    nand g2831(n5476 ,n5298 ,n5399);
    nand g2832(n2243 ,n2133 ,n2181);
    nand g2833(n4440 ,n21[5] ,n4365);
    nand g2834(n1150 ,n6[6] ,n713);
    nand g2835(n4854 ,n4423 ,n4458);
    dff g2836(.RN(n1), .SN(1'b1), .CK(n0), .D(n1243), .Q(n31[5]));
    not g2837(n5870 ,n5869);
    xnor g2838(n5433 ,n5161 ,n4877);
    nand g2839(n3157 ,n3107 ,n3141);
    nor g2840(n270 ,n202 ,n236);
    or g2841(n793 ,n637 ,n721);
    xnor g2842(n3452 ,n3447 ,n19[2]);
    nand g2843(n3321 ,n6584 ,n6572);
    nand g2844(n2096 ,n6540 ,n2085);
    nand g2845(n2209 ,n2094 ,n2161);
    nor g2846(n2278 ,n2109 ,n2229);
    nand g2847(n914 ,n30[7] ,n723);
    xnor g2848(n4141 ,n4063 ,n3939);
    xnor g2849(n375 ,n295 ,n184);
    nor g2850(n1966 ,n1789 ,n1937);
    xnor g2851(n5930 ,n5818 ,n5836);
    not g2852(n5545 ,n5544);
    xnor g2853(n2861 ,n2787 ,n2737);
    nand g2854(n4600 ,n4382 ,n20[2]);
    xnor g2855(n2039 ,n2025 ,n2019);
    not g2856(n1559 ,n37[7]);
    nor g2857(n2534 ,n2454 ,n2509);
    or g2858(n3196 ,n3158 ,n3179);
    xnor g2859(n5773 ,n5623 ,n5687);
    nor g2860(n2789 ,n2598 ,n2699);
    xnor g2861(n3122 ,n6559 ,n6582);
    not g2862(n6226 ,n25[2]);
    xnor g2863(n5553 ,n5305 ,n5099);
    or g2864(n6134 ,n6070 ,n6116);
    nand g2865(n2130 ,n6539 ,n2123);
    nand g2866(n143 ,n32[6] ,n142);
    nand g2867(n3643 ,n3474 ,n3486);
    xnor g2868(n5928 ,n5773 ,n5837);
    xnor g2869(n4184 ,n4097 ,n4080);
    nand g2870(n1369 ,n632 ,n758);
    nor g2871(n2026 ,n2006 ,n2013);
    nand g2872(n2428 ,n2396 ,n2399);
    nand g2873(n5582 ,n5339 ,n5476);
    dff g2874(.RN(n1), .SN(1'b1), .CK(n0), .D(n1340), .Q(n24[2]));
    nand g2875(n3512 ,n3460 ,n3481);
    xnor g2876(n41[7] ,n6176 ,n6185);
    xnor g2877(n511 ,n477 ,n461);
    or g2878(n5926 ,n5800 ,n5871);
    not g2879(n166 ,n36[3]);
    nor g2880(n1625 ,n1601 ,n1614);
    nor g2881(n2902 ,n2808 ,n2880);
    nand g2882(n1000 ,n4[3] ,n713);
    nand g2883(n5252 ,n4420 ,n5077);
    xnor g2884(n2948 ,n2864 ,n2900);
    xnor g2885(n6494 ,n3221 ,n3245);
    xnor g2886(n2426 ,n2368 ,n2295);
    xnor g2887(n2285 ,n2246 ,n2118);
    nand g2888(n4273 ,n4240 ,n4253);
    nand g2889(n5708 ,n5542 ,n5615);
    xnor g2890(n3938 ,n3763 ,n3611);
    nand g2891(n3084 ,n3058 ,n3083);
    nor g2892(n5321 ,n5182 ,n5179);
    nor g2893(n4519 ,n4407 ,n4416);
    nor g2894(n2329 ,n2268 ,n2311);
    nand g2895(n2892 ,n2777 ,n2806);
    not g2896(n2123 ,n2124);
    nand g2897(n6414 ,n6273 ,n6322);
    xnor g2898(n1314 ,n715 ,n24[0]);
    nand g2899(n420 ,n336 ,n384);
    or g2900(n577 ,n22[2] ,n22[3]);
    nand g2901(n6242 ,n41[5] ,n6595);
    nand g2902(n1704 ,n1584 ,n1675);
    buf g2903(n14[4], n10[4]);
    nand g2904(n4317 ,n4280 ,n4311);
    xor g2905(n4926 ,n4518 ,n4591);
    nor g2906(n2767 ,n2614 ,n2684);
    or g2907(n4148 ,n4060 ,n4104);
    xnor g2908(n4179 ,n4113 ,n4091);
    nand g2909(n1724 ,n1576 ,n1677);
    nor g2910(n5729 ,n5687 ,n5624);
    or g2911(n2838 ,n2786 ,n2760);
    dff g2912(.RN(n1), .SN(1'b1), .CK(n0), .D(n1296), .Q(n1509));
    nand g2913(n2942 ,n2830 ,n2907);
    xnor g2914(n1616 ,n1570 ,n19[2]);
    nand g2915(n3081 ,n3063 ,n3080);
    nand g2916(n5942 ,n5850 ,n5880);
    nand g2917(n5807 ,n5566 ,n5712);
    dff g2918(.RN(n1), .SN(1'b1), .CK(n0), .D(n1270), .Q(n1505));
    or g2919(n1981 ,n1922 ,n1951);
    nand g2920(n771 ,n724 ,n693);
    buf g2921(n37[7] ,n1507);
    nand g2922(n6365 ,n39[4] ,n6248);
    xnor g2923(n2025 ,n1988 ,n1965);
    dff g2924(.RN(n1), .SN(1'b1), .CK(n0), .D(n1227), .Q(n27[1]));
    nand g2925(n1632 ,n1600 ,n1611);
    nor g2926(n2995 ,n2924 ,n2949);
    xnor g2927(n3069 ,n3040 ,n3030);
    xnor g2928(n2914 ,n2863 ,n2798);
    nand g2929(n2140 ,n6538 ,n2121);
    xnor g2930(n6139 ,n6093 ,n6115);
    xnor g2931(n3914 ,n3772 ,n3573);
    nor g2932(n4877 ,n4655 ,n4656);
    xnor g2933(n1923 ,n1871 ,n1785);
    nand g2934(n4829 ,n4563 ,n4440);
    nand g2935(n950 ,n35[8] ,n712);
    nand g2936(n5683 ,n5500 ,n5539);
    nand g2937(n3227 ,n3177 ,n3225);
    or g2938(n4716 ,n4483 ,n4595);
    nand g2939(n3019 ,n2960 ,n2987);
    not g2940(n2785 ,n2784);
    nor g2941(n3397 ,n6561 ,n6546);
    nand g2942(n1091 ,n33[11] ,n710);
    nand g2943(n1771 ,n1694 ,n1712);
    xnor g2944(n1828 ,n1772 ,n1645);
    dff g2945(.RN(n1), .SN(1'b1), .CK(n0), .D(n1440), .Q(n17[0]));
    nand g2946(n541 ,n521 ,n540);
    nand g2947(n6263 ,n6556 ,n6251);
    nand g2948(n3534 ,n3482 ,n19[2]);
    nand g2949(n3823 ,n3624 ,n3705);
    nand g2950(n5500 ,n5270 ,n5371);
    xnor g2951(n6503 ,n3070 ,n3077);
    or g2952(n6190 ,n6165 ,n6183);
    or g2953(n4313 ,n4286 ,n4309);
    not g2954(n3265 ,n3264);
    or g2955(n5275 ,n5068 ,n5074);
    xnor g2956(n6497 ,n2912 ,n2849);
    nor g2957(n2720 ,n2566 ,n2622);
    nand g2958(n3609 ,n3466 ,n3481);
    xnor g2959(n6140 ,n6117 ,n6023);
    xnor g2960(n1814 ,n1747 ,n1749);
    xnor g2961(n6066 ,n5996 ,n6008);
    dff g2962(.RN(n1), .SN(1'b1), .CK(n0), .D(n1478), .Q(n17[3]));
    nand g2963(n2964 ,n2929 ,n2920);
    nand g2964(n534 ,n517 ,n523);
    or g2965(n4775 ,n4593 ,n4431);
    nand g2966(n5726 ,n5553 ,n5670);
    nand g2967(n6301 ,n40[5] ,n6250);
    xnor g2968(n5190 ,n4948 ,n4601);
    not g2969(n2855 ,n2847);
    nor g2970(n615 ,n23[6] ,n34[6]);
    nor g2971(n4054 ,n3883 ,n4024);
    xnor g2972(n3885 ,n3758 ,n3601);
    nand g2973(n624 ,n17[6] ,n26[6]);
    nand g2974(n4001 ,n3659 ,n3934);
    nor g2975(n2710 ,n2565 ,n2629);
    nor g2976(n2977 ,n2918 ,n2950);
    xnor g2977(n2378 ,n2321 ,n2282);
    nand g2978(n4987 ,n4672 ,n4866);
    nor g2979(n3421 ,n3392 ,n3420);
    xnor g2980(n1753 ,n1656 ,n1648);
    nand g2981(n35[15] ,n6470 ,n6483);
    nand g2982(n1153 ,n23[12] ,n716);
    nand g2983(n5795 ,n5582 ,n5739);
    nand g2984(n3845 ,n3672 ,n3826);
    nand g2985(n1134 ,n22[5] ,n720);
    not g2986(n2324 ,n2323);
    xnor g2987(n2544 ,n2527 ,n2502);
    nand g2988(n6220 ,n6219 ,n6162);
    xor g2989(n4952 ,n4524 ,n4615);
    nand g2990(n6463 ,n6379 ,n6444);
    nor g2991(n2314 ,n2273 ,n2283);
    nor g2992(n3618 ,n3492 ,n3494);
    nand g2993(n1075 ,n10[5] ,n555);
    nand g2994(n1600 ,n1562 ,n1568);
    xor g2995(n1519 ,n444 ,n552);
    xnor g2996(n3939 ,n3762 ,n3551);
    not g2997(n1746 ,n1747);
    nand g2998(n5254 ,n4784 ,n5084);
    not g2999(n567 ,n17[3]);
    nand g3000(n6273 ,n6562 ,n6251);
    nand g3001(n207 ,n163 ,n146);
    nand g3002(n3698 ,n3517 ,n3594);
    nor g3003(n2476 ,n2459 ,n2462);
    not g3004(n2229 ,n2230);
    or g3005(n3150 ,n3120 ,n3097);
    nor g3006(n2725 ,n2566 ,n2626);
    nand g3007(n1353 ,n1107 ,n906);
    not g3008(n5573 ,n5572);
    nand g3009(n3249 ,n3200 ,n3248);
    nand g3010(n6434 ,n6368 ,n6366);
    nand g3011(n3289 ,n3283 ,n3265);
    xnor g3012(n5914 ,n5807 ,n5825);
    not g3013(n4404 ,n20[4]);
    dff g3014(.RN(n1), .SN(1'b1), .CK(n0), .D(n1309), .Q(n10[13]));
    xor g3015(n39[0] ,n6618 ,n38[0]);
    xnor g3016(n2486 ,n2415 ,n2448);
    not g3017(n1564 ,n1563);
    nand g3018(n2584 ,n40[0] ,n6511);
    nand g3019(n5267 ,n5118 ,n5107);
    xnor g3020(n2973 ,n2940 ,n2939);
    nand g3021(n4472 ,n4386 ,n20[0]);
    not g3022(n1909 ,n1908);
    dff g3023(.RN(n1), .SN(1'b1), .CK(n0), .D(n1465), .Q(n28[7]));
    not g3024(n5615 ,n5614);
    nor g3025(n2721 ,n2568 ,n2620);
    nand g3026(n861 ,n1515 ,n714);
    or g3027(n4763 ,n4445 ,n4470);
    nand g3028(n2144 ,n6537 ,n2121);
    dff g3029(.RN(n1), .SN(1'b1), .CK(n0), .D(n1398), .Q(n27[11]));
    nor g3030(n769 ,n612 ,n720);
    xnor g3031(n4023 ,n3880 ,n3872);
    nand g3032(n708 ,n569 ,n588);
    not g3033(n2664 ,n2663);
    nand g3034(n5983 ,n5853 ,n5937);
    xnor g3035(n6582 ,n2044 ,n2032);
    nand g3036(n1145 ,n22[0] ,n720);
    nand g3037(n1051 ,n1527 ,n716);
    nand g3038(n97 ,n92 ,n96);
    nor g3039(n3016 ,n2967 ,n2999);
    nor g3040(n1837 ,n1636 ,n1826);
    not g3041(n1563 ,n37[4]);
    nor g3042(n2897 ,n2824 ,n2884);
    nand g3043(n1414 ,n981 ,n1170);
    or g3044(n4766 ,n4478 ,n4493);
    buf g3045(n13[9], n10[9]);
    nand g3046(n3062 ,n3028 ,n3039);
    dff g3047(.RN(n1), .SN(1'b1), .CK(n0), .D(n1414), .Q(n20[4]));
    xnor g3048(n1793 ,n1726 ,n1646);
    xnor g3049(n669 ,n21[2] ,n30[2]);
    xnor g3050(n1824 ,n1645 ,n1770);
    nor g3051(n2674 ,n2568 ,n2593);
    nand g3052(n4167 ,n4083 ,n4114);
    nand g3053(n6209 ,n6182 ,n6207);
    nand g3054(n915 ,n23[15] ,n715);
    nor g3055(n2016 ,n1986 ,n1996);
    xnor g3056(n2473 ,n2370 ,n2426);
    nand g3057(n4578 ,n21[7] ,n4367);
    nor g3058(n1894 ,n1832 ,n1838);
    xnor g3059(n3174 ,n3124 ,n38[4]);
    not g3060(n715 ,n716);
    nor g3061(n4171 ,n4049 ,n4122);
    nand g3062(n801 ,n26[2] ,n723);
    nand g3063(n3310 ,n3291 ,n3309);
    nand g3064(n3206 ,n3160 ,n3171);
    not g3065(n3270 ,n36[7]);
    nand g3066(n1142 ,n33[9] ,n555);
    nand g3067(n4824 ,n4484 ,n4479);
    nor g3068(n2470 ,n2415 ,n2449);
    xnor g3069(n4185 ,n4094 ,n4048);
    xor g3070(n4883 ,n4648 ,n4595);
    nand g3071(n218 ,n169 ,n146);
    nand g3072(n1297 ,n1052 ,n874);
    or g3073(n3065 ,n3027 ,n3036);
    nand g3074(n6269 ,n40[12] ,n6250);
    nand g3075(n5750 ,n5569 ,n5610);
    nor g3076(n5837 ,n5707 ,n5774);
    nand g3077(n4487 ,n21[5] ,n4380);
    xnor g3078(n6532 ,n4263 ,n4358);
    dff g3079(.RN(n1), .SN(1'b1), .CK(n0), .D(n1446), .Q(n12[5]));
    nor g3080(n4670 ,n4412 ,n4413);
    nand g3081(n6325 ,n38[8] ,n6246);
    not g3082(n2501 ,n2500);
    xnor g3083(n5875 ,n5764 ,n5549);
    nand g3084(n1640 ,n1606 ,n1630);
    nand g3085(n197 ,n159 ,n153);
    dff g3086(.RN(n1), .SN(1'b1), .CK(n0), .D(n1461), .Q(n22[7]));
    nand g3087(n1723 ,n1620 ,n1698);
    nand g3088(n6277 ,n6550 ,n6251);
    nand g3089(n6079 ,n5981 ,n6042);
    nor g3090(n2737 ,n2567 ,n2621);
    xnor g3091(n5186 ,n4893 ,n4493);
    nand g3092(n4193 ,n4130 ,n4163);
    not g3093(n3735 ,n3710);
    nand g3094(n1148 ,n6[7] ,n713);
    or g3095(n4774 ,n4425 ,n4644);
    nand g3096(n4526 ,n21[5] ,n4374);
    dff g3097(.RN(n1), .SN(1'b1), .CK(n0), .D(n1329), .Q(n10[2]));
    nor g3098(n4509 ,n4408 ,n4416);
    nand g3099(n5705 ,n5646 ,n5672);
    nand g3100(n5404 ,n4977 ,n5264);
    nand g3101(n3645 ,n3470 ,n3484);
    nand g3102(n4019 ,n3903 ,n3973);
    nand g3103(n654 ,n16[8] ,n23[8]);
    nor g3104(n3690 ,n3565 ,n3641);
    xnor g3105(n697 ,n23[5] ,n16[5]);
    nand g3106(n5498 ,n5261 ,n5356);
    xnor g3107(n2951 ,n2856 ,n2910);
    nand g3108(n3458 ,n3450 ,n3457);
    xnor g3109(n5885 ,n5760 ,n5754);
    dff g3110(.RN(n1), .SN(1'b1), .CK(n0), .D(n1459), .Q(n30[6]));
    nand g3111(n4427 ,n20[2] ,n4369);
    or g3112(n3963 ,n3843 ,n3898);
    nand g3113(n6221 ,n6169 ,n6220);
    not g3114(n3499 ,n19[5]);
    nand g3115(n5023 ,n4510 ,n4806);
    or g3116(n4726 ,n4582 ,n4637);
    xor g3117(n5781 ,n5597 ,n5507);
    nand g3118(n349 ,n286 ,n317);
    nand g3119(n3620 ,n3485 ,n19[7]);
    nand g3120(n5850 ,n5747 ,n5794);
    xnor g3121(n6087 ,n5968 ,n6051);
    nand g3122(n4516 ,n21[1] ,n4378);
    nand g3123(n3346 ,n6566 ,n3345);
    or g3124(n1855 ,n1828 ,n1806);
    nor g3125(n4511 ,n4409 ,n4399);
    nand g3126(n5052 ,n4525 ,n4823);
    nand g3127(n4995 ,n4689 ,n4808);
    nor g3128(n2786 ,n2606 ,n2700);
    nor g3129(n2514 ,n2470 ,n2499);
    nand g3130(n868 ,n1512 ,n714);
    dff g3131(.RN(n1), .SN(1'b1), .CK(n0), .D(n1314), .Q(n24[0]));
    nand g3132(n2847 ,n2797 ,n2761);
    nand g3133(n1266 ,n846 ,n1010);
    nand g3134(n3619 ,n3470 ,n3481);
    or g3135(n416 ,n308 ,n370);
    nand g3136(n1209 ,n34[5] ,n833);
    nand g3137(n2185 ,n6533 ,n2148);
    or g3138(n2819 ,n2743 ,n2765);
    nand g3139(n1012 ,n12[10] ,n555);
    nor g3140(n612 ,n21[5] ,n30[5]);
    nand g3141(n2131 ,n6535 ,n2122);
    nor g3142(n2385 ,n2237 ,n2355);
    xnor g3143(n5691 ,n5491 ,n5570);
    xnor g3144(n5226 ,n4918 ,n4558);
    nand g3145(n6402 ,n6285 ,n6329);
    nor g3146(n5057 ,n4981 ,n4963);
    xnor g3147(n5644 ,n5425 ,n5192);
    nand g3148(n232 ,n165 ,n150);
    nor g3149(n1751 ,n1667 ,n1734);
    nor g3150(n1655 ,n1612 ,n1641);
    nand g3151(n4495 ,n20[3] ,n4365);
    or g3152(n2558 ,n2538 ,n2557);
    not g3153(n4412 ,n21[6]);
    nor g3154(n730 ,n611 ,n555);
    xnor g3155(n5221 ,n4899 ,n4497);
    xnor g3156(n5299 ,n4927 ,n4432);
    xnor g3157(n38[12] ,n2545 ,n2557);
    nand g3158(n5141 ,n4759 ,n4987);
    nand g3159(n472 ,n389 ,n449);
    nor g3160(n3860 ,n3679 ,n3821);
    not g3161(n5289 ,n5288);
    nand g3162(n3931 ,n3795 ,n3855);
    not g3163(n4878 ,n4877);
    nor g3164(n2741 ,n2645 ,n2713);
    not g3165(n1812 ,n1811);
    not g3166(n137 ,n136);
    xnor g3167(n2423 ,n2375 ,n2291);
    nor g3168(n2747 ,n2644 ,n2681);
    not g3169(n1562 ,n1561);
    xnor g3170(n5603 ,n5442 ,n5290);
    or g3171(n3105 ,n38[2] ,n6575);
    nand g3172(n800 ,n26[3] ,n723);
    or g3173(n3102 ,n6577 ,n6554);
    not g3174(n1194 ,n1141);
    nand g3175(n4870 ,n4469 ,n4456);
    nand g3176(n3248 ,n3195 ,n3247);
    nand g3177(n1288 ,n1042 ,n866);
    nand g3178(n4423 ,n21[7] ,n4388);
    nand g3179(n5671 ,n5453 ,n5546);
    nand g3180(n5390 ,n5201 ,n5204);
    nand g3181(n5146 ,n4796 ,n4989);
    xnor g3182(n6085 ,n6030 ,n5992);
    or g3183(n4717 ,n4568 ,n4453);
    nand g3184(n1598 ,n1570 ,n1574);
    dff g3185(.RN(n1), .SN(1'b1), .CK(n0), .D(n1280), .Q(n1500));
    nor g3186(n4778 ,n4526 ,n4666);
    xnor g3187(n692 ,n26[5] ,n22[5]);
    nand g3188(n5042 ,n4521 ,n4873);
    nand g3189(n4315 ,n4285 ,n4305);
    xnor g3190(n5155 ,n4963 ,n4435);
    xnor g3191(n6604 ,n3403 ,n3425);
    nand g3192(n1329 ,n1085 ,n928);
    or g3193(n2358 ,n2233 ,n2292);
    xnor g3194(n2241 ,n2120 ,n2128);
    nor g3195(n198 ,n177 ,n176);
    not g3196(n3894 ,n3893);
    or g3197(n4312 ,n4272 ,n4303);
    xnor g3198(n4177 ,n4109 ,n4000);
    nand g3199(n35[10] ,n6465 ,n6464);
    not g3200(n2364 ,n2351);
    or g3201(n3058 ,n3032 ,n3037);
    nand g3202(n5856 ,n5735 ,n5775);
    xnor g3203(n4208 ,n4138 ,n4115);
    xnor g3204(n6578 ,n1970 ,n2007);
    nand g3205(n4534 ,n20[0] ,n4374);
    nand g3206(n5131 ,n4753 ,n5036);
    xnor g3207(n3912 ,n3775 ,n3784);
    xnor g3208(n2865 ,n2784 ,n2735);
    nand g3209(n3116 ,n38[13] ,n6586);
    xnor g3210(n1527 ,n508 ,n518);
    nor g3211(n5377 ,n5138 ,n5282);
    nand g3212(n3382 ,n3320 ,n3381);
    dff g3213(.RN(n1), .SN(1'b1), .CK(n0), .D(n1454), .Q(n31[6]));
    xnor g3214(n6492 ,n3219 ,n3241);
    nand g3215(n1977 ,n1964 ,n1921);
    nand g3216(n913 ,n22[7] ,n719);
    nand g3217(n1233 ,n1022 ,n728);
    nand g3218(n4993 ,n4554 ,n4843);
    dff g3219(.RN(n1), .SN(1'b1), .CK(n0), .D(n1347), .Q(n23[14]));
    nor g3220(n406 ,n290 ,n368);
    nand g3221(n4652 ,n21[6] ,n4367);
    not g3222(n3262 ,n37[2]);
    nand g3223(n707 ,n562 ,n622);
    nand g3224(n3525 ,n3484 ,n19[1]);
    xor g3225(n4139 ,n4062 ,n4088);
    nand g3226(n4121 ,n4081 ,n4059);
    nand g3227(n3083 ,n3043 ,n3082);
    nand g3228(n5045 ,n4685 ,n4869);
    nand g3229(n2351 ,n2289 ,n2287);
    xnor g3230(n2916 ,n2877 ,n2729);
    xor g3231(n1532 ,n248 ,n210);
    xnor g3232(n2293 ,n2118 ,n2224);
    or g3233(n5715 ,n5640 ,n5656);
    nand g3234(n3015 ,n2942 ,n2984);
    xnor g3235(n6588 ,n1969 ,n2057);
    xnor g3236(n2238 ,n2118 ,n2129);
    nand g3237(n2201 ,n2101 ,n2173);
    nand g3238(n2336 ,n2260 ,n2314);
    nor g3239(n4122 ,n4021 ,n4090);
    not g3240(n2379 ,n2378);
    xnor g3241(n5157 ,n4942 ,n4702);
    nand g3242(n3981 ,n3849 ,n3922);
    not g3243(n2703 ,n2702);
    not g3244(n2759 ,n2758);
    nand g3245(n2159 ,n6534 ,n2127);
    not g3246(n5543 ,n5542);
    xnor g3247(n3829 ,n3569 ,n3571);
    xnor g3248(n84 ,n63 ,n45);
    nand g3249(n4288 ,n4230 ,n4274);
    nor g3250(n3352 ,n3344 ,n3351);
    xor g3251(n3952 ,n3860 ,n3873);
    xnor g3252(n1928 ,n1879 ,n1824);
    nand g3253(n1094 ,n33[6] ,n710);
    xnor g3254(n6008 ,n5911 ,n5829);
    xnor g3255(n6586 ,n2053 ,n2022);
    xnor g3256(n5198 ,n4919 ,n4588);
    nand g3257(n1129 ,n20[7] ,n722);
    nor g3258(n139 ,n132 ,n138);
    xnor g3259(n4918 ,n4629 ,n4424);
    nor g3260(n2882 ,n2766 ,n2826);
    xnor g3261(n5539 ,n5313 ,n5084);
    or g3262(n5558 ,n5172 ,n5459);
    nor g3263(n586 ,n33[1] ,n35[1]);
    not g3264(n2728 ,n2727);
    nand g3265(n2217 ,n6533 ,n2178);
    nor g3266(n415 ,n289 ,n369);
    nand g3267(n3529 ,n3478 ,n19[0]);
    xnor g3268(n2896 ,n2804 ,n2741);
    not g3269(n58 ,n36[7]);
    nor g3270(n2005 ,n1949 ,n1978);
    nand g3271(n1259 ,n843 ,n1002);
    not g3272(n1572 ,n1571);
    or g3273(n4329 ,n4320 ,n4302);
    or g3274(n4737 ,n4487 ,n4488);
    not g3275(n3474 ,n3473);
    xor g3276(n4914 ,n4522 ,n4491);
    or g3277(n5796 ,n5644 ,n5728);
    nand g3278(n4580 ,n21[1] ,n4382);
    dff g3279(.RN(n1), .SN(1'b1), .CK(n0), .D(n1307), .Q(n10[15]));
    nor g3280(n1961 ,n1867 ,n1928);
    nor g3281(n2687 ,n2565 ,n2623);
    nand g3282(n3826 ,n3568 ,n3713);
    nand g3283(n1773 ,n1666 ,n1707);
    nor g3284(n2723 ,n2568 ,n2627);
    not g3285(n560 ,n17[2]);
    nand g3286(n852 ,n1504 ,n714);
    nand g3287(n4839 ,n4457 ,n4450);
    xnor g3288(n2526 ,n2485 ,n2438);
    not g3289(n73 ,n72);
    xnor g3290(n3033 ,n2911 ,n3001);
    dff g3291(.RN(n1), .SN(1'b1), .CK(n0), .D(n1277), .Q(n16[1]));
    nand g3292(n639 ,n33[5] ,n35[5]);
    xnor g3293(n4097 ,n3971 ,n4045);
    or g3294(n6015 ,n5951 ,n5989);
    or g3295(n2579 ,n40[4] ,n6515);
    nand g3296(n6377 ,n6545 ,n6248);
    nand g3297(n3322 ,n6573 ,n6565);
    nand g3298(n701 ,n582 ,n581);
    or g3299(n5709 ,n5552 ,n5654);
    dff g3300(.RN(n1), .SN(1'b1), .CK(n0), .D(n1364), .Q(n23[7]));
    xnor g3301(n1802 ,n1745 ,n1646);
    not g3302(n2893 ,n2888);
    not g3303(n4798 ,n4430);
    or g3304(n3964 ,n3848 ,n3890);
    not g3305(n56 ,n37[1]);
    nand g3306(n4604 ,n4376 ,n20[4]);
    nor g3307(n382 ,n219 ,n343);
    not g3308(n3260 ,n37[5]);
    nor g3309(n2033 ,n1989 ,n2030);
    nand g3310(n5483 ,n5146 ,n5383);
    nand g3311(n2070 ,n20[2] ,n20[1]);
    nand g3312(n3245 ,n3205 ,n3244);
    nand g3313(n1461 ,n1130 ,n1380);
    nand g3314(n2193 ,n6536 ,n2148);
    nand g3315(n321 ,n231 ,n291);
    nand g3316(n2247 ,n2176 ,n2187);
    nand g3317(n222 ,n159 ,n146);
    not g3318(n2340 ,n2058);
    nand g3319(n4489 ,n21[0] ,n4389);
    not g3320(n4084 ,n4083);
    nand g3321(n5406 ,n5064 ,n5249);
    not g3322(n1995 ,n1994);
    nand g3323(n4571 ,n21[2] ,n4373);
    nand g3324(n1422 ,n799 ,n1177);
    nand g3325(n3324 ,n6587 ,n41[14]);
    not g3326(n4965 ,n4964);
    nor g3327(n2607 ,n2567 ,n2587);
    xor g3328(n5863 ,n5779 ,n5753);
    nor g3329(n128 ,n24[5] ,n127);
    xnor g3330(n3767 ,n3586 ,n3595);
    nand g3331(n1206 ,n815 ,n744);
    nand g3332(n4353 ,n4352 ,n4327);
    nand g3333(n5345 ,n5101 ,n5275);
    not g3334(n173 ,n36[1]);
    nand g3335(n4219 ,n4167 ,n4187);
    nand g3336(n4826 ,n4473 ,n4604);
    nand g3337(n6013 ,n5951 ,n5989);
    nand g3338(n1733 ,n1577 ,n1700);
    nor g3339(n2604 ,n2567 ,n2584);
    xor g3340(n6533 ,n3283 ,n3265);
    or g3341(n480 ,n450 ,n465);
    nand g3342(n974 ,n20[7] ,n714);
    nand g3343(n5910 ,n5740 ,n5842);
    dff g3344(.RN(n1), .SN(1'b1), .CK(n0), .D(n1216), .Q(n30[3]));
    dff g3345(.RN(n1), .SN(1'b1), .CK(n0), .D(n1217), .Q(n30[1]));
    nand g3346(n1713 ,n1582 ,n1676);
    nor g3347(n2807 ,n2669 ,n2763);
    nor g3348(n4782 ,n4652 ,n4700);
    nand g3349(n4149 ,n4067 ,n4107);
    dff g3350(.RN(n1), .SN(1'b1), .CK(n0), .D(n1394), .Q(n21[6]));
    or g3351(n3678 ,n3590 ,n3528);
    or g3352(n5272 ,n5133 ,n5071);
    not g3353(n3366 ,n3365);
    xnor g3354(n5770 ,n5607 ,n5634);
    nand g3355(n6335 ,n6491 ,n6253);
    xnor g3356(n5437 ,n5280 ,n5148);
    nand g3357(n35[13] ,n6467 ,n6484);
    not g3358(n1565 ,n37[0]);
    not g3359(n1578 ,n36[6]);
    dff g3360(.RN(n1), .SN(1'b1), .CK(n0), .D(n1326), .Q(n34[9]));
    or g3361(n2984 ,n2938 ,n2953);
    nand g3362(n3790 ,n3544 ,n3689);
    nand g3363(n3325 ,n6583 ,n6571);
    nand g3364(n4850 ,n4425 ,n4644);
    nand g3365(n6312 ,n6579 ,n6247);
    nand g3366(n6097 ,n6004 ,n6066);
    or g3367(n3056 ,n3031 ,n3035);
    dff g3368(.RN(n1), .SN(1'b1), .CK(n0), .D(n1219), .Q(n34[0]));
    or g3369(n4733 ,n4467 ,n4575);
    nand g3370(n4647 ,n21[2] ,n4374);
    xnor g3371(n1646 ,n1632 ,n1605);
    xnor g3372(n1945 ,n1884 ,n1917);
    xnor g3373(n2299 ,n2120 ,n2250);
    nand g3374(n4863 ,n4496 ,n4465);
    dff g3375(.RN(n1), .SN(1'b1), .CK(n0), .D(n1215), .Q(n30[5]));
    xnor g3376(n430 ,n376 ,n375);
    xor g3377(n3945 ,n3841 ,n3875);
    nand g3378(n413 ,n386 ,n372);
    nand g3379(n1257 ,n844 ,n1004);
    nand g3380(n1055 ,n2[0] ,n557);
    nand g3381(n3148 ,n38[3] ,n3100);
    nor g3382(n3288 ,n3275 ,n3257);
    nand g3383(n5033 ,n4698 ,n4864);
    nand g3384(n5579 ,n5333 ,n5490);
    xnor g3385(n4933 ,n4624 ,n4455);
    xnor g3386(n5200 ,n4884 ,n4638);
    nand g3387(n3521 ,n3472 ,n3478);
    or g3388(n3671 ,n3501 ,n3591);
    nand g3389(n1750 ,n1672 ,n1735);
    xnor g3390(n5598 ,n5056 ,n5462);
    nand g3391(n2069 ,n20[6] ,n20[5]);
    nor g3392(n1867 ,n1794 ,n1831);
    nand g3393(n2839 ,n2732 ,n2792);
    not g3394(n3785 ,n3784);
    xnor g3395(n1975 ,n1875 ,n1932);
    nand g3396(n4239 ,n4154 ,n4207);
    not g3397(n3900 ,n3899);
    nor g3398(n4119 ,n4044 ,n4078);
    nor g3399(n6484 ,n6422 ,n6473);
    xnor g3400(n2323 ,n2118 ,n2239);
    nor g3401(n3097 ,n6574 ,n6551);
    dff g3402(.RN(n1), .SN(1'b1), .CK(n0), .D(n1447), .Q(n12[3]));
    or g3403(n6132 ,n6029 ,n6112);
    buf g3404(n14[9], n11[9]);
    nand g3405(n5493 ,n5271 ,n5336);
    nand g3406(n1229 ,n999 ,n949);
    xnor g3407(n5455 ,n5155 ,n4787);
    nand g3408(n1451 ,n822 ,n1335);
    not g3409(n3497 ,n19[1]);
    not g3410(n4405 ,n20[6]);
    nand g3411(n1619 ,n1579 ,n1612);
    nand g3412(n6316 ,n6587 ,n6247);
    xnor g3413(n3883 ,n3743 ,n3535);
    xnor g3414(n1606 ,n1568 ,n19[5]);
    not g3415(n561 ,n17[5]);
    xnor g3416(n6158 ,n6065 ,n6127);
    nand g3417(n4272 ,n4214 ,n4255);
    not g3418(n3564 ,n3563);
    nand g3419(n5104 ,n4845 ,n4969);
    nand g3420(n5041 ,n4667 ,n4854);
    nand g3421(n1438 ,n932 ,n1212);
    nand g3422(n922 ,n30[3] ,n723);
    xnor g3423(n2321 ,n2119 ,n2255);
    xnor g3424(n1806 ,n1648 ,n1764);
    or g3425(n6199 ,n6180 ,n6187);
    dff g3426(.RN(n1), .SN(1'b1), .CK(n0), .D(n1354), .Q(n32[6]));
    nand g3427(n999 ,n12[15] ,n711);
    xor g3428(n6618 ,n6573 ,n6565);
    not g3429(n4370 ,n37[0]);
    nand g3430(n2626 ,n2590 ,n2580);
    nand g3431(n4358 ,n4288 ,n4357);
    or g3432(n1857 ,n1802 ,n1801);
    nand g3433(n282 ,n188 ,n227);
    or g3434(n3652 ,n3583 ,n3596);
    nand g3435(n3706 ,n3603 ,n3513);
    nor g3436(n4160 ,n4000 ,n4110);
    nand g3437(n1161 ,n33[15] ,n710);
    xor g3438(n6534 ,n3298 ,n3289);
    dff g3439(.RN(n1), .SN(1'b1), .CK(n0), .D(n1342), .Q(n33[10]));
    nand g3440(n3989 ,n3891 ,n3904);
    nor g3441(n2693 ,n2568 ,n2617);
    dff g3442(.RN(n1), .SN(1'b1), .CK(n0), .D(n18[0]), .Q(n15[4]));
    nand g3443(n3623 ,n3480 ,n19[0]);
    xnor g3444(n3300 ,n3279 ,n3261);
    nand g3445(n3455 ,n3449 ,n3454);
    not g3446(n3282 ,n36[0]);
    nand g3447(n6477 ,n6372 ,n6438);
    nand g3448(n3616 ,n3470 ,n3482);
    nand g3449(n952 ,n35[10] ,n712);
    nor g3450(n2506 ,n2460 ,n2476);
    nand g3451(n285 ,n223 ,n211);
    xnor g3452(n3130 ,n6581 ,n6558);
    nor g3453(n2739 ,n2567 ,n2629);
    not g3454(n3445 ,n3444);
    xnor g3455(n4092 ,n3883 ,n4023);
    xnor g3456(n6540 ,n3297 ,n3316);
    nand g3457(n1406 ,n969 ,n1162);
    nand g3458(n4608 ,n20[1] ,n4369);
    not g3459(n1584 ,n1583);
    nand g3460(n3944 ,n3790 ,n3833);
    xnor g3461(n1947 ,n1906 ,n1557);
    nand g3462(n5003 ,n4519 ,n4820);
    nand g3463(n802 ,n26[1] ,n723);
    or g3464(n2571 ,n40[6] ,n6517);
    dff g3465(.RN(n1), .SN(1'b1), .CK(n0), .D(n1235), .Q(n12[2]));
    not g3466(n2670 ,n2669);
    xnor g3467(n3751 ,n3511 ,n3604);
    nand g3468(n5736 ,n5578 ,n5613);
    not g3469(n4689 ,n4688);
    nand g3470(n4844 ,n4481 ,n4432);
    nand g3471(n1384 ,n629 ,n773);
    nand g3472(n3709 ,n3539 ,n3599);
    nor g3473(n2520 ,n2500 ,n2491);
    xnor g3474(n1817 ,n1766 ,n1648);
    nand g3475(n4589 ,n21[5] ,n4384);
    dff g3476(.RN(n1), .SN(1'b1), .CK(n0), .D(n1491), .Q(n18[2]));
    nand g3477(n1728 ,n1623 ,n1686);
    nand g3478(n5953 ,n5839 ,n5904);
    nor g3479(n6091 ,n6038 ,n6061);
    nand g3480(n2627 ,n2589 ,n2575);
    nand g3481(n1107 ,n32[7] ,n710);
    not g3482(n5527 ,n5526);
    nand g3483(n1130 ,n22[7] ,n720);
    or g3484(n4753 ,n4567 ,n4590);
    nor g3485(n2829 ,n2706 ,n2754);
    nor g3486(n76 ,n63 ,n45);
    nor g3487(n2883 ,n2798 ,n2840);
    not g3488(n4384 ,n4383);
    nand g3489(n2158 ,n6538 ,n2127);
    xnor g3490(n357 ,n335 ,n230);
    nand g3491(n5505 ,n5267 ,n5364);
    xnor g3492(n2415 ,n2371 ,n2294);
    nand g3493(n1392 ,n945 ,n1148);
    nand g3494(n1216 ,n922 ,n765);
    nor g3495(n4522 ,n4395 ,n4415);
    xnor g3496(n4066 ,n3951 ,n3850);
    or g3497(n4279 ,n4227 ,n4267);
    xnor g3498(n5228 ,n4903 ,n4454);
    or g3499(n3106 ,n6579 ,n6556);
    dff g3500(.RN(n1), .SN(1'b1), .CK(n0), .D(n1224), .Q(n27[7]));
    nand g3501(n3808 ,n3555 ,n3715);
    xor g3502(n5215 ,n4936 ,n4600);
    nand g3503(n3147 ,n38[5] ,n3104);
    nand g3504(n3573 ,n3476 ,n19[2]);
    nand g3505(n1079 ,n10[3] ,n555);
    nand g3506(n5094 ,n4876 ,n5054);
    nand g3507(n3615 ,n3486 ,n19[4]);
    xor g3508(n39[4] ,n38[4] ,n6614);
    nand g3509(n3027 ,n2994 ,n3015);
    xnor g3510(n4268 ,n4223 ,n4151);
    xnor g3511(n2859 ,n2756 ,n2704);
    nand g3512(n1111 ,n32[4] ,n710);
    nand g3513(n2226 ,n2137 ,n2184);
    xnor g3514(n2879 ,n2762 ,n2669);
    nand g3515(n4679 ,n21[6] ,n4374);
    not g3516(n3737 ,n3719);
    nand g3517(n1294 ,n873 ,n1048);
    nand g3518(n6049 ,n5909 ,n6000);
    nand g3519(n5004 ,n4524 ,n4867);
    nand g3520(n4484 ,n21[1] ,n4363);
    or g3521(n732 ,n711 ,n677);
    xnor g3522(n391 ,n346 ,n288);
    xnor g3523(n4096 ,n3944 ,n4025);
    nand g3524(n1631 ,n1598 ,n1610);
    nand g3525(n6382 ,n6489 ,n6253);
    not g3526(n67 ,n66);
    xnor g3527(n318 ,n232 ,n187);
    nand g3528(n6289 ,n6563 ,n6251);
    nor g3529(n6070 ,n6052 ,n6033);
    nand g3530(n248 ,n161 ,n157);
    nand g3531(n5071 ,n4751 ,n5001);
    nor g3532(n6260 ,n6234 ,n6252);
    nand g3533(n4199 ,n4120 ,n4161);
    nand g3534(n5148 ,n4739 ,n4984);
    nand g3535(n4463 ,n20[6] ,n4361);
    dff g3536(.RN(n1), .SN(1'b1), .CK(n0), .D(n1284), .Q(n1513));
    xnor g3537(n2441 ,n2397 ,n2399);
    nor g3538(n6261 ,n6235 ,n6252);
    or g3539(n5344 ,n5128 ,n5157);
    not g3540(n2004 ,n2003);
    xor g3541(n4902 ,n4658 ,n4568);
    nand g3542(n6181 ,n6174 ,n6163);
    not g3543(n6227 ,n25[0]);
    nand g3544(n4614 ,n21[6] ,n4388);
    nand g3545(n2184 ,n6537 ,n2150);
    not g3546(n60 ,n36[4]);
    nand g3547(n3554 ,n3486 ,n19[6]);
    nand g3548(n1224 ,n970 ,n746);
    nand g3549(n3513 ,n3460 ,n3478);
    or g3550(n4760 ,n4448 ,n4589);
    xor g3551(n6529 ,n3452 ,n3456);
    nand g3552(n4528 ,n4389 ,n20[3]);
    not g3553(n3500 ,n19[6]);
    xnor g3554(n3182 ,n3131 ,n38[12]);
    xnor g3555(n5606 ,n5443 ,n5287);
    nand g3556(n5387 ,n5200 ,n5199);
    or g3557(n95 ,n90 ,n94);
    nor g3558(n2053 ,n2052 ,n2028);
    not g3559(n1583 ,n36[1]);
    nand g3560(n6191 ,n6179 ,n6173);
    dff g3561(.RN(n1), .SN(1'b1), .CK(n0), .D(n1337), .Q(n24[4]));
    nand g3562(n3505 ,n3460 ,n3482);
    nand g3563(n6211 ,n6210 ,n6191);
    xnor g3564(n5996 ,n5908 ,n5932);
    or g3565(n5657 ,n5453 ,n5546);
    nand g3566(n439 ,n225 ,n418);
    nand g3567(n4253 ,n4200 ,n4241);
    nand g3568(n5355 ,n5149 ,n5272);
    xor g3569(n4925 ,n4649 ,n4609);
    nor g3570(n716 ,n18[2] ,n621);
    nand g3571(n5271 ,n5079 ,n5119);
    or g3572(n4758 ,n4616 ,n4472);
    nor g3573(n2462 ,n2395 ,n2436);
    nand g3574(n3926 ,n3684 ,n3844);
    nand g3575(n1226 ,n979 ,n790);
    xnor g3576(n5218 ,n4889 ,n4614);
    xor g3577(n5779 ,n5602 ,n5493);
    nand g3578(n1228 ,n985 ,n788);
    nand g3579(n4830 ,n4602 ,n4587);
    xnor g3580(n4949 ,n4585 ,n4608);
    nand g3581(n3646 ,n3484 ,n19[0]);
    nand g3582(n493 ,n429 ,n462);
    nor g3583(n2275 ,n2229 ,n2232);
    nor g3584(n4978 ,n4435 ,n4788);
    xor g3585(n4884 ,n4661 ,n4576);
    xnor g3586(n682 ,n35[6] ,n33[6]);
    nand g3587(n341 ,n271 ,n326);
    nand g3588(n4806 ,n4442 ,n4459);
    nand g3589(n246 ,n167 ,n153);
    not g3590(n6094 ,n6093);
    nand g3591(n1439 ,n933 ,n1213);
    nand g3592(n3811 ,n3632 ,n3718);
    xnor g3593(n3022 ,n2973 ,n2956);
    xnor g3594(n6589 ,n3253 ,n3211);
    nor g3595(n1552 ,n128 ,n130);
    nand g3596(n1404 ,n654 ,n783);
    xnor g3597(n3169 ,n3128 ,n38[5]);
    not g3598(n2851 ,n2850);
    nand g3599(n3354 ,n6577 ,n3353);
    nand g3600(n6228 ,n6226 ,n6225);
    nand g3601(n195 ,n161 ,n152);
    or g3602(n1979 ,n1956 ,n1923);
    or g3603(n412 ,n382 ,n374);
    xnor g3604(n4974 ,n4632 ,n4480);
    xor g3605(n6515 ,n6554 ,n6577);
    nand g3606(n1282 ,n861 ,n1034);
    nand g3607(n1298 ,n1054 ,n804);
    xnor g3608(n1757 ,n1636 ,n1679);
    nand g3609(n5563 ,n5393 ,n5461);
    nor g3610(n2688 ,n2565 ,n2630);
    xnor g3611(n2273 ,n2108 ,n2208);
    nand g3612(n5677 ,n5576 ,n5579);
    nor g3613(n6482 ,n6439 ,n6477);
    xnor g3614(n41[4] ,n6084 ,n6016);
    nand g3615(n1275 ,n639 ,n729);
    not g3616(n563 ,n18[2]);
    nor g3617(n2409 ,n2339 ,n2390);
    xnor g3618(n5288 ,n4946 ,n4442);
    xnor g3619(n5639 ,n5435 ,n5129);
    nand g3620(n2072 ,n20[0] ,n21[0]);
    nand g3621(n3856 ,n3531 ,n3781);
    nand g3622(n1795 ,n1648 ,n1753);
    nand g3623(n3563 ,n3484 ,n19[6]);
    or g3624(n5887 ,n5780 ,n5832);
    nand g3625(n633 ,n33[8] ,n35[8]);
    nand g3626(n1307 ,n1065 ,n953);
    nand g3627(n4852 ,n4607 ,n4643);
    nand g3628(n6017 ,n5940 ,n5980);
    nand g3629(n1077 ,n27[13] ,n718);
    not g3630(n1927 ,n1926);
    nor g3631(n587 ,n34[0] ,n34[12]);
    not g3632(n555 ,n712);
    nand g3633(n6426 ,n6290 ,n6357);
    nand g3634(n190 ,n165 ,n146);
    xnor g3635(n1994 ,n1904 ,n1944);
    buf g3636(n13[6], n11[6]);
    nand g3637(n4338 ,n4316 ,n4325);
    nor g3638(n6460 ,n6420 ,n6419);
    dff g3639(.RN(n1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n23[10]));
    nor g3640(n2306 ,n2152 ,n2266);
    or g3641(n885 ,n555 ,n673);
    or g3642(n446 ,n388 ,n430);
    nand g3643(n2027 ,n2020 ,n1993);
    nand g3644(n5152 ,n4721 ,n5027);
    nand g3645(n4318 ,n4293 ,n4306);
    nand g3646(n1081 ,n27[9] ,n718);
    xnor g3647(n5724 ,n5509 ,n5590);
    nand g3648(n6000 ,n5873 ,n5973);
    nor g3649(n4694 ,n4415 ,n4407);
    nand g3650(n889 ,n33[6] ,n712);
    xnor g3651(n3002 ,n2970 ,n2914);
    or g3652(n4705 ,n4564 ,n4485);
    nand g3653(n6299 ,n41[4] ,n6254);
    nand g3654(n492 ,n403 ,n474);
    nand g3655(n3597 ,n3460 ,n3486);
    nor g3656(n3617 ,n3491 ,n3495);
    nand g3657(n6378 ,n6510 ,n6249);
    nand g3658(n1898 ,n1558 ,n1854);
    nand g3659(n6401 ,n6277 ,n6326);
    nand g3660(n1446 ,n1024 ,n1275);
    nor g3661(n734 ,n586 ,n555);
    xnor g3662(n6057 ,n5931 ,n6019);
    not g3663(n5635 ,n5634);
    xnor g3664(n5211 ,n4926 ,n4562);
    nand g3665(n6432 ,n6293 ,n6364);
    nand g3666(n3729 ,n3579 ,n3527);
    nand g3667(n1390 ,n1091 ,n957);
    not g3668(n564 ,n34[7]);
    nand g3669(n6395 ,n6271 ,n6323);
    nand g3670(n6435 ,n6299 ,n6369);
    nor g3671(n2961 ,n2940 ,n2939);
    or g3672(n759 ,n720 ,n698);
    nor g3673(n2496 ,n2406 ,n2473);
    or g3674(n1935 ,n1903 ,n1905);
    xnor g3675(n4176 ,n4069 ,n4111);
    nand g3676(n1762 ,n1664 ,n1719);
    nor g3677(n2833 ,n2707 ,n2753);
    xnor g3678(n3333 ,n41[12] ,n6585);
    nand g3679(n6476 ,n6380 ,n6430);
    nand g3680(n1011 ,n3[7] ,n713);
    nand g3681(n5650 ,n5547 ,n5523);
    nor g3682(n2699 ,n2565 ,n2619);
    nand g3683(n3246 ,n3192 ,n3245);
    nor g3684(n2555 ,n2539 ,n2554);
    nand g3685(n814 ,n34[5] ,n717);
    nand g3686(n881 ,n1549 ,n712);
    nand g3687(n856 ,n1501 ,n714);
    not g3688(n164 ,n36[6]);
    nand g3689(n2596 ,n40[13] ,n6524);
    xnor g3690(n6177 ,n6121 ,n6145);
    nand g3691(n6041 ,n5991 ,n6003);
    not g3692(n2363 ,n2346);
    not g3693(n63 ,n62);
    nor g3694(n2608 ,n2567 ,n2594);
    nand g3695(n6318 ,n40[8] ,n6250);
    nand g3696(n3711 ,n3512 ,n3536);
    nand g3697(n3810 ,n3558 ,n3717);
    or g3698(n4715 ,n4614 ,n4444);
    nand g3699(n4191 ,n4079 ,n4153);
    nand g3700(n3839 ,n3685 ,n3783);
    nand g3701(n4073 ,n3900 ,n4022);
    nand g3702(n1770 ,n1695 ,n1709);
    nor g3703(n742 ,n660 ,n717);
    nand g3704(n3385 ,n3336 ,n3384);
    xnor g3705(n4055 ,n3946 ,n3890);
    xnor g3706(n2921 ,n2862 ,n2892);
    xor g3707(n40[10] ,n6601 ,n38[11]);
    nor g3708(n4227 ,n4144 ,n4204);
    xnor g3709(n2925 ,n2876 ,n2768);
    nand g3710(n6341 ,n6488 ,n6253);
    nand g3711(n1462 ,n923 ,n1381);
    nand g3712(n1518 ,n439 ,n553);
    nand g3713(n5076 ,n4711 ,n5014);
    dff g3714(.RN(n1), .SN(1'b1), .CK(n0), .D(n1399), .Q(n21[4]));
    nor g3715(n2718 ,n2566 ,n2620);
    not g3716(n142 ,n141);
    nand g3717(n408 ,n308 ,n370);
    nand g3718(n2480 ,n2423 ,n2447);
    nand g3719(n2174 ,n6540 ,n2126);
    not g3720(n2952 ,n2951);
    nand g3721(n4246 ,n4191 ,n4213);
    xnor g3722(n6611 ,n3329 ,n3368);
    not g3723(n5352 ,n5351);
    xnor g3724(n3331 ,n6572 ,n6584);
    xnor g3725(n2398 ,n2326 ,n2320);
    not g3726(n1847 ,n1557);
    xor g3727(n4888 ,n4505 ,n4636);
    nand g3728(n5103 ,n4830 ,n4965);
    xnor g3729(n6605 ,n3414 ,n3423);
    nand g3730(n1088 ,n1552 ,n716);
    nand g3731(n5814 ,n5676 ,n5743);
    xnor g3732(n6564 ,n4298 ,n4356);
    nand g3733(n5259 ,n5081 ,n5125);
    nand g3734(n136 ,n32[2] ,n135);
    xnor g3735(n5830 ,n5698 ,n5640);
    nand g3736(n4189 ,n4172 ,n4146);
    not g3737(n5541 ,n5540);
    nand g3738(n4823 ,n4605 ,n4599);
    or g3739(n5515 ,n5498 ,n5496);
    nand g3740(n5364 ,n5144 ,n5241);
    nand g3741(n221 ,n170 ,n152);
    xnor g3742(n5535 ,n5307 ,n5090);
    nand g3743(n3607 ,n3466 ,n3484);
    or g3744(n4120 ,n4025 ,n4057);
    nor g3745(n3390 ,n6560 ,n6545);
    not g3746(n559 ,n18[1]);
    nand g3747(n4126 ,n3939 ,n4063);
    xnor g3748(n2440 ,n2393 ,n2327);
    not g3749(n5409 ,n5387);
    not g3750(n5132 ,n5131);
    nor g3751(n2540 ,n2502 ,n2526);
    nand g3752(n5990 ,n5893 ,n5946);
    nand g3753(n1754 ,n1659 ,n1739);
    xnor g3754(n5997 ,n5879 ,n5953);
    nand g3755(n5347 ,n5115 ,n5175);
    xor g3756(n40[5] ,n38[6] ,n6606);
    or g3757(n5901 ,n5779 ,n5830);
    nand g3758(n2223 ,n2134 ,n2180);
    nand g3759(n4585 ,n20[0] ,n4373);
    nand g3760(n4996 ,n4696 ,n4816);
    nand g3761(n4460 ,n21[1] ,n4367);
    nor g3762(n3858 ,n3695 ,n3799);
    nand g3763(n4856 ,n4491 ,n4482);
    not g3764(n3632 ,n3631);
    or g3765(n4757 ,n4501 ,n4573);
    nand g3766(n3142 ,n38[6] ,n3106);
    xnor g3767(n2489 ,n2443 ,n2427);
    nand g3768(n6194 ,n6172 ,n6181);
    nand g3769(n1351 ,n642 ,n751);
    nand g3770(n2585 ,n40[1] ,n6512);
    not g3771(n3136 ,n3135);
    nand g3772(n3113 ,n38[10] ,n6560);
    nand g3773(n6412 ,n6239 ,n6258);
    xnor g3774(n3303 ,n3277 ,n3267);
    nand g3775(n5002 ,n4561 ,n4819);
    nand g3776(n279 ,n186 ,n216);
    nand g3777(n1449 ,n813 ,n1330);
    xor g3778(n428 ,n355 ,n366);
    nand g3779(n3547 ,n3466 ,n3482);
    nand g3780(n1039 ,n2[5] ,n557);
    xnor g3781(n4094 ,n3899 ,n4022);
    xnor g3782(n2448 ,n2284 ,n2413);
    xnor g3783(n2466 ,n2424 ,n2400);
    xnor g3784(n5826 ,n5699 ,n5531);
    not g3785(n2362 ,n2344);
    nand g3786(n2511 ,n2483 ,n2489);
    nand g3787(n2197 ,n6539 ,n2150);
    nor g3788(n4506 ,n4400 ,n4413);
    xnor g3789(n1551 ,n24[6] ,n129);
    nand g3790(n1772 ,n1692 ,n1737);
    nand g3791(n1069 ,n10[11] ,n711);
    nand g3792(n5565 ,n5494 ,n5499);
    nand g3793(n1454 ,n1117 ,n1365);
    nand g3794(n1141 ,n20[4] ,n722);
    not g3795(n4377 ,n36[4]);
    xnor g3796(n3954 ,n3829 ,n3867);
    or g3797(n3663 ,n3538 ,n3505);
    nand g3798(n2249 ,n2171 ,n2220);
    xor g3799(n4936 ,n4657 ,n4641);
    nor g3800(n604 ,n22[1] ,n26[1]);
    nand g3801(n5734 ,n5571 ,n5688);
    or g3802(n1516 ,n32[6] ,n119);
    xnor g3803(n1529 ,n460 ,n457);
    nand g3804(n6374 ,n39[5] ,n6248);
    nand g3805(n1668 ,n1579 ,n1651);
    nor g3806(n2831 ,n2734 ,n2778);
    xnor g3807(n2971 ,n2943 ,n2925);
    nand g3808(n141 ,n32[5] ,n139);
    nand g3809(n4448 ,n21[1] ,n4376);
    xnor g3810(n5287 ,n4951 ,n4691);
    or g3811(n3418 ,n3408 ,n3417);
    nand g3812(n1896 ,n1790 ,n1845);
    nand g3813(n893 ,n23[10] ,n715);
    nand g3814(n6349 ,n6497 ,n6249);
    xnor g3815(n5623 ,n5427 ,n5185);
    xnor g3816(n6554 ,n4251 ,n4220);
    nand g3817(n6358 ,n38[10] ,n6246);
    nand g3818(n3720 ,n3532 ,n3529);
    dff g3819(.RN(n1), .SN(1'b1), .CK(n0), .D(n1271), .Q(n16[3]));
    xnor g3820(n2530 ,n2482 ,n2489);
    nand g3821(n211 ,n169 ,n152);
    nand g3822(n3077 ,n3054 ,n3076);
    nand g3823(n275 ,n180 ,n222);
    nand g3824(n1416 ,n987 ,n1175);
    dff g3825(.RN(n1), .SN(1'b1), .CK(n0), .D(n1310), .Q(n10[12]));
    nor g3826(n2600 ,n2567 ,n2595);
    or g3827(n4164 ,n4086 ,n4119);
    nand g3828(n3795 ,n3605 ,n3691);
    nand g3829(n118 ,n32[5] ,n117);
    nand g3830(n2222 ,n2156 ,n2216);
    xnor g3831(n3405 ,n39[2] ,n6551);
    nand g3832(n1680 ,n1586 ,n1654);
    nand g3833(n4494 ,n21[4] ,n4382);
    not g3834(n2311 ,n2310);
    nand g3835(n483 ,n470 ,n467);
    not g3836(n2922 ,n2921);
    xnor g3837(n3123 ,n6576 ,n6553);
    nand g3838(n902 ,n23[14] ,n715);
    nand g3839(n6359 ,n6498 ,n6249);
    xnor g3840(n4968 ,n4697 ,n4651);
    nand g3841(n1057 ,n11[5] ,n711);
    nor g3842(n3669 ,n3598 ,n3593);
    nand g3843(n4814 ,n4562 ,n4591);
    xnor g3844(n3329 ,n41[7] ,n6580);
    or g3845(n4749 ,n4437 ,n4596);
    xnor g3846(n5172 ,n4911 ,n4645);
    xnor g3847(n1805 ,n1760 ,n1646);
    xnor g3848(n3453 ,n3443 ,n19[1]);
    nand g3849(n5348 ,n5099 ,n5273);
    or g3850(n703 ,n22[1] ,n577);
    nor g3851(n724 ,n18[0] ,n663);
    nand g3852(n626 ,n17[4] ,n26[4]);
    nand g3853(n1427 ,n802 ,n1183);
    not g3854(n3343 ,n3342);
    xnor g3855(n1528 ,n496 ,n494);
    nand g3856(n3144 ,n38[4] ,n3102);
    not g3857(n240 ,n239);
    nor g3858(n2691 ,n2566 ,n2621);
    nand g3859(n1942 ,n1883 ,n1903);
    nand g3860(n4320 ,n4283 ,n4307);
    nand g3861(n1116 ,n1526 ,n716);
    xnor g3862(n2871 ,n2779 ,n2672);
    nand g3863(n4560 ,n21[3] ,n4369);
    nor g3864(n2681 ,n2568 ,n2623);
    xnor g3865(n2023 ,n1985 ,n1996);
    xnor g3866(n6160 ,n6105 ,n6138);
    dff g3867(.RN(n1), .SN(1'b1), .CK(n0), .D(n1327), .Q(n10[3]));
    nand g3868(n516 ,n480 ,n501);
    nand g3869(n355 ,n251 ,n323);
    nand g3870(n6157 ,n6097 ,n6135);
    nand g3871(n6168 ,n6150 ,n6157);
    xnor g3872(n2292 ,n2248 ,n2120);
    xnor g3873(n4924 ,n4611 ,n4597);
    nor g3874(n2820 ,n2672 ,n2780);
    nand g3875(n1441 ,n1006 ,n1260);
    nand g3876(n6399 ,n6276 ,n6325);
    nand g3877(n4630 ,n20[5] ,n4361);
    nand g3878(n5378 ,n5138 ,n5282);
    not g3879(n5592 ,n5554);
    nand g3880(n5263 ,n5108 ,n5085);
    or g3881(n4751 ,n4581 ,n4586);
    nand g3882(n6357 ,n39[3] ,n6248);
    nand g3883(n630 ,n22[0] ,n26[0]);
    nand g3884(n443 ,n380 ,n395);
    nand g3885(n1403 ,n1161 ,n953);
    nor g3886(n5713 ,n5540 ,n5629);
    not g3887(n372 ,n371);
    xnor g3888(n477 ,n451 ,n459);
    xnor g3889(n38[7] ,n2530 ,n2546);
    nand g3890(n3115 ,n6580 ,n6557);
    or g3891(n4145 ,n4070 ,n4101);
    nand g3892(n6308 ,n40[11] ,n6250);
    nor g3893(n4674 ,n4392 ,n4402);
    nand g3894(n6062 ,n5966 ,n6031);
    or g3895(n255 ,n190 ,n181);
    not g3896(n2418 ,n2417);
    xnor g3897(n5836 ,n5692 ,n5508);
    nand g3898(n930 ,n29[4] ,n721);
    not g3899(n1925 ,n1924);
    not g3900(n4390 ,n37[1]);
    xnor g3901(n5696 ,n5544 ,n5517);
    nor g3902(n291 ,n247 ,n200);
    nor g3903(n3425 ,n3395 ,n3424);
    nand g3904(n5384 ,n5187 ,n5186);
    nor g3905(n2276 ,n2231 ,n2230);
    nand g3906(n442 ,n379 ,n412);
    xnor g3907(n2086 ,n20[5] ,n21[5]);
    nor g3908(n1593 ,n1560 ,n19[7]);
    or g3909(n2431 ,n2391 ,n2396);
    or g3910(n6043 ,n5972 ,n6002);
    xnor g3911(n5869 ,n5767 ,n5815);
    not g3912(n6225 ,n25[1]);
    nor g3913(n2790 ,n2639 ,n2698);
    nand g3914(n932 ,n29[2] ,n721);
    nand g3915(n4076 ,n4002 ,n4018);
    nand g3916(n5492 ,n5265 ,n5325);
    xnor g3917(n709 ,n23[0] ,n16[0]);
    nand g3918(n187 ,n159 ,n148);
    nand g3919(n1383 ,n657 ,n769);
    nand g3920(n1119 ,n1529 ,n716);
    nor g3921(n2610 ,n2567 ,n2582);
    nand g3922(n1984 ,n1942 ,n1957);
    nand g3923(n4196 ,n4102 ,n4162);
    nand g3924(n4835 ,n4611 ,n4597);
    xnor g3925(n3070 ,n3035 ,n3031);
    not g3926(n3272 ,n36[4]);
    not g3927(n1974 ,n1973);
    xnor g3928(n5156 ,n4916 ,n4968);
    nand g3929(n5935 ,n5778 ,n5872);
    or g3930(n3387 ,n6551 ,n39[2]);
    nand g3931(n3535 ,n3486 ,n19[0]);
    not g3932(n2780 ,n2779);
    nand g3933(n410 ,n362 ,n373);
    xnor g3934(n5772 ,n5603 ,n5636);
    nand g3935(n326 ,n205 ,n285);
    nand g3936(n3203 ,n3161 ,n3174);
    xnor g3937(n3020 ,n2982 ,n2983);
    nand g3938(n1038 ,n11[15] ,n710);
    or g3939(n5732 ,n5592 ,n5642);
    nand g3940(n5689 ,n5376 ,n5563);
    xnor g3941(n3127 ,n6579 ,n6556);
    nand g3942(n2254 ,n2168 ,n2193);
    xnor g3943(n4881 ,n4492 ,n4434);
    nand g3944(n5258 ,n5069 ,n5075);
    nand g3945(n839 ,n25[0] ,n714);
    or g3946(n5238 ,n5137 ,n5126);
    not g3947(n3470 ,n3469);
    nand g3948(n4071 ,n4043 ,n3972);
    dff g3949(.RN(n1), .SN(1'b1), .CK(n0), .D(n1300), .Q(n11[6]));
    nand g3950(n1095 ,n1518 ,n716);
    not g3951(n3334 ,n3333);
    dff g3952(.RN(n1), .SN(1'b1), .CK(n0), .D(n1287), .Q(n11[14]));
    not g3953(n3848 ,n3847);
    nand g3954(n3508 ,n3466 ,n3476);
    nand g3955(n5499 ,n5257 ,n5340);
    xnor g3956(n6112 ,n6055 ,n6036);
    nand g3957(n1220 ,n938 ,n753);
    nand g3958(n4256 ,n4197 ,n4239);
    nand g3959(n1002 ,n4[2] ,n713);
    xnor g3960(n6109 ,n6004 ,n6066);
    or g3961(n5899 ,n5823 ,n5852);
    or g3962(n5481 ,n5293 ,n5377);
    xnor g3963(n82 ,n61 ,n47);
    nand g3964(n6151 ,n6138 ,n6105);
    xnor g3965(n5424 ,n5170 ,n5171);
    xnor g3966(n5859 ,n5784 ,n5805);
    not g3967(n3478 ,n3477);
    xnor g3968(n1554 ,n24[3] ,n124);
    not g3969(n83 ,n82);
    xnor g3970(n3372 ,n6581 ,n3370);
    nor g3971(n2758 ,n2643 ,n2685);
    nand g3972(n1486 ,n791 ,n1434);
    xnor g3973(n5638 ,n5431 ,n5139);
    nand g3974(n5948 ,n5813 ,n5899);
    not g3975(n4542 ,n4541);
    nand g3976(n6398 ,n6341 ,n6340);
    nor g3977(n2359 ,n2306 ,n2320);
    nand g3978(n2154 ,n6541 ,n2127);
    nand g3979(n4574 ,n21[3] ,n4382);
    nor g3980(n2827 ,n2708 ,n2802);
    nand g3981(n3205 ,n3162 ,n3175);
    nand g3982(n1893 ,n1784 ,n1863);
    or g3983(n2848 ,n2744 ,n2772);
    nand g3984(n2453 ,n2412 ,n2431);
    nor g3985(n2742 ,n2605 ,n2680);
    nand g3986(n1683 ,n1588 ,n1655);
    nand g3987(n1659 ,n1579 ,n1649);
    or g3988(n5327 ,n5208 ,n5207);
    nor g3989(n2214 ,n2061 ,n2177);
    nand g3990(n6350 ,n6506 ,n6249);
    dff g3991(.RN(n1), .SN(1'b1), .CK(n0), .D(n1254), .Q(n19[4]));
    not g3992(n4374 ,n4390);
    nand g3993(n3542 ,n3481 ,n19[3]);
    nand g3994(n5717 ,n5641 ,n5658);
    not g3995(n4365 ,n4364);
    xnor g3996(n1537 ,n100 ,n88);
    xnor g3997(n5292 ,n4950 ,n4440);
    nand g3998(n4843 ,n4569 ,n4601);
    not g3999(n1575 ,n36[7]);
    dff g4000(.RN(n1), .SN(1'b1), .CK(n0), .D(n1338), .Q(n33[14]));
    xnor g4001(n1543 ,n32[7] ,n143);
    xnor g4002(n5308 ,n5100 ,n5135);
    or g4003(n6189 ,n6179 ,n6173);
    nand g4004(n6268 ,n40[7] ,n6250);
    xnor g4005(n3941 ,n3767 ,n3629);
    xnor g4006(n3068 ,n3038 ,n3029);
    xnor g4007(n5219 ,n4896 ,n4642);
    nor g4008(n2756 ,n2599 ,n2679);
    nand g4009(n241 ,n172 ,n148);
    buf g4010(n15[7], 1'b0);
    xnor g4011(n2269 ,n2108 ,n2200);
    nand g4012(n3549 ,n3480 ,n19[7]);
    nand g4013(n343 ,n258 ,n331);
    nand g4014(n956 ,n35[14] ,n712);
    xor g4015(n6514 ,n6576 ,n6553);
    or g4016(n4746 ,n4496 ,n4465);
    xnor g4017(n6055 ,n5990 ,n6020);
    nor g4018(n3976 ,n3866 ,n3885);
    nor g4019(n105 ,n85 ,n104);
    xor g4020(n38[1] ,n2271 ,n2153);
    or g4021(n3187 ,n3157 ,n3172);
    not g4022(n146 ,n145);
    nand g4023(n1097 ,n33[5] ,n555);
    xnor g4024(n299 ,n192 ,n226);
    xnor g4025(n1803 ,n1773 ,n1646);
    nand g4026(n4556 ,n21[3] ,n4374);
    xnor g4027(n2545 ,n2521 ,n2533);
    nand g4028(n2256 ,n2169 ,n2190);
    not g4029(n1586 ,n1585);
    xnor g4030(n6559 ,n4342 ,n4346);
    xnor g4031(n4326 ,n4297 ,n4287);
    nand g4032(n4866 ,n4623 ,n4592);
    or g4033(n6133 ,n6103 ,n6114);
    nand g4034(n1843 ,n1774 ,n1823);
    not g4035(n3783 ,n3782);
    nor g4036(n3667 ,n3584 ,n3547);
    nand g4037(n2943 ,n2805 ,n2908);
    nor g4038(n2821 ,n2660 ,n2746);
    nand g4039(n2888 ,n2852 ,n2843);
    nand g4040(n4817 ,n4461 ,n4594);
    nand g4041(n5472 ,n5295 ,n5385);
    nand g4042(n1386 ,n627 ,n776);
    xor g4043(n4913 ,n4515 ,n4443);
    nand g4044(n1330 ,n636 ,n757);
    dff g4045(.RN(n1), .SN(1'b1), .CK(n0), .D(n1426), .Q(n19[7]));
    nand g4046(n3156 ,n3114 ,n3150);
    xnor g4047(n5312 ,n5074 ,n5101);
    xnor g4048(n3349 ,n6575 ,n3347);
    nand g4049(n1308 ,n1066 ,n956);
    dff g4050(.RN(n1), .SN(1'b1), .CK(n0), .D(n1429), .Q(n19[5]));
    xnor g4051(n2417 ,n2365 ,n2285);
    xnor g4052(n4892 ,n4577 ,n4449);
    nand g4053(n339 ,n269 ,n310);
    nand g4054(n6039 ,n5972 ,n6002);
    or g4055(n4731 ,n4580 ,n4499);
    dff g4056(.RN(n1), .SN(1'b1), .CK(n0), .D(n1411), .Q(n20[6]));
    not g4057(n3323 ,n3322);
    nand g4058(n1256 ,n841 ,n1073);
    nand g4059(n6360 ,n6490 ,n6253);
    nand g4060(n6080 ,n6010 ,n6049);
    not g4061(n5456 ,n5455);
    nand g4062(n1152 ,n6[5] ,n713);
    xnor g4063(n6616 ,n3349 ,n6567);
    not g4064(n163 ,n162);
    xnor g4065(n2955 ,n2872 ,n2909);
    nand g4066(n1313 ,n1071 ,n951);
    nand g4067(n652 ,n20[2] ,n28[2]);
    or g4068(n3100 ,n6576 ,n6553);
    nor g4069(n1866 ,n1818 ,n1799);
    xnor g4070(n6510 ,n3091 ,n3066);
    nand g4071(n1087 ,n1551 ,n716);
    xnor g4072(n3052 ,n3007 ,n3025);
    dff g4073(.RN(n1), .SN(1'b1), .CK(n0), .D(n1234), .Q(n12[4]));
    nor g4074(n104 ,n76 ,n103);
    nor g4075(n1989 ,n1912 ,n1976);
    nand g4076(n6213 ,n6212 ,n6199);
    nand g4077(n468 ,n417 ,n448);
    nor g4078(n2461 ,n2398 ,n2419);
    xnor g4079(n6614 ,n3355 ,n41[4]);
    dff g4080(.RN(n1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n23[13]));
    xnor g4081(n5416 ,n5156 ,n5198);
    not g4082(n1561 ,n37[6]);
    xnor g4083(n5975 ,n5862 ,n5833);
    nand g4084(n2517 ,n2481 ,n2495);
    nand g4085(n6418 ,n6284 ,n6345);
    xnor g4086(n4111 ,n4016 ,n3942);
    not g4087(n2484 ,n2480);
    xnor g4088(n512 ,n476 ,n462);
    nor g4089(n884 ,n571 ,n720);
    dff g4090(.RN(n1), .SN(1'b1), .CK(n0), .D(n1261), .Q(n19[1]));
    nand g4091(n3585 ,n3468 ,n3478);
    nand g4092(n6419 ,n6298 ,n6347);
    nand g4093(n6245 ,n41[7] ,n6593);
    nand g4094(n1105 ,n1522 ,n716);
    nor g4095(n4672 ,n4398 ,n4396);
    or g4096(n5245 ,n5110 ,n5135);
    nand g4097(n6429 ,n6241 ,n6259);
    xnor g4098(n5602 ,n5404 ,n5503);
    or g4099(n782 ,n711 ,n685);
    nand g4100(n1163 ,n1555 ,n716);
    nand g4101(n655 ,n16[6] ,n23[6]);
    xnor g4102(n4151 ,n4052 ,n4089);
    nand g4103(n3929 ,n3863 ,n3861);
    nand g4104(n3501 ,n3464 ,n3484);
    nor g4105(n6466 ,n6435 ,n6433);
    or g4106(n1865 ,n1701 ,n1820);
    nand g4107(n5360 ,n5102 ,n5236);
    nor g4108(n1937 ,n1786 ,n1910);
    nor g4109(n2433 ,n2276 ,n2402);
    nor g4110(n662 ,n563 ,n18[1]);
    or g4111(n3919 ,n3684 ,n3844);
    xnor g4112(n2535 ,n2490 ,n2514);
    xor g4113(n40[1] ,n6610 ,n38[2]);
    nand g4114(n4434 ,n21[0] ,n4365);
    nor g4115(n2884 ,n2770 ,n2821);
    xnor g4116(n2938 ,n2875 ,n2767);
    xnor g4117(n6027 ,n5955 ,n5995);
    nand g4118(n978 ,n20[5] ,n714);
    or g4119(n792 ,n652 ,n721);
    nand g4120(n1447 ,n1030 ,n1278);
    xnor g4121(n3335 ,n41[14] ,n6587);
    xnor g4122(n3134 ,n6561 ,n6584);
    nand g4123(n6136 ,n6123 ,n6111);
    or g4124(n5986 ,n5879 ,n5930);
    xnor g4125(n5964 ,n5871 ,n5799);
    nor g4126(n2677 ,n2566 ,n2628);
    nand g4127(n4549 ,n21[0] ,n4386);
    nor g4128(n3432 ,n3412 ,n3431);
    dff g4129(.RN(n1), .SN(1'b1), .CK(n0), .D(n1291), .Q(n11[11]));
    nand g4130(n803 ,n26[0] ,n723);
    nor g4131(n2931 ,n2809 ,n2902);
    nand g4132(n386 ,n257 ,n348);
    nand g4133(n6217 ,n6216 ,n6202);
    nand g4134(n525 ,n507 ,n512);
    nand g4135(n5667 ,n5351 ,n5520);
    nand g4136(n1270 ,n850 ,n1016);
    xor g4137(n4897 ,n4694 ,n4581);
    xor g4138(n39[1] ,n6617 ,n38[1]);
    xnor g4139(n4939 ,n4610 ,n4598);
    not g4140(n1953 ,n1952);
    nand g4141(n1181 ,n4[7] ,n557);
    xnor g4142(n3067 ,n3039 ,n3028);
    or g4143(n4773 ,n4577 ,n4449);
    nand g4144(n3589 ,n3464 ,n3486);
    nor g4145(n6149 ,n6130 ,n6094);
    xnor g4146(n691 ,n562 ,n26[1]);
    nand g4147(n1065 ,n10[15] ,n711);
    nand g4148(n2082 ,n21[6] ,n2067);
    xnor g4149(n1603 ,n19[3] ,n19[4]);
    nand g4150(n4047 ,n3926 ,n3961);
    nand g4151(n4873 ,n4566 ,n4476);
    nand g4152(n894 ,n28[0] ,n717);
    xnor g4153(n5819 ,n5620 ,n5722);
    nor g4154(n2792 ,n2654 ,n2718);
    or g4155(n5339 ,n5284 ,n5287);
    xnor g4156(n3342 ,n6571 ,n6583);
    nand g4157(n5503 ,n5255 ,n5375);
    nand g4158(n4628 ,n21[2] ,n4376);
    nand g4159(n6274 ,n6558 ,n6251);
    xnor g4160(n6569 ,n6186 ,n6201);
    xnor g4161(n3741 ,n3539 ,n3599);
    xnor g4162(n2291 ,n2247 ,n2118);
    dff g4163(.RN(n1), .SN(1'b1), .CK(n0), .D(n1294), .Q(n1510));
    not g4164(n4410 ,n4384);
    not g4165(n4367 ,n4366);
    nand g4166(n6291 ,n6553 ,n6251);
    nand g4167(n1693 ,n1579 ,n1654);
    xnor g4168(n3972 ,n3745 ,n3851);
    not g4169(n4397 ,n20[5]);
    nor g4170(n4032 ,n3911 ,n4003);
    or g4171(n5463 ,n5227 ,n5410);
    nand g4172(n1024 ,n12[5] ,n710);
    nor g4173(n605 ,n17[6] ,n26[6]);
    xnor g4174(n5315 ,n5117 ,n5088);
    not g4175(n51 ,n50);
    or g4176(n4777 ,n4460 ,n4571);
    nor g4177(n2656 ,n2565 ,n2591);
    nor g4178(n2482 ,n2342 ,n2458);
    nand g4179(n3089 ,n3042 ,n3088);
    or g4180(n3186 ,n3153 ,n3170);
    nand g4181(n3966 ,n3850 ,n3920);
    nand g4182(n6121 ,n6075 ,n6104);
    buf g4183(n13[11], n10[11]);
    nand g4184(n2622 ,n2586 ,n2570);
    nand g4185(n1114 ,n1525 ,n716);
    nand g4186(n827 ,n17[3] ,n721);
    nor g4187(n2686 ,n2565 ,n2620);
    nand g4188(n4592 ,n21[4] ,n4369);
    nand g4189(n5896 ,n5780 ,n5832);
    nor g4190(n2380 ,n2300 ,n2330);
    nor g4191(n2472 ,n2451 ,n2417);
    nand g4192(n323 ,n245 ,n287);
    or g4193(n778 ,n717 ,n679);
    nand g4194(n2138 ,n6537 ,n2122);
    xnor g4195(n4022 ,n3882 ,n3687);
    xnor g4196(n476 ,n429 ,n456);
    nand g4197(n2334 ,n2119 ,n2294);
    nor g4198(n3992 ,n3794 ,n3910);
    nand g4199(n1165 ,n5[7] ,n713);
    nand g4200(n5754 ,n5561 ,n5679);
    nor g4201(n4793 ,n4504 ,n4543);
    xnor g4202(n1783 ,n1636 ,n1728);
    nor g4203(n2531 ,n2514 ,n2490);
    nor g4204(n2040 ,n1990 ,n2033);
    or g4205(n5890 ,n5841 ,n5855);
    nand g4206(n1147 ,n23[15] ,n716);
    dff g4207(.RN(n1), .SN(1'b1), .CK(n0), .D(n1262), .Q(n19[0]));
    xnor g4208(n3039 ,n3002 ,n2921);
    nand g4209(n1402 ,n966 ,n1157);
    xnor g4210(n5445 ,n5166 ,n5146);
    or g4211(n3101 ,n38[10] ,n6560);
    nand g4212(n3970 ,n3835 ,n3921);
    xnor g4213(n3294 ,n3273 ,n3259);
    not g4214(n172 ,n171);
    nand g4215(n1943 ,n1860 ,n1916);
    xnor g4216(n696 ,n561 ,n26[5]);
    xnor g4217(n4333 ,n4320 ,n4302);
    xnor g4218(n5612 ,n5430 ,n5228);
    nand g4219(n5093 ,n4746 ,n5000);
    nand g4220(n274 ,n182 ,n194);
    nand g4221(n4499 ,n4378 ,n20[2]);
    nor g4222(n780 ,n606 ,n717);
    xnor g4223(n1811 ,n1765 ,n1646);
    nand g4224(n79 ,n65 ,n55);
    nand g4225(n5806 ,n5660 ,n5715);
    nor g4226(n2546 ,n2496 ,n2536);
    xnor g4227(n3175 ,n3133 ,n38[10]);
    xor g4228(n40[2] ,n6609 ,n38[3]);
    nand g4229(n1187 ,n4[5] ,n713);
    nand g4230(n1639 ,n1605 ,n1632);
    nand g4231(n4858 ,n4616 ,n4472);
    nand g4232(n6298 ,n40[2] ,n6250);
    nand g4233(n5560 ,n5169 ,n5455);
    or g4234(n4285 ,n4229 ,n4269);
    nand g4235(n6371 ,n6584 ,n6247);
    xnor g4236(n5818 ,n5751 ,n5632);
    nor g4237(n6479 ,n6383 ,n6463);
    or g4238(n5326 ,n5200 ,n5199);
    xnor g4239(n2419 ,n2372 ,n2322);
    nand g4240(n2274 ,n2117 ,n2239);
    xnor g4241(n5998 ,n5906 ,n5952);
    xnor g4242(n5614 ,n5429 ,n5353);
    nor g4243(n5774 ,n5551 ,n5704);
    not g4244(n2052 ,n2051);
    nand g4245(n1355 ,n893 ,n1108);
    not g4246(n711 ,n712);
    nand g4247(n5000 ,n4669 ,n4863);
    not g4248(n4517 ,n4516);
    not g4249(n5206 ,n5205);
    dff g4250(.RN(n1), .SN(1'b1), .CK(n0), .D(n1295), .Q(n11[9]));
    xnor g4251(n3908 ,n3757 ,n3517);
    xnor g4252(n2525 ,n2493 ,n2504);
    xnor g4253(n5425 ,n5193 ,n5297);
    nand g4254(n5488 ,n5402 ,n5289);
    xnor g4255(n5758 ,n5605 ,n5606);
    nand g4256(n1263 ,n648 ,n770);
    nand g4257(n4215 ,n4194 ,n4184);
    not g4258(n3903 ,n3902);
    xnor g4259(n4953 ,n4679 ,n4675);
    xnor g4260(n431 ,n357 ,n291);
    nor g4261(n2562 ,n2561 ,n2531);
    nand g4262(n1067 ,n10[13] ,n711);
    nand g4263(n4569 ,n4389 ,n20[5]);
    nand g4264(n1271 ,n851 ,n1018);
    not g4265(n3495 ,n19[3]);
    nand g4266(n6016 ,n5921 ,n5978);
    nand g4267(n5367 ,n5128 ,n5157);
    xnor g4268(n6114 ,n6057 ,n5970);
    not g4269(n3886 ,n3885);
    nand g4270(n1371 ,n820 ,n1122);
    dff g4271(.RN(n1), .SN(1'b1), .CK(n0), .D(n1433), .Q(n10[7]));
    not g4272(n4409 ,n21[3]);
    nand g4273(n1763 ,n1696 ,n1704);
    nand g4274(n5992 ,n5894 ,n5943);
    nand g4275(n3590 ,n3472 ,n3484);
    nand g4276(n6330 ,n38[14] ,n6246);
    xnor g4277(n6557 ,n4323 ,n4331);
    nand g4278(n5923 ,n5876 ,n5868);
    nand g4279(n3595 ,n3466 ,n3486);
    nand g4280(n4458 ,n20[3] ,n4367);
    xnor g4281(n5646 ,n5419 ,n5202);
    nand g4282(n3114 ,n6574 ,n6551);
    or g4283(n469 ,n389 ,n449);
    nand g4284(n5085 ,n4766 ,n5013);
    nand g4285(n2389 ,n2270 ,n2348);
    nand g4286(n1621 ,n1584 ,n1612);
    xnor g4287(n449 ,n393 ,n370);
    xnor g4288(n6187 ,n6160 ,n6147);
    not g4289(n4007 ,n3991);
    not g4290(n2999 ,n2991);
    not g4291(n3634 ,n3633);
    xnor g4292(n5313 ,n5150 ,n4784);
    not g4293(n157 ,n156);
    nand g4294(n1455 ,n1120 ,n1368);
    nor g4295(n6248 ,n25[0] ,n6222);
    nand g4296(n925 ,n34[9] ,n717);
    nand g4297(n1015 ,n12[9] ,n711);
    nor g4298(n2811 ,n2735 ,n2785);
    nand g4299(n3565 ,n3468 ,n3476);
    nand g4300(n5790 ,n5621 ,n5722);
    nand g4301(n4197 ,n4118 ,n4169);
    not g4302(n713 ,n714);
    xnor g4303(n4233 ,n4178 ,n4172);
    xnor g4304(n4057 ,n3948 ,n3908);
    not g4305(n5083 ,n5082);
    not g4306(n3482 ,n3487);
    nand g4307(n1035 ,n31[5] ,n720);
    nand g4308(n2099 ,n2080 ,n2073);
    xnor g4309(n6579 ,n2008 ,n2030);
    xnor g4310(n5529 ,n5308 ,n5110);
    nand g4311(n4640 ,n4378 ,n20[3]);
    xnor g4312(n6549 ,n3386 ,n3328);
    nand g4313(n842 ,n19[3] ,n714);
    nand g4314(n4330 ,n4320 ,n4302);
    xnor g4315(n3403 ,n6556 ,n39[7]);
    or g4316(n2575 ,n40[5] ,n6516);
    nand g4317(n553 ,n438 ,n552);
    nand g4318(n4621 ,n4389 ,n20[1]);
    dff g4319(.RN(n1), .SN(1'b1), .CK(n0), .D(n1362), .Q(n23[8]));
    nor g4320(n6485 ,n6431 ,n6475);
    not g4321(n1850 ,n1843);
    not g4322(n1955 ,n1954);
    nand g4323(n81 ,n67 ,n49);
    xnor g4324(n6126 ,n6095 ,n6106);
    nand g4325(n6393 ,n6270 ,n6321);
    nand g4326(n1123 ,n31[1] ,n720);
    dff g4327(.RN(n1), .SN(1'b1), .CK(n0), .D(n1442), .Q(n12[11]));
    nor g4328(n2735 ,n2567 ,n2628);
    xnor g4329(n5302 ,n5113 ,n5086);
    not g4330(n4781 ,n4780);
    xnor g4331(n6552 ,n4092 ,n4046);
    nand g4332(n6012 ,n5934 ,n5995);
    dff g4333(.RN(n1), .SN(1'b1), .CK(n0), .D(n1274), .Q(n16[2]));
    nor g4334(n2880 ,n2800 ,n2807);
    nor g4335(n1891 ,n1809 ,n1851);
    not g4336(n4958 ,n4957);
    xnor g4337(n6591 ,n3223 ,n3249);
    nor g4338(n735 ,n589 ,n710);
    nor g4339(n6541 ,n3287 ,n3317);
    nand g4340(n4464 ,n21[7] ,n4365);
    xnor g4341(n2298 ,n2245 ,n2120);
    xnor g4342(n6593 ,n3217 ,n3237);
    nand g4343(n1769 ,n1693 ,n1716);
    not g4344(n5162 ,n5161);
    nand g4345(n936 ,n34[11] ,n717);
    nor g4346(n766 ,n595 ,n723);
    xor g4347(n4915 ,n4525 ,n4599);
    or g4348(n6090 ,n6004 ,n6066);
    xnor g4349(n5521 ,n5310 ,n5107);
    or g4350(n2813 ,n2732 ,n2792);
    nand g4351(n5010 ,n4678 ,n4846);
    xnor g4352(n2075 ,n20[1] ,n21[1]);
    nor g4353(n3371 ,n6581 ,n3370);
    xnor g4354(n1604 ,n19[2] ,n19[1]);
    nor g4355(n6450 ,n6402 ,n6401);
    dff g4356(.RN(n1), .SN(1'b1), .CK(n0), .D(n1366), .Q(n23[6]));
    nand g4357(n1155 ,n6[4] ,n713);
    nor g4358(n6246 ,n25[0] ,n6223);
    nand g4359(n6082 ,n5999 ,n6046);
    or g4360(n790 ,n715 ,n704);
    nor g4361(n6470 ,n6408 ,n6390);
    nor g4362(n4780 ,n4548 ,n4664);
    not g4363(n3276 ,n36[3]);
    xnor g4364(n4935 ,n4633 ,n4489);
    nand g4365(n4985 ,n4542 ,n4800);
    xnor g4366(n3221 ,n3164 ,n3181);
    nand g4367(n3983 ,n3843 ,n3898);
    xnor g4368(n1954 ,n1900 ,n1846);
    nand g4369(n1457 ,n1123 ,n1372);
    nor g4370(n2454 ,n2400 ,n2425);
    nand g4371(n3164 ,n3113 ,n3146);
    nand g4372(n3871 ,n3666 ,n3813);
    nand g4373(n658 ,n16[2] ,n23[2]);
    xnor g4374(n3214 ,n3158 ,n3179);
    nand g4375(n35[12] ,n6454 ,n6486);
    not g4376(n566 ,n17[4]);
    nor g4377(n2613 ,n2565 ,n2584);
    xnor g4378(n3899 ,n3744 ,n3572);
    xnor g4379(n5776 ,n5601 ,n5589);
    nand g4380(n5568 ,n5342 ,n5482);
    xnor g4381(n2890 ,n2675 ,n2799);
    xnor g4382(n1550 ,n24[7] ,n131);
    or g4383(n5239 ,n4793 ,n5067);
    not g4384(n4402 ,n20[7]);
    xnor g4385(n689 ,n23[5] ,n34[5]);
    nand g4386(n5947 ,n5816 ,n5886);
    or g4387(n3693 ,n3546 ,n3502);
    xnor g4388(n5209 ,n4895 ,n4513);
    not g4389(n2791 ,n2790);
    xnor g4390(n86 ,n69 ,n57);
    xnor g4391(n6116 ,n6056 ,n6005);
    dff g4392(.RN(n1), .SN(1'b1), .CK(n0), .D(n1223), .Q(n28[1]));
    nand g4393(n1682 ,n1586 ,n1655);
    nand g4394(n1393 ,n947 ,n1149);
    not g4395(n351 ,n350);
    xnor g4396(n3888 ,n3753 ,n3631);
    nand g4397(n6391 ,n6334 ,n6333);
    or g4398(n3675 ,n3575 ,n3580);
    or g4399(n4053 ,n3900 ,n4022);
    nand g4400(n6244 ,n41[6] ,n6594);
    nand g4401(n4349 ,n4348 ,n4337);
    xnor g4402(n4178 ,n4104 ,n4060);
    xnor g4403(n462 ,n425 ,n356);
    nand g4404(n5954 ,n5845 ,n5890);
    not g4405(n1976 ,n1975);
    nand g4406(n1157 ,n6[3] ,n713);
    nand g4407(n3503 ,n3472 ,n3485);
    nor g4408(n6110 ,n6106 ,n6096);
    not g4409(n4417 ,n21[7]);
    not g4410(n155 ,n154);
    nor g4411(n3394 ,n6562 ,n6547);
    xnor g4412(n4941 ,n4476 ,n4566);
    nand g4413(n1085 ,n10[2] ,n555);
    or g4414(n4742 ,n4579 ,n4451);
    nand g4415(n6302 ,n6532 ,n6251);
    nand g4416(n5043 ,n4552 ,n4859);
    dff g4417(.RN(n1), .SN(1'b1), .CK(n0), .D(n1395), .Q(n21[5]));
    or g4418(n1861 ,n1749 ,n1805);
    nand g4419(n2993 ,n2925 ,n2955);
    or g4420(n617 ,n22[4] ,n22[5]);
    nand g4421(n1023 ,n3[3] ,n557);
    dff g4422(.RN(n1), .SN(1'b1), .CK(n0), .D(n1242), .Q(n33[0]));
    xnor g4423(n4250 ,n4210 ,n4185);
    xnor g4424(n6175 ,n6154 ,n6113);
    nand g4425(n5265 ,n5114 ,n5109);
    nand g4426(n189 ,n170 ,n144);
    nand g4427(n2593 ,n40[7] ,n6518);
    nand g4428(n3815 ,n3550 ,n3722);
    nand g4429(n905 ,n34[15] ,n717);
    not g4430(n52 ,n37[0]);
    nand g4431(n5113 ,n4762 ,n5011);
    xnor g4432(n5350 ,n5055 ,n5094);
    nand g4433(n1122 ,n1530 ,n716);
    nand g4434(n621 ,n18[0] ,n559);
    nand g4435(n1020 ,n12[7] ,n710);
    xor g4436(n39[3] ,n6615 ,n38[3]);
    buf g4437(n13[5], n11[5]);
    nand g4438(n1171 ,n5[3] ,n557);
    xor g4439(n4900 ,n4547 ,n4438);
    xor g4440(n6610 ,n6550 ,n39[1]);
    nand g4441(n5673 ,n5522 ,n5521);
    or g4442(n6150 ,n6079 ,n6128);
    nand g4443(n4597 ,n20[5] ,n4371);
    nand g4444(n3229 ,n3198 ,n3228);
    xor g4445(n1833 ,n1784 ,n1751);
    not g4446(n3267 ,n3266);
    xor g4447(n3766 ,n3561 ,n3540);
    nor g4448(n1890 ,n1813 ,n1849);
    not g4449(n2794 ,n2793);
    dff g4450(.RN(n1), .SN(1'b1), .CK(n0), .D(n1230), .Q(n12[14]));
    xnor g4451(n5453 ,n5230 ,n5141);
    nand g4452(n4594 ,n20[2] ,n4373);
    nor g4453(n5655 ,n5517 ,n5545);
    xnor g4454(n4230 ,n4093 ,n4198);
    nand g4455(n6045 ,n5949 ,n6006);
    nand g4456(n4558 ,n20[1] ,n4374);
    nor g4457(n3423 ,n3399 ,n3422);
    nand g4458(n2095 ,n6538 ,n2085);
    nand g4459(n3824 ,n3562 ,n3732);
    not g4460(n5581 ,n5580);
    nor g4461(n2455 ,n2401 ,n2424);
    nand g4462(n5561 ,n5404 ,n5493);
    nand g4463(n4497 ,n21[5] ,n4363);
    xnor g4464(n2074 ,n21[4] ,n21[3]);
    nand g4465(n6354 ,n6583 ,n6247);
    nand g4466(n4816 ,n4598 ,n4610);
    nand g4467(n2989 ,n2927 ,n2954);
    or g4468(n4327 ,n4318 ,n4310);
    nand g4469(n6423 ,n6291 ,n6353);
    nor g4470(n2438 ,n2353 ,n2404);
    xnor g4471(n312 ,n247 ,n200);
    nand g4472(n3591 ,n3484 ,n19[4]);
    or g4473(n2930 ,n2854 ,n2910);
    nor g4474(n3635 ,n3491 ,n3493);
    not g4475(n245 ,n244);
    nor g4476(n5654 ,n5501 ,n5531);
    xnor g4477(n667 ,n19[5] ,n27[5]);
    xnor g4478(n5880 ,n5769 ,n5551);
    nand g4479(n994 ,n19[5] ,n556);
    nand g4480(n649 ,n19[2] ,n27[2]);
    xnor g4481(n3131 ,n6585 ,n6562);
    nand g4482(n1749 ,n1665 ,n1732);
    xnor g4483(n6083 ,n6025 ,n6035);
    nand g4484(n1765 ,n1687 ,n1718);
    nand g4485(n278 ,n193 ,n217);
    nor g4486(n6161 ,n6115 ,n6149);
    nand g4487(n951 ,n35[9] ,n554);
    nand g4488(n4859 ,n4489 ,n4633);
    nand g4489(n650 ,n16[4] ,n23[4]);
    nand g4490(n4695 ,n21[3] ,n4386);
    nand g4491(n1478 ,n827 ,n1252);
    nand g4492(n3291 ,n3277 ,n3267);
    not g4493(n3471 ,n37[3]);
    nand g4494(n2051 ,n2027 ,n2050);
    nand g4495(n98 ,n79 ,n97);
    nand g4496(n546 ,n534 ,n545);
    nand g4497(n4478 ,n21[4] ,n4367);
    nand g4498(n3942 ,n3671 ,n3857);
    nor g4499(n2680 ,n2565 ,n2633);
    nand g4500(n887 ,n27[13] ,n715);
    not g4501(n3469 ,n37[0]);
    nand g4502(n1672 ,n1580 ,n1649);
    nand g4503(n843 ,n19[2] ,n556);
    nand g4504(n1117 ,n31[6] ,n720);
    xor g4505(n4938 ,n4546 ,n4462);
    or g4506(n3189 ,n3163 ,n3176);
    nand g4507(n3592 ,n3466 ,n3478);
    nand g4508(n1466 ,n937 ,n1385);
    nand g4509(n4441 ,n20[0] ,n4371);
    nand g4510(n35[1] ,n6456 ,n6455);
    nor g4511(n6456 ,n6398 ,n6413);
    nand g4512(n5397 ,n5286 ,n5159);
    nor g4513(n3396 ,n6563 ,n6548);
    or g4514(n5842 ,n5718 ,n5786);
    xnor g4515(n5534 ,n5304 ,n5133);
    not g4516(n4369 ,n4368);
    nor g4517(n1842 ,n1774 ,n1823);
    nand g4518(n4426 ,n4382 ,n20[5]);
    nand g4519(n505 ,n456 ,n484);
    nand g4520(n2387 ,n2322 ,n2349);
    xnor g4521(n4973 ,n4470 ,n4502);
    nor g4522(n2653 ,n2565 ,n2595);
    not g4523(n3281 ,n3280);
    nand g4524(n5075 ,n4745 ,n4992);
    or g4525(n4290 ,n4245 ,n4270);
    xnor g4526(n5829 ,n5700 ,n5688);
    nand g4527(n3560 ,n3474 ,n3481);
    nand g4528(n1238 ,n1094 ,n748);
    not g4529(n719 ,n720);
    xnor g4530(n5353 ,n4971 ,n5142);
    xor g4531(n5622 ,n5432 ,n5213);
    not g4532(n3550 ,n3549);
    or g4533(n4721 ,n4638 ,n4576);
    nand g4534(n1666 ,n1588 ,n1651);
    nand g4535(n5578 ,n5338 ,n5483);
    xnor g4536(n3777 ,n3638 ,n3625);
    xnor g4537(n5824 ,n5702 ,n5519);
    nor g4538(n729 ,n572 ,n710);
    nand g4539(n5398 ,n5198 ,n5156);
    not g4540(n1882 ,n1881);
    dff g4541(.RN(n1), .SN(1'b1), .CK(n0), .D(n1258), .Q(n19[3]));
    nor g4542(n2277 ,n2108 ,n2230);
    nand g4543(n2245 ,n2138 ,n2198);
    xnor g4544(n4907 ,n4461 ,n4594);
    nand g4545(n3364 ,n6579 ,n3363);
    nand g4546(n3556 ,n3485 ,n19[0]);
    xnor g4547(n4951 ,n4618 ,n4427);
    nand g4548(n6400 ,n6267 ,n6327);
    nand g4549(n5080 ,n4719 ,n5005);
    nand g4550(n4801 ,n4498 ,n4500);
    not g4551(n4383 ,n36[3]);
    nor g4552(n5791 ,n5666 ,n5724);
    nand g4553(n6370 ,n39[1] ,n6248);
    not g4554(n5195 ,n5194);
    xnor g4555(n5293 ,n4912 ,n4688);
    nand g4556(n2199 ,n6538 ,n2149);
    nor g4557(n3997 ,n3865 ,n3886);
    or g4558(n5672 ,n5547 ,n5523);
    xnor g4559(n5690 ,n5496 ,n5587);
    xor g4560(n2085 ,n21[0] ,n20[0]);
    nand g4561(n1089 ,n1553 ,n716);
    nand g4562(n1218 ,n926 ,n771);
    nor g4563(n738 ,n618 ,n717);
    nand g4564(n5564 ,n5168 ,n5456);
    nand g4565(n3836 ,n3682 ,n3780);
    xnor g4566(n5429 ,n5174 ,n5115);
    nand g4567(n35[4] ,n6466 ,n6485);
    xnor g4568(n3759 ,n3527 ,n3579);
    nand g4569(n2204 ,n6541 ,n2149);
    xnor g4570(n373 ,n305 ,n204);
    nand g4571(n3234 ,n3191 ,n3233);
    nand g4572(n1044 ,n11[12] ,n711);
    nand g4573(n4841 ,n4579 ,n4451);
    nand g4574(n1040 ,n11[14] ,n710);
    or g4575(n3833 ,n3793 ,n3786);
    nand g4576(n6278 ,n6551 ,n6251);
    nand g4577(n3232 ,n3190 ,n3231);
    nand g4578(n3837 ,n3683 ,n3779);
    nor g4579(n2935 ,n2842 ,n2909);
    nand g4580(n5066 ,n4792 ,n4955);
    xnor g4581(n497 ,n403 ,n474);
    nand g4582(n5039 ,n4547 ,n4871);
    or g4583(n3676 ,n3539 ,n3599);
    nand g4584(n1431 ,n995 ,n1186);
    nand g4585(n6431 ,n6294 ,n6365);
    nand g4586(n3571 ,n3474 ,n3482);
    nand g4587(n226 ,n170 ,n150);
    nand g4588(n4344 ,n4314 ,n4339);
    dff g4589(.RN(n1), .SN(1'b1), .CK(n0), .D(n1236), .Q(n12[0]));
    xnor g4590(n2875 ,n2790 ,n2665);
    xnor g4591(n3881 ,n3786 ,n3543);
    xnor g4592(n5694 ,n5522 ,n5521);
    or g4593(n5987 ,n5908 ,n5932);
    xnor g4594(n38[10] ,n2544 ,n2553);
    or g4595(n1596 ,n1570 ,n1574);
    xnor g4596(n3892 ,n3771 ,n3567);
    not g4597(n2401 ,n2400);
    nor g4598(n1549 ,n135 ,n133);
    nor g4599(n2733 ,n2567 ,n2627);
    nor g4600(n834 ,n566 ,n721);
    not g4601(n4790 ,n4789);
    or g4602(n753 ,n717 ,n689);
    nand g4603(n2103 ,n2069 ,n2082);
    nand g4604(n5843 ,n5631 ,n5776);
    not g4605(n6130 ,n6129);
    nor g4606(n592 ,n21[0] ,n30[0]);
    xnor g4607(n5220 ,n4909 ,n4560);
    not g4608(n5881 ,n5880);
    nand g4609(n6342 ,n38[15] ,n6246);
    nand g4610(n6007 ,n5918 ,n5965);
    nand g4611(n931 ,n29[3] ,n721);
    nand g4612(n5853 ,n5734 ,n5795);
    nand g4613(n35[9] ,n6461 ,n6457);
    xnor g4614(n4138 ,n4064 ,n3999);
    xor g4615(n5214 ,n4914 ,n4482);
    nor g4616(n3799 ,n3628 ,n3738);
    xnor g4617(n6489 ,n3212 ,n3227);
    nand g4618(n2221 ,n2146 ,n2186);
    or g4619(n4714 ,n4484 ,n4479);
    xnor g4620(n6615 ,n3344 ,n3351);
    buf g4621(n37[3] ,n1503);
    nand g4622(n3079 ,n3056 ,n3078);
    or g4623(n4117 ,n4062 ,n4061);
    nand g4624(n5686 ,n5502 ,n5555);
    nand g4625(n5802 ,n5673 ,n5703);
    buf g4626(n14[10], n11[10]);
    nor g4627(n1734 ,n1589 ,n1699);
    or g4628(n4242 ,n4185 ,n4210);
    nand g4629(n2206 ,n6541 ,n2150);
    nand g4630(n3141 ,n6552 ,n3105);
    nor g4631(n3821 ,n3615 ,n3735);
    nand g4632(n1064 ,n11[0] ,n710);
    nand g4633(n6237 ,n6226 ,n6227);
    xor g4634(n40[6] ,n38[7] ,n6605);
    xnor g4635(n5307 ,n5070 ,n5080);
    nor g4636(n2709 ,n2567 ,n2616);
    dff g4637(.RN(n1), .SN(1'b1), .CK(n0), .D(n1445), .Q(n12[8]));
    nor g4638(n4155 ,n4054 ,n4099);
    nand g4639(n2980 ,n2966 ,n2944);
    dff g4640(.RN(n1), .SN(1'b1), .CK(n0), .D(n1415), .Q(n20[3]));
    not g4641(n2117 ,n2118);
    nor g4642(n2753 ,n2600 ,n2719);
    nand g4643(n3117 ,n6576 ,n6553);
    xnor g4644(n1523 ,n538 ,n544);
    dff g4645(.RN(n1), .SN(1'b1), .CK(n0), .D(n1420), .Q(n26[5]));
    nor g4646(n2832 ,n2658 ,n2748);
    nand g4647(n4200 ,n4117 ,n4159);
    nand g4648(n3369 ,n3330 ,n3368);
    nand g4649(n3570 ,n3470 ,n3478);
    xnor g4650(n2024 ,n1987 ,n1966);
    not g4651(n3406 ,n3405);
    nand g4652(n3158 ,n3115 ,n3137);
    not g4653(n3275 ,n3274);
    or g4654(n3659 ,n3608 ,n3504);
    nor g4655(n4034 ,n3909 ,n4005);
    nand g4656(n1093 ,n33[7] ,n555);
    nor g4657(n1592 ,n1574 ,n19[1]);
    nand g4658(n4867 ,n4615 ,n4471);
    not g4659(n2661 ,n2660);
    xnor g4660(n5204 ,n4920 ,n4604);
    not g4661(n5197 ,n5196);
    nor g4662(n2714 ,n2565 ,n2626);
    nand g4663(n985 ,n27[0] ,n715);
    not g4664(n3778 ,n3777);
    nand g4665(n184 ,n172 ,n152);
    nand g4666(n3231 ,n3202 ,n3230);
    nand g4667(n1344 ,n1142 ,n951);
    nand g4668(n5479 ,n5089 ,n5358);
    nand g4669(n4615 ,n4384 ,n20[6]);
    nand g4670(n5136 ,n4763 ,n5021);
    nand g4671(n4158 ,n4084 ,n4113);
    xnor g4672(n3037 ,n3006 ,n2968);
    not g4673(n150 ,n149);
    nand g4674(n5798 ,n5643 ,n5710);
    or g4675(n3190 ,n3161 ,n3174);
    xnor g4676(n1524 ,n537 ,n542);
    nand g4677(n4465 ,n21[3] ,n4389);
    nand g4678(n1125 ,n31[0] ,n720);
    nand g4679(n6293 ,n40[10] ,n6250);
    nand g4680(n4280 ,n4227 ,n4267);
    nand g4681(n1179 ,n29[4] ,n724);
    xnor g4682(n1920 ,n1778 ,n1881);
    nand g4683(n5026 ,n4649 ,n4853);
    not g4684(n4366 ,n37[4]);
    nor g4685(n2638 ,n2566 ,n2588);
    not g4686(n2316 ,n2315);
    xor g4687(n366 ,n302 ,n207);
    nor g4688(n591 ,n22[4] ,n26[4]);
    nand g4689(n1047 ,n11[10] ,n555);
    nor g4690(n1901 ,n1778 ,n1882);
    xor g4691(n4893 ,n4511 ,n4478);
    nor g4692(n2603 ,n2567 ,n2586);
    nand g4693(n1617 ,n1586 ,n1612);
    nand g4694(n4347 ,n4334 ,n4346);
    nor g4695(n5720 ,n5607 ,n5635);
    not g4696(n2494 ,n2493);
    xor g4697(n40[13] ,n6598 ,n38[14]);
    nand g4698(n2084 ,n21[4] ,n2066);
    not g4699(n721 ,n722);
    not g4700(n4375 ,n36[7]);
    nor g4701(n3029 ,n2981 ,n3010);
    nand g4702(n1494 ,n1063 ,n1488);
    nand g4703(n4083 ,n3957 ,n4033);
    nand g4704(n4146 ,n4060 ,n4104);
    nor g4705(n2646 ,n2566 ,n2589);
    nand g4706(n536 ,n515 ,n522);
    xor g4707(n1542 ,n71 ,n53);
    xnor g4708(n2305 ,n2230 ,n2109);
    nand g4709(n1895 ,n1829 ,n1858);
    not g4710(n4005 ,n3989);
    nand g4711(n3064 ,n3029 ,n3038);
    nand g4712(n858 ,n16[1] ,n714);
    not g4713(n1569 ,n37[2]);
    nand g4714(n2194 ,n6534 ,n2148);
    xnor g4715(n3770 ,n3516 ,n3548);
    not g4716(n2408 ,n2407);
    xnor g4717(n5871 ,n5768 ,n5645);
    xor g4718(n6567 ,n5866 ,n5689);
    nor g4719(n2383 ,n2298 ,n2362);
    xnor g4720(n5769 ,n5618 ,n5529);
    xnor g4721(n3889 ,n3760 ,n3644);
    not g4722(n92 ,n91);
    nand g4723(n6381 ,n39[6] ,n6248);
    or g4724(n520 ,n516 ,n510);
    nand g4725(n4833 ,n4632 ,n4480);
    xnor g4726(n4909 ,n4460 ,n4571);
    nor g4727(n3028 ,n2977 ,n3016);
    dff g4728(.RN(n1), .SN(1'b1), .CK(n0), .D(n18[1]), .Q(n15[5]));
    nand g4729(n4477 ,n4384 ,n20[4]);
    xnor g4730(n5695 ,n5580 ,n5583);
    nor g4731(n5512 ,n5497 ,n5492);
    nand g4732(n5396 ,n5210 ,n5283);
    xor g4733(n4944 ,n4540 ,n4446);
    xnor g4734(n3882 ,n3787 ,n3576);
    nor g4735(n3562 ,n3496 ,n3500);
    not g4736(n2377 ,n2376);
    xnor g4737(n451 ,n391 ,n341);
    xnor g4738(n1641 ,n1618 ,n1613);
    nor g4739(n3350 ,n6567 ,n3349);
    nor g4740(n2694 ,n2568 ,n2622);
    xnor g4741(n4014 ,n3914 ,n3865);
    nand g4742(n80 ,n73 ,n51);
    nand g4743(n5110 ,n4727 ,n5050);
    nand g4744(n5991 ,n5844 ,n5916);
    xnor g4745(n681 ,n35[2] ,n31[2]);
    nand g4746(n1102 ,n33[2] ,n710);
    xnor g4747(n3898 ,n3759 ,n3636);
    nand g4748(n101 ,n89 ,n100);
    xnor g4749(n5210 ,n4932 ,n4662);
    nand g4750(n831 ,n34[1] ,n717);
    xnor g4751(n5765 ,n5641 ,n5535);
    xnor g4752(n1874 ,n1809 ,n1818);
    xnor g4753(n6570 ,n6196 ,n6209);
    nor g4754(n289 ,n203 ,n201);
    nor g4755(n4678 ,n4402 ,n4399);
    xnor g4756(n529 ,n513 ,n511);
    xnor g4757(n6571 ,n6203 ,n6211);
    nor g4758(n2437 ,n2058 ,n2408);
    not g4759(n130 ,n129);
    nor g4760(n2901 ,n2831 ,n2893);
    or g4761(n407 ,n342 ,n367);
    dff g4762(.RN(n1), .SN(1'b1), .CK(n0), .D(n1468), .Q(n22[1]));
    nand g4763(n5376 ,n5278 ,n5181);
    or g4764(n2573 ,n40[12] ,n6523);
    nand g4765(n200 ,n163 ,n153);
    nor g4766(n2335 ,n2260 ,n2314);
    nand g4767(n2188 ,n6534 ,n2149);
    xnor g4768(n5461 ,n5232 ,n5224);
    nand g4769(n6411 ,n6280 ,n6338);
    nand g4770(n3984 ,n3888 ,n3887);
    nand g4771(n2183 ,n6534 ,n2150);
    nand g4772(n3398 ,n6552 ,n39[3]);
    dff g4773(.RN(n1), .SN(1'b1), .CK(n0), .D(n1496), .Q(n18[1]));
    xnor g4774(n3296 ,n3275 ,n3257);
    xnor g4775(n6490 ,n3213 ,n3229);
    nand g4776(n1213 ,n34[1] ,n836);
    nand g4777(n3506 ,n3476 ,n19[7]);
    not g4778(n1931 ,n1930);
    nand g4779(n1335 ,n649 ,n742);
    xnor g4780(n5912 ,n5820 ,n5838);
    nand g4781(n3707 ,n3530 ,n3537);
    xnor g4782(n5642 ,n5433 ,n5151);
    not g4783(n3261 ,n3260);
    nand g4784(n5794 ,n5756 ,n5744);
    nand g4785(n5048 ,n4531 ,n4872);
    nand g4786(n1309 ,n1067 ,n955);
    dff g4787(.RN(n1), .SN(1'b1), .CK(n0), .D(n1237), .Q(n33[7]));
    xnor g4788(n38[2] ,n2373 ,n2319);
    nand g4789(n6292 ,n6571 ,n6254);
    nor g4790(n620 ,n563 ,n18[0]);
    nor g4791(n2614 ,n2565 ,n2588);
    nand g4792(n1222 ,n941 ,n778);
    xnor g4793(n5632 ,n5428 ,n5217);
    nand g4794(n134 ,n32[1] ,n32[0]);
    not g4795(n45 ,n44);
    nand g4796(n6184 ,n6151 ,n6164);
    nand g4797(n5379 ,n5280 ,n5158);
    nand g4798(n1225 ,n973 ,n880);
    nand g4799(n883 ,n34[12] ,n717);
    dff g4800(.RN(n1), .SN(1'b1), .CK(n0), .D(n1396), .Q(n27[13]));
    nand g4801(n4278 ,n4242 ,n4258);
    nand g4802(n2160 ,n6536 ,n2127);
    nand g4803(n5024 ,n4648 ,n4849);
    not g4804(n153 ,n175);
    nand g4805(n965 ,n27[9] ,n715);
    buf g4806(n14[0], n11[0]);
    nand g4807(n1124 ,n1532 ,n716);
    nand g4808(n194 ,n163 ,n155);
    nor g4809(n6001 ,n5933 ,n5975);
    not g4810(n2406 ,n2405);
    xnor g4811(n3126 ,n6564 ,n6587);
    nand g4812(n957 ,n35[11] ,n554);
    nand g4813(n1031 ,n3[0] ,n557);
    xor g4814(n4898 ,n4653 ,n4477);
    xnor g4815(n1797 ,n1747 ,n1750);
    not g4816(n46 ,n37[4]);
    nor g4817(n5247 ,n5139 ,n5134);
    nand g4818(n636 ,n19[6] ,n27[6]);
    nand g4819(n1342 ,n1139 ,n952);
    nand g4820(n6383 ,n6309 ,n6381);
    dff g4821(.RN(n1), .SN(1'b1), .CK(n0), .D(n1283), .Q(n1514));
    nand g4822(n4042 ,n3913 ,n3987);
    dff g4823(.RN(n1), .SN(1'b1), .CK(n0), .D(n1288), .Q(n11[13]));
    not g4824(n4962 ,n4961);
    not g4825(n5410 ,n5388);
    nand g4826(n4504 ,n21[4] ,n4374);
    xnor g4827(n5443 ,n5298 ,n5284);
    nor g4828(n4540 ,n4412 ,n4416);
    nand g4829(n2135 ,n6535 ,n2121);
    not g4830(n1567 ,n37[5]);
    nand g4831(n5789 ,n5620 ,n5723);
    nand g4832(n5354 ,n5093 ,n5239);
    nand g4833(n273 ,n229 ,n184);
    xnor g4834(n6488 ,n3226 ,n3154);
    xnor g4835(n394 ,n290 ,n353);
    nand g4836(n4611 ,n4386 ,n20[4]);
    nand g4837(n2002 ,n1919 ,n1981);
    xnor g4838(n5878 ,n5761 ,n5523);
    xnor g4839(n523 ,n498 ,n475);
    nor g4840(n2769 ,n2649 ,n2697);
    nand g4841(n400 ,n342 ,n367);
    nand g4842(n2592 ,n40[2] ,n6513);
    xnor g4843(n3171 ,n3126 ,n38[14]);
    xnor g4844(n6129 ,n6083 ,n6107);
    nand g4845(n5044 ,n4690 ,n4840);
    xor g4846(n39[2] ,n38[2] ,n6616);
    nand g4847(n6362 ,n38[13] ,n6246);
    nand g4848(n656 ,n22[1] ,n26[1]);
    nand g4849(n1707 ,n1584 ,n1676);
    nand g4850(n3042 ,n3008 ,n3024);
    not g4851(n556 ,n557);
    nand g4852(n1916 ,n1865 ,n1887);
    nor g4853(n2307 ,n2151 ,n2265);
    nand g4854(n1790 ,n1647 ,n1756);
    nand g4855(n5946 ,n5814 ,n5891);
    xnor g4856(n38[14] ,n2525 ,n2562);
    nor g4857(n3026 ,n2986 ,n3017);
    nor g4858(n3965 ,n3888 ,n3887);
    xnor g4859(n4008 ,n3904 ,n3891);
    nand g4860(n4127 ,n4062 ,n4061);
    nand g4861(n6375 ,n6578 ,n6247);
    nand g4862(n4865 ,n4494 ,n4572);
    xnor g4863(n2974 ,n2926 ,n2827);
    nand g4864(n4002 ,n3789 ,n3931);
    or g4865(n4335 ,n4319 ,n4324);
    nand g4866(n346 ,n249 ,n334);
    xnor g4867(n1956 ,n1814 ,n1910);
    nor g4868(n596 ,n9[3] ,n9[2]);
    nor g4869(n3679 ,n3521 ,n3589);
    dff g4870(.RN(n1), .SN(1'b1), .CK(n0), .D(n1272), .Q(n1504));
    xnor g4871(n4093 ,n3972 ,n4043);
    xnor g4872(n3911 ,n3773 ,n3554);
    or g4873(n789 ,n555 ,n687);
    not g4874(n3462 ,n3461);
    nand g4875(n4795 ,n4621 ,n4422);
    xor g4876(n4929 ,n4512 ,n4488);
    nand g4877(n5060 ,n4779 ,n4953);
    dff g4878(.RN(n1), .SN(1'b1), .CK(n0), .D(n1228), .Q(n27[0]));
    nand g4879(n4644 ,n21[3] ,n4367);
    nand g4880(n647 ,n21[7] ,n30[7]);
    or g4881(n5891 ,n5781 ,n5835);
    nor g4882(n5805 ,n5651 ,n5706);
    not g4883(n5279 ,n5278);
    or g4884(n755 ,n720 ,n692);
    nand g4885(n5941 ,n5757 ,n5887);
    or g4886(n4754 ,n4636 ,n4452);
    xnor g4887(n2077 ,n21[7] ,n20[7]);
    xnor g4888(n3038 ,n3003 ,n2919);
    nand g4889(n3727 ,n3645 ,n3646);
    not g4890(n1700 ,n1699);
    xnor g4891(n1784 ,n1648 ,n1725);
    xnor g4892(n5610 ,n5426 ,n5072);
    nor g4893(n3428 ,n3404 ,n3427);
    nand g4894(n4261 ,n4220 ,n4235);
    nand g4895(n6138 ,n6064 ,n6118);
    nor g4896(n3692 ,n3616 ,n3640);
    nand g4897(n1231 ,n1003 ,n885);
    nor g4898(n2062 ,n20[5] ,n21[5]);
    nand g4899(n230 ,n161 ,n150);
    or g4900(n6164 ,n6147 ,n6144);
    nand g4901(n1046 ,n11[11] ,n710);
    not g4902(n4552 ,n4551);
    nand g4903(n2990 ,n2928 ,n2947);
    nand g4904(n5031 ,n4514 ,n4848);
    not g4905(n5811 ,n5810);
    nand g4906(n5257 ,n5139 ,n5134);
    nand g4907(n3975 ,n3661 ,n3932);
    not g4908(n44 ,n37[6]);
    nand g4909(n579 ,n558 ,n559);
    xnor g4910(n3404 ,n6542 ,n6557);
    nand g4911(n4855 ,n4466 ,n4606);
    nand g4912(n1456 ,n1121 ,n1369);
    nand g4913(n4874 ,n4487 ,n4488);
    xnor g4914(n461 ,n421 ,n405);
    nand g4915(n5139 ,n4725 ,n5004);
    nand g4916(n334 ,n235 ,n274);
    nand g4917(n3509 ,n3462 ,n3486);
    nor g4918(n2598 ,n2567 ,n2585);
    nor g4919(n1678 ,n1637 ,n1653);
    or g4920(n4741 ,n4618 ,n4427);
    nor g4921(n2683 ,n2568 ,n2629);
    or g4922(n484 ,n429 ,n462);
    nor g4923(n4100 ,n3999 ,n4064);
    nor g4924(n1962 ,n1868 ,n1929);
    nor g4925(n745 ,n26[0] ,n706);
    nand g4926(n4187 ,n4091 ,n4158);
    or g4927(n5236 ,n5108 ,n5085);
    nand g4928(n3835 ,n3733 ,n3778);
    xnor g4929(n4029 ,n3916 ,n3852);
    nand g4930(n642 ,n31[1] ,n35[1]);
    nand g4931(n1434 ,n718 ,n1198);
    or g4932(n470 ,n417 ,n448);
    nor g4933(n1915 ,n1834 ,n1894);
    not g4934(n1986 ,n1985);
    nand g4935(n1159 ,n6[2] ,n713);
    nand g4936(n2142 ,n6534 ,n2122);
    nand g4937(n5358 ,n5073 ,n5194);
    dff g4938(.RN(n1), .SN(1'b1), .CK(n0), .D(n1315), .Q(n33[13]));
    or g4939(n1595 ,n1564 ,n1572);
    nand g4940(n6101 ,n6058 ,n6082);
    xnor g4941(n5305 ,n5081 ,n5125);
    nor g4942(n722 ,n18[2] ,n623);
    nand g4943(n5127 ,n4748 ,n4985);
    or g4944(n532 ,n515 ,n522);
    not g4945(n1614 ,n1613);
    xnor g4946(n2295 ,n2242 ,n2118);
    nand g4947(n550 ,n514 ,n549);
    xnor g4948(n1520 ,n497 ,n550);
    nand g4949(n1026 ,n3[2] ,n557);
    nand g4950(n4483 ,n21[7] ,n4386);
    nand g4951(n859 ,n21[2] ,n714);
    xnor g4952(n3907 ,n3774 ,n3580);
    nand g4953(n3201 ,n3153 ,n3170);
    xor g4954(n6535 ,n3302 ,n3306);
    not g4955(n1191 ,n1129);
    nand g4956(n4031 ,n3871 ,n3996);
    nand g4957(n1721 ,n1619 ,n1688);
    nand g4958(n1175 ,n1534 ,n557);
    xnor g4959(n1922 ,n1878 ,n1807);
    xnor g4960(n5229 ,n4885 ,n4426);
    xnor g4961(n38[0] ,n2108 ,n2125);
    nand g4962(n6403 ,n6318 ,n6328);
    nor g4963(n2657 ,n2565 ,n2587);
    nand g4964(n4422 ,n20[3] ,n4371);
    xnor g4965(n3764 ,n3596 ,n3583);
    nand g4966(n4292 ,n4226 ,n4273);
    nand g4967(n5400 ,n5096 ,n5253);
    buf g4968(n14[6], n10[6]);
    nor g4969(n1786 ,n1746 ,n1749);
    xnor g4970(n4901 ,n4579 ,n4451);
    nand g4971(n5548 ,n5320 ,n5473);
    dff g4972(.RN(n1), .SN(1'b1), .CK(n0), .D(n1356), .Q(n32[5]));
    not g4973(n4385 ,n36[1]);
    or g4974(n2903 ,n2789 ,n2873);
    nand g4975(n6137 ,n6029 ,n6112);
    nor g4976(n836 ,n562 ,n721);
    nand g4977(n3921 ,n3852 ,n3832);
    nor g4978(n2910 ,n2836 ,n2886);
    xnor g4979(n3224 ,n3160 ,n3171);
    nor g4980(n2471 ,n2450 ,n2418);
    nand g4981(n1146 ,n33[12] ,n710);
    dff g4982(.RN(n1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n32[1]));
    nand g4983(n6380 ,n6509 ,n6249);
    nand g4984(n1354 ,n1082 ,n907);
    nand g4985(n1495 ,n916 ,n1489);
    xor g4986(n39[7] ,n6611 ,n38[7]);
    dff g4987(.RN(n1), .SN(1'b1), .CK(n0), .D(n1439), .Q(n29[1]));
    nand g4988(n5566 ,n5497 ,n5492);
    nor g4989(n1904 ,n1840 ,n1890);
    nand g4990(n117 ,n115 ,n116);
    nor g4991(n1950 ,n1938 ,n1933);
    not g4992(n3258 ,n37[4]);
    nand g4993(n1324 ,n1084 ,n919);
    nand g4994(n5906 ,n5790 ,n5846);
    xnor g4995(n1752 ,n1657 ,n1646);
    or g4996(n6142 ,n6127 ,n6065);
    nor g4997(n1834 ,n1775 ,n1821);
    not g4998(n3624 ,n3623);
    xnor g4999(n6613 ,n3360 ,n41[5]);
    not g5000(n42 ,n37[7]);
    nand g5001(n1982 ,n1922 ,n1951);
    nand g5002(n513 ,n493 ,n505);
    xnor g5003(n2982 ,n2894 ,n2941);
    nor g5004(n127 ,n120 ,n126);
    not g5005(n3830 ,n3829);
    nand g5006(n871 ,n33[10] ,n712);
    not g5007(n3734 ,n3733);
    not g5008(n5411 ,n5392);
    xnor g5009(n1970 ,n1908 ,n1930);
    xnor g5010(n4207 ,n4143 ,n4085);
    nand g5011(n3543 ,n3486 ,n19[3]);
    not g5012(n5412 ,n5395);
    nand g5013(n5250 ,n5141 ,n5060);
    nor g5014(n5847 ,n5806 ,n5783);
    nand g5015(n1200 ,n584 ,n745);
    xor g5016(n6526 ,n6588 ,n6532);
    or g5017(n5338 ,n5166 ,n5165);
    or g5018(n3054 ,n3030 ,n3040);
    not g5019(n3523 ,n3522);
    xnor g5020(n5430 ,n5199 ,n5200);
    not g5021(n4373 ,n4372);
    nand g5022(n1628 ,n1608 ,n1602);
    nand g5023(n126 ,n24[3] ,n125);
    not g5024(n4703 ,n4702);
    nand g5025(n1252 ,n28[3] ,n1190);
    nand g5026(n2202 ,n2093 ,n2159);
    dff g5027(.RN(n1), .SN(1'b1), .CK(n0), .D(n1196), .Q(n10[8]));
    xnor g5028(n5780 ,n5594 ,n5505);
    nand g5029(n870 ,n33[11] ,n712);
    nand g5030(n2163 ,n6537 ,n2127);
    nand g5031(n3704 ,n3524 ,n3542);
    nand g5032(n6064 ,n6026 ,n6035);
    not g5033(n2341 ,n2334);
    nor g5034(n610 ,n33[8] ,n35[8]);
    nand g5035(n3375 ,n3338 ,n3374);
    xor g5036(n3758 ,n3562 ,n3582);
    nand g5037(n6295 ,n40[13] ,n6250);
    nor g5038(n1998 ,n1955 ,n1984);
    xnor g5039(n316 ,n242 ,n246);
    nor g5040(n3788 ,n3525 ,n3680);
    nand g5041(n4475 ,n20[7] ,n4374);
    dff g5042(.RN(n1), .SN(1'b1), .CK(n0), .D(n1317), .Q(n34[15]));
    nand g5043(n1671 ,n1588 ,n1649);
    nor g5044(n4553 ,n4408 ,n4399);
    nand g5045(n193 ,n165 ,n148);
    nor g5046(n2771 ,n2611 ,n2722);
    nand g5047(n3504 ,n3482 ,n19[5]);
    nor g5048(n2841 ,n2668 ,n2782);
    nand g5049(n5388 ,n5171 ,n5170);
    nand g5050(n6324 ,n6581 ,n6247);
    nand g5051(n3091 ,n3060 ,n3090);
    nand g5052(n4170 ,n4001 ,n4128);
    nand g5053(n5583 ,n5328 ,n5472);
    nand g5054(n4428 ,n4389 ,n20[4]);
    nor g5055(n2795 ,n2607 ,n2682);
    nand g5056(n5489 ,n5296 ,n5389);
    dff g5057(.RN(n1), .SN(1'b1), .CK(n0), .D(n1239), .Q(n33[5]));
    xnor g5058(n4103 ,n4014 ,n3885);
    nor g5059(n2835 ,n2736 ,n2784);
    not g5060(n1590 ,n36[4]);
    nor g5061(n595 ,n17[2] ,n26[2]);
    nand g5062(n5357 ,n5130 ,n5196);
    nand g5063(n4421 ,n21[2] ,n4361);
    nand g5064(n4168 ,n4000 ,n4110);
    nand g5065(n6345 ,n6543 ,n6248);
    buf g5066(n14[15], n11[15]);
    nand g5067(n3873 ,n3668 ,n3819);
    nand g5068(n3726 ,n3585 ,n3607);
    not g5069(n4550 ,n4549);
    nand g5070(n1832 ,n1678 ,n1781);
    nor g5071(n757 ,n593 ,n717);
    dff g5072(.RN(n1), .SN(1'b1), .CK(n0), .D(n1207), .Q(n34[1]));
    or g5073(n3104 ,n6578 ,n6555);
    xnor g5074(n3297 ,n3271 ,n3255);
    nand g5075(n3520 ,n3485 ,n19[4]);
    nand g5076(n3209 ,n3164 ,n3181);
    nand g5077(n5747 ,n5603 ,n5637);
    nand g5078(n4198 ,n4134 ,n4165);
    nand g5079(n4433 ,n21[7] ,n4382);
    xnor g5080(n5605 ,n5444 ,n5281);
    or g5081(n4739 ,n4443 ,n4447);
    xnor g5082(n5163 ,n4935 ,n4551);
    or g5083(n1864 ,n1751 ,n1798);
    nand g5084(n1699 ,n19[7] ,n1650);
    nand g5085(n3237 ,n3204 ,n3236);
    nor g5086(n6255 ,n6231 ,n6252);
    nand g5087(n2775 ,n2662 ,n2729);
    nand g5088(n2018 ,n1980 ,n2001);
    nand g5089(n1251 ,n28[4] ,n1194);
    xnor g5090(n2126 ,n2105 ,n2097);
    nor g5091(n6249 ,n25[0] ,n6224);
    nor g5092(n5401 ,n5123 ,n5290);
    nand g5093(n6141 ,n6127 ,n6065);
    nand g5094(n5576 ,n5335 ,n5486);
    xnor g5095(n4104 ,n4009 ,n3943);
    nand g5096(n4437 ,n4386 ,n20[3]);
    nand g5097(n3602 ,n3462 ,n3478);
    or g5098(n256 ,n229 ,n184);
    not g5099(n120 ,n24[4]);
    nand g5100(n1679 ,n1576 ,n1655);
    xnor g5101(n530 ,n510 ,n516);
    nand g5102(n5072 ,n4744 ,n5009);
    nand g5103(n119 ,n113 ,n118);
    nor g5104(n5838 ,n5655 ,n5791);
    nand g5105(n6389 ,n6266 ,n6313);
    nand g5106(n5105 ,n4841 ,n4962);
    nor g5107(n3689 ,n3619 ,n3612);
    or g5108(n3978 ,n3841 ,n3897);
    nand g5109(n3090 ,n3065 ,n3089);
    xnor g5110(n6502 ,n3069 ,n3075);
    or g5111(n5341 ,n5220 ,n5240);
    xnor g5112(n1782 ,n1636 ,n1730);
    or g5113(n5892 ,n5807 ,n5825);
    or g5114(n3655 ,n3503 ,n3519);
    nor g5115(n712 ,n563 ,n661);
    nand g5116(n2549 ,n2517 ,n2548);
    nand g5117(n2413 ,n2352 ,n2389);
    xnor g5118(n5868 ,n5762 ,n5625);
    nand g5119(n2959 ,n2838 ,n2930);
    nand g5120(n4846 ,n4433 ,n4565);
    nor g5121(n5058 ,n4980 ,n4970);
    xor g5122(n2975 ,n2901 ,n2927);
    nand g5123(n1137 ,n22[3] ,n720);
    nand g5124(n4194 ,n4129 ,n4145);
    nand g5125(n4488 ,n20[7] ,n4367);
    nand g5126(n3233 ,n3203 ,n3232);
    nand g5127(n1844 ,n1818 ,n1799);
    nand g5128(n3166 ,n3119 ,n3142);
    xnor g5129(n5702 ,n5351 ,n5553);
    xnor g5130(n3935 ,n3764 ,n3692);
    nand g5131(n991 ,n19[7] ,n714);
    xnor g5132(n2487 ,n2452 ,n2423);
    nand g5133(n3702 ,n3518 ,n3535);
    nand g5134(n4567 ,n21[1] ,n4388);
    nand g5135(n4588 ,n4389 ,n20[6]);
    or g5136(n4255 ,n4202 ,n4232);
    nand g5137(n4469 ,n21[6] ,n4380);
    nand g5138(n1740 ,n1660 ,n1714);
    nand g5139(n1302 ,n1058 ,n807);
    or g5140(n3657 ,n3512 ,n3536);
    xnor g5141(n5828 ,n5701 ,n5538);
    nand g5142(n2957 ,n2818 ,n2933);
    buf g5143(n14[14], n11[14]);
    xnor g5144(n2368 ,n2302 ,n2309);
    dff g5145(.RN(n1), .SN(1'b1), .CK(n0), .D(n1441), .Q(n12[12]));
    nand g5146(n901 ,n30[6] ,n723);
    nand g5147(n933 ,n29[1] ,n721);
    nand g5148(n3586 ,n3472 ,n3481);
    nor g5149(n2488 ,n2438 ,n2471);
    nand g5150(n3163 ,n3111 ,n3145);
    nor g5151(n6496 ,n2849 ,n2828);
    xnor g5152(n6600 ,n3415 ,n3433);
    or g5153(n5318 ,n5160 ,n5211);
    or g5154(n949 ,n710 ,n664);
    nor g5155(n269 ,n243 ,n206);
    nor g5156(n2678 ,n2568 ,n2619);
    nand g5157(n1286 ,n860 ,n1029);
    nand g5158(n5555 ,n5172 ,n5459);
    nor g5159(n2605 ,n2567 ,n2583);
    or g5160(n414 ,n362 ,n373);
    xnor g5161(n1886 ,n1815 ,n1816);
    dff g5162(.RN(n1), .SN(1'b1), .CK(n0), .D(n1391), .Q(n27[15]));
    dff g5163(.RN(n1), .SN(1'b1), .CK(n0), .D(n1233), .Q(n12[6]));
    nand g5164(n3053 ,n3030 ,n3040);
    not g5165(n4535 ,n4534);
    nand g5166(n4491 ,n4382 ,n20[6]);
    xnor g5167(n5177 ,n4938 ,n4620);
    nand g5168(n5557 ,n5406 ,n5465);
    nand g5169(n1768 ,n1690 ,n1703);
    nand g5170(n3986 ,n3896 ,n3895);
    nand g5171(n5917 ,n5831 ,n5877);
    nand g5172(n6243 ,n41[14] ,n6590);
    nand g5173(n2388 ,n2059 ,n2331);
    nand g5174(n94 ,n74 ,n93);
    nor g5175(n140 ,n32[5] ,n139);
    nand g5176(n4245 ,n4166 ,n4216);
    nor g5177(n5649 ,n5548 ,n5524);
    xnor g5178(n2267 ,n2108 ,n2202);
    nor g5179(n2761 ,n2597 ,n2720);
    nand g5180(n488 ,n451 ,n461);
    not g5181(n132 ,n32[4]);
    nand g5182(n5687 ,n5451 ,n5557);
    xnor g5183(n1645 ,n1631 ,n1615);
    nand g5184(n4566 ,n21[1] ,n4389);
    nor g5185(n4649 ,n4394 ,n4415);
    not g5186(n57 ,n56);
    nor g5187(n2510 ,n2483 ,n2489);
    xnor g5188(n5911 ,n5824 ,n5809);
    nor g5189(n6454 ,n6400 ,n6414);
    nand g5190(n5799 ,n5659 ,n5717);
    nor g5191(n2836 ,n2666 ,n2790);
    nand g5192(n3533 ,n3460 ,n3484);
    xnor g5193(n1876 ,n1645 ,n1813);
    nand g5194(n1664 ,n1582 ,n1652);
    dff g5195(.RN(n1), .SN(1'b1), .CK(n0), .D(n1204), .Q(n34[7]));
    xnor g5196(n6580 ,n2023 ,n2040);
    xnor g5197(n5831 ,n5695 ,n5573);
    not g5198(n4788 ,n4787);
    nand g5199(n661 ,n18[1] ,n558);
    nor g5200(n6254 ,n6227 ,n6223);
    not g5201(n4967 ,n4966);
    xnor g5202(n3744 ,n3520 ,n3597);
    not g5203(n3463 ,n37[4]);
    nand g5204(n988 ,n20[1] ,n714);
    not g5205(n4413 ,n4363);
    nand g5206(n4545 ,n21[4] ,n4371);
    or g5207(n1594 ,n1562 ,n1568);
    xnor g5208(n1779 ,n1636 ,n1723);
    xnor g5209(n5283 ,n4940 ,n4964);
    nor g5210(n5362 ,n5111 ,n5203);
    xnor g5211(n6507 ,n3068 ,n3085);
    buf g5212(n13[1], n10[1]);
    nand g5213(n1424 ,n800 ,n1179);
    nand g5214(n5751 ,n5516 ,n5668);
    xor g5215(n6617 ,n6566 ,n3345);
    buf g5216(n37[5] ,n1505);
    nand g5217(n3400 ,n6550 ,n39[1]);
    nand g5218(n1657 ,n1586 ,n1651);
    xnor g5219(n2399 ,n2328 ,n2292);
    or g5220(n4735 ,n4469 ,n4456);
    nor g5221(n882 ,n614 ,n711);
    nand g5222(n1100 ,n33[3] ,n710);
    nor g5223(n2538 ,n2522 ,n2533);
    not g5224(n5950 ,n5949);
    nand g5225(n3111 ,n38[12] ,n6585);
    nand g5226(n201 ,n159 ,n157);
    not g5227(n3443 ,n3442);
    or g5228(n258 ,n193 ,n217);
    nand g5229(n3099 ,n38[8] ,n6581);
    dff g5230(.RN(n1), .SN(1'b1), .CK(n0), .D(n1205), .Q(n34[5]));
    nand g5231(n4572 ,n20[3] ,n4363);
    nand g5232(n1378 ,n823 ,n1127);
    xnor g5233(n4265 ,n4229 ,n4247);
    nor g5234(n2900 ,n2815 ,n2889);
    xnor g5235(n2868 ,n2772 ,n2674);
    not g5236(n2707 ,n2706);
    nand g5237(n5248 ,n5147 ,n5066);
    xnor g5238(n6595 ,n3215 ,n3233);
    nand g5239(n1005 ,n4[1] ,n557);
    nand g5240(n4587 ,n4388 ,n20[3]);
    nor g5241(n598 ,n23[4] ,n34[4]);
    xnor g5242(n1650 ,n1639 ,n1593);
    nand g5243(n4496 ,n21[0] ,n4382);
    nand g5244(n2104 ,n2071 ,n2084);
    nand g5245(n2210 ,n6541 ,n2148);
    xnor g5246(n1521 ,n519 ,n548);
    not g5247(n4503 ,n4502);
    xnor g5248(n6602 ,n3409 ,n3429);
    xnor g5249(n1952 ,n1797 ,n1918);
    nand g5250(n1336 ,n898 ,n1088);
    nand g5251(n3832 ,n3734 ,n3777);
    or g5252(n5916 ,n5847 ,n5885);
    dff g5253(.RN(n1), .SN(1'b1), .CK(n0), .D(n1467), .Q(n28[4]));
    nand g5254(n3601 ,n3464 ,n3485);
    nand g5255(n1101 ,n20[3] ,n722);
    nand g5256(n6319 ,n39[7] ,n6248);
    xnor g5257(n2528 ,n2487 ,n2447);
    nand g5258(n1474 ,n980 ,n1413);
    nand g5259(n4165 ,n4087 ,n4126);
    not g5260(n3552 ,n3551);
    nand g5261(n623 ,n18[0] ,n18[1]);
    nand g5262(n4520 ,n21[0] ,n4384);
    xnor g5263(n2926 ,n2865 ,n2874);
    or g5264(n2946 ,n2929 ,n2920);
    nand g5265(n2212 ,n6534 ,n2178);
    nand g5266(n5936 ,n5777 ,n4359);
    nand g5267(n4037 ,n3935 ,n3969);
    nor g5268(n2020 ,n1971 ,n1999);
    nand g5269(n2034 ,n2019 ,n2025);
    nor g5270(n4654 ,n4414 ,n4402);
    xnor g5271(n4964 ,n4647 ,n4660);
    not g5272(n4110 ,n4109);
    nand g5273(n4257 ,n4193 ,n4231);
    nor g5274(n4658 ,n4409 ,n4413);
    not g5275(n4381 ,n36[5]);
    xnor g5276(n4324 ,n4299 ,n4275);
    xnor g5277(n5620 ,n5438 ,n5204);
    nor g5278(n2355 ,n2235 ,n2316);
    nor g5279(n112 ,n24[7] ,n111);
    or g5280(n750 ,n711 ,n681);
    xnor g5281(n1544 ,n32[6] ,n141);
    nand g5282(n6348 ,n6504 ,n6249);
    xnor g5283(n4228 ,n4174 ,n4153);
    xnor g5284(n1969 ,n1934 ,n1886);
    nand g5285(n4446 ,n21[7] ,n4363);
    nand g5286(n5016 ,n4533 ,n4837);
    nor g5287(n4020 ,n3914 ,n3997);
    xnor g5288(n665 ,n19[4] ,n27[4]);
    dff g5289(.RN(n1), .SN(1'b1), .CK(n0), .D(n1477), .Q(n17[4]));
    nand g5290(n5516 ,n5206 ,n5457);
    nand g5291(n1738 ,n1579 ,n1675);
    xor g5292(n3747 ,n3566 ,n3536);
    or g5293(n3185 ,n3156 ,n3173);
    nand g5294(n4234 ,n4071 ,n4212);
    xnor g5295(n2443 ,n2058 ,n2407);
    or g5296(n4736 ,n4492 ,n4434);
    or g5297(n4710 ,n4433 ,n4565);
    nand g5298(n5727 ,n5508 ,n5653);
    xor g5299(n6518 ,n6580 ,n6557);
    or g5300(n4711 ,n4611 ,n4597);
    or g5301(n3195 ,n3159 ,n3182);
    dff g5302(.RN(n1), .SN(1'b1), .CK(n0), .D(n1298), .Q(n11[7]));
    not g5303(n1581 ,n36[5]);
    nand g5304(n960 ,n33[3] ,n554);
    xnor g5305(n6504 ,n3067 ,n3079);
    nand g5306(n388 ,n261 ,n349);
    nand g5307(n2940 ,n2813 ,n2904);
    xnor g5308(n6197 ,n6165 ,n6183);
    nand g5309(n1135 ,n20[5] ,n722);
    nand g5310(n1205 ,n814 ,n733);
    nand g5311(n4078 ,n3980 ,n4039);
    nand g5312(n5934 ,n5851 ,n5881);
    or g5313(n5918 ,n5831 ,n5877);
    xnor g5314(n4343 ,n4316 ,n4325);
    dff g5315(.RN(n1), .SN(1'b1), .CK(n0), .D(n1453), .Q(n33[1]));
    xnor g5316(n2304 ,n2235 ,n2237);
    nand g5317(n5449 ,n5343 ,n5353);
    or g5318(n262 ,n178 ,n215);
    nand g5319(n4662 ,n4384 ,n20[0]);
    xnor g5320(n1932 ,n1874 ,n1799);
    nand g5321(n1034 ,n2[7] ,n713);
    nand g5322(n3825 ,n3639 ,n3702);
    xnor g5323(n670 ,n35[14] ,n33[14]);
    nand g5324(n3636 ,n3481 ,n19[6]);
    xnor g5325(n2009 ,n1984 ,n1954);
    xnor g5326(n5286 ,n4941 ,n4520);
    nor g5327(n2651 ,n2565 ,n2596);
    nand g5328(n4625 ,n4388 ,n20[0]);
    xor g5329(n693 ,n26[0] ,n17[0]);
    nand g5330(n1050 ,n11[9] ,n710);
    dff g5331(.RN(n1), .SN(1'b1), .CK(n0), .D(n1417), .Q(n20[2]));
    xnor g5332(n1815 ,n1646 ,n1741);
    nand g5333(n3622 ,n3470 ,n3486);
    nand g5334(n928 ,n33[2] ,n712);
    not g5335(n1885 ,n1884);
    nor g5336(n1963 ,n1902 ,n1940);
    not g5337(n3256 ,n37[6]);
    xnor g5338(n6029 ,n5962 ,n5973);
    buf g5339(n14[13], n11[13]);
    nand g5340(n6275 ,n6531 ,n6250);
    nand g5341(n5995 ,n5896 ,n5941);
    nand g5342(n4827 ,n4463 ,n4446);
    nand g5343(n454 ,n400 ,n442);
    nor g5344(n2500 ,n2465 ,n2479);
    nand g5345(n6367 ,n6577 ,n6247);
    nor g5346(n3353 ,n3318 ,n3352);
    nand g5347(n6018 ,n5922 ,n5983);
    nand g5348(n810 ,n35[1] ,n554);
    or g5349(n2045 ,n2026 ,n2044);
    xnor g5350(n88 ,n67 ,n49);
    nor g5351(n2634 ,n2568 ,n2588);
    xnor g5352(n3410 ,n6548 ,n6563);
    not g5353(n4681 ,n4680);
    xor g5354(n6565 ,n5153 ,n4625);
    xnor g5355(n4140 ,n4070 ,n3970);
    nand g5356(n3384 ,n3327 ,n3383);
    nand g5357(n4432 ,n20[3] ,n4361);
    not g5358(n4779 ,n4778);
    nor g5359(n6458 ,n6405 ,n6396);
    nor g5360(n4538 ,n4400 ,n4416);
    nand g5361(n4321 ,n4286 ,n4309);
    xnor g5362(n4972 ,n4682 ,n4593);
    nand g5363(n552 ,n492 ,n551);
    xnor g5364(n3763 ,n3598 ,n3593);
    nand g5365(n2502 ,n2445 ,n2469);
    or g5366(n3980 ,n3860 ,n3941);
    nand g5367(n401 ,n350 ,n365);
    nand g5368(n4471 ,n4378 ,n20[5]);
    nand g5369(n4596 ,n20[3] ,n4374);
    nand g5370(n228 ,n169 ,n155);
    dff g5371(.RN(n1), .SN(1'b1), .CK(n0), .D(n1334), .Q(n24[6]));
    nand g5372(n1794 ,n1645 ,n1755);
    nand g5373(n3207 ,n3167 ,n3169);
    dff g5374(.RN(n1), .SN(1'b1), .CK(n0), .D(n1470), .Q(n28[0]));
    nand g5375(n3625 ,n3468 ,n3482);
    nand g5376(n5965 ,n5883 ,n5917);
    nand g5377(n1177 ,n29[5] ,n724);
    nand g5378(n6266 ,n40[14] ,n6250);
    nand g5379(n4357 ,n4282 ,n4356);
    nand g5380(n3961 ,n3854 ,n3919);
    nand g5381(n4258 ,n4211 ,n4244);
    xnor g5382(n305 ,n223 ,n211);
    xnor g5383(n1875 ,n1774 ,n1823);
    nand g5384(n4319 ,n4294 ,n4308);
    nand g5385(n4311 ,n4257 ,n4291);
    nand g5386(n4339 ,n4312 ,n4331);
    nand g5387(n702 ,n587 ,n583);
    dff g5388(.RN(n1), .SN(1'b1), .CK(n0), .D(n1421), .Q(n20[1]));
    not g5389(n3738 ,n3721);
    nand g5390(n3449 ,n3445 ,n19[0]);
    nand g5391(n4354 ,n4328 ,n4353);
    nand g5392(n2337 ,n2308 ,n2290);
    nor g5393(n2724 ,n2566 ,n2630);
    xnor g5394(n5310 ,n5118 ,n5144);
    nand g5395(n2559 ,n2558 ,n2537);
    nand g5396(n5793 ,n5632 ,n5751);
    nor g5397(n2327 ,n2324 ,n2299);
    or g5398(n5938 ,n5802 ,n5875);
    nand g5399(n3082 ,n3047 ,n3081);
    dff g5400(.RN(n1), .SN(1'b1), .CK(n0), .D(n1299), .Q(n1508));
    nand g5401(n5147 ,n4772 ,n4975);
    nand g5402(n4802 ,n4629 ,n4424);
    nand g5403(n1688 ,n1582 ,n1655);
    not g5404(n4112 ,n4111);
    nor g5405(n338 ,n267 ,n313);
    nand g5406(n2252 ,n2165 ,n2189);
    nand g5407(n1306 ,n1064 ,n811);
    xnor g5408(n2317 ,n2119 ,n2256);
    nand g5409(n6396 ,n6272 ,n6316);
    nand g5410(n2219 ,n6540 ,n2148);
    xor g5411(n1642 ,n1628 ,n1605);
    nand g5412(n6407 ,n6335 ,n6356);
    xnor g5413(n3772 ,n3609 ,n3602);
    nand g5414(n3870 ,n3674 ,n3812);
    xnor g5415(n5173 ,n4947 ,n4479);
    xnor g5416(n3036 ,n3005 ,n2969);
    xnor g5417(n5627 ,n5422 ,n5178);
    nor g5418(n2816 ,n2665 ,n2791);
    nand g5419(n6074 ,n5993 ,n6043);
    not g5420(n2503 ,n2502);
    or g5421(n5340 ,n5292 ,n5247);
    xnor g5422(n38[11] ,n2543 ,n2555);
    or g5423(n4724 ,n4428 ,n4438);
    xnor g5424(n4231 ,n4176 ,n4186);
    xnor g5425(n370 ,n301 ,n227);
    xnor g5426(n6065 ,n5998 ,n5929);
    dff g5427(.RN(n1), .SN(1'b1), .CK(n0), .D(n1475), .Q(n29[7]));
    nand g5428(n5574 ,n5337 ,n5487);
    xnor g5429(n3831 ,n3605 ,n3690);
    nand g5430(n3719 ,n3597 ,n3520);
    not g5431(n5575 ,n5574);
    xnor g5432(n5537 ,n5303 ,n5126);
    or g5433(n4750 ,n4497 ,n4578);
    nand g5434(n4551 ,n4388 ,n20[2]);
    xnor g5435(n5817 ,n5631 ,n5752);
    nand g5436(n990 ,n16[7] ,n714);
    xnor g5437(n376 ,n312 ,n267);
    xor g5438(n3765 ,n3635 ,n3537);
    or g5439(n5244 ,n4784 ,n5084);
    xnor g5440(n2366 ,n2287 ,n2289);
    nand g5441(n6201 ,n6167 ,n6193);
    nand g5442(n1223 ,n943 ,n741);
    xnor g5443(n5625 ,n5417 ,n5216);
    nand g5444(n2110 ,n2077 ,n2103);
    nand g5445(n4811 ,n4564 ,n4485);
    or g5446(n3651 ,n3604 ,n3511);
    nand g5447(n5368 ,n5095 ,n5274);
    nand g5448(n4130 ,n3999 ,n4064);
    nand g5449(n2386 ,n2272 ,n2356);
    nand g5450(n6170 ,n6156 ,n6141);
    dff g5451(.RN(n1), .SN(1'b1), .CK(n0), .D(n1319), .Q(n34[14]));
    xnor g5452(n5768 ,n5610 ,n5568);
    nand g5453(n4438 ,n20[6] ,n4371);
    or g5454(n2818 ,n2797 ,n2761);
    nand g5455(n3108 ,n38[14] ,n6587);
    xnor g5456(n5523 ,n5315 ,n5076);
    xnor g5457(n1830 ,n1648 ,n1756);
    xnor g5458(n5428 ,n5188 ,n5082);
    nand g5459(n3060 ,n3027 ,n3036);
    xnor g5460(n5457 ,n5154 ,n4785);
    nand g5461(n4356 ,n4355 ,n4321);
    nor g5462(n4505 ,n4412 ,n4406);
    nand g5463(n5070 ,n4718 ,n4994);
    nand g5464(n5984 ,n5906 ,n5928);
    not g5465(n3868 ,n3867);
    nand g5466(n4992 ,n4537 ,n4798);
    nand g5467(n818 ,n23[5] ,n715);
    not g5468(n4024 ,n4023);
    xnor g5469(n4205 ,n4142 ,n4086);
    xnor g5470(n465 ,n428 ,n404);
    xnor g5471(n5161 ,n4933 ,n4684);
    nand g5472(n1428 ,n993 ,n1184);
    nand g5473(n2589 ,n40[5] ,n6516);
    buf g5474(n15[0], n15[4]);
    xnor g5475(n4269 ,n4225 ,n4205);
    nand g5476(n5385 ,n5285 ,n5190);
    nand g5477(n4275 ,n4215 ,n4254);
    nand g5478(n3708 ,n3588 ,n3506);
    not g5479(n419 ,n418);
    nand g5480(n6287 ,n6568 ,n6254);
    xnor g5481(n41[14] ,n6175 ,n6219);
    nand g5482(n5731 ,n5534 ,n5633);
    nand g5483(n4424 ,n20[0] ,n4369);
    nor g5484(n6478 ,n6427 ,n6426);
    nand g5485(n3381 ,n3334 ,n3380);
    nand g5486(n3198 ,n3156 ,n3173);
    nand g5487(n5719 ,n5543 ,n5614);
    or g5488(n3095 ,n38[9] ,n6582);
    xnor g5489(n3909 ,n3768 ,n3524);
    or g5490(n5999 ,n5931 ,n5971);
    xnor g5491(n5957 ,n5874 ,n5828);
    nor g5492(n622 ,n17[2] ,n17[3]);
    not g5493(n165 ,n164);
    nand g5494(n1685 ,n1584 ,n1655);
    nand g5495(n5102 ,n4730 ,n4990);
    not g5496(n5078 ,n5077);
    nand g5497(n963 ,n27[10] ,n715);
    or g5498(n2570 ,n40[9] ,n6520);
    nand g5499(n1059 ,n27[15] ,n718);
    nand g5500(n35[0] ,n6452 ,n6450);
    nor g5501(n4661 ,n4397 ,n4390);
    nor g5502(n2650 ,n2565 ,n2590);
    nand g5503(n1845 ,n1830 ,n1812);
    nand g5504(n6355 ,n38[3] ,n6246);
    xor g5505(n4887 ,n4699 ,n4628);
    not g5506(n4416 ,n4361);
    nand g5507(n35[2] ,n6460 ,n6459);
    nand g5508(n3875 ,n3657 ,n3818);
    or g5509(n4752 ,n4457 ,n4450);
    xnor g5510(n41[13] ,n6197 ,n6217);
    nand g5511(n5030 ,n4509 ,n4831);
    xor g5512(n4012 ,n3905 ,n3913);
    nand g5513(n4461 ,n4378 ,n20[1]);
    nand g5514(n243 ,n169 ,n157);
    xor g5515(n3756 ,n3618 ,n3590);
    nand g5516(n1138 ,n33[8] ,n711);
    xnor g5517(n2956 ,n2895 ,n2733);
    nand g5518(n5356 ,n5090 ,n5235);
    nand g5519(n5134 ,n4729 ,n5006);
    nand g5520(n2891 ,n2776 ,n2848);
    xnor g5521(n4270 ,n4224 ,n4233);
    nand g5522(n2475 ,n2429 ,n2453);
    not g5523(n1577 ,n1590);
    nor g5524(n1888 ,n1810 ,n1839);
    nor g5525(n3561 ,n3492 ,n3495);
    buf g5526(n37[4] ,n1504);
    nand g5527(n4447 ,n20[4] ,n4373);
    xnor g5528(n320 ,n213 ,n214);
    not g5529(n2522 ,n2521);
    nand g5530(n942 ,n24[1] ,n715);
    nor g5531(n3791 ,n3576 ,n3688);
    xnor g5532(n6025 ,n5964 ,n5857);
    xnor g5533(n6575 ,n1877 ,n1832);
    xnor g5534(n4060 ,n3955 ,n3898);
    nand g5535(n1207 ,n831 ,n787);
    not g5536(n48 ,n37[5]);
    nand g5537(n3152 ,n3108 ,n3138);
    nor g5538(n2360 ,n2282 ,n2321);
    xor g5539(n1651 ,n1633 ,n1640);
    nand g5540(n5133 ,n4761 ,n5003);
    dff g5541(.RN(n1), .SN(1'b1), .CK(n0), .D(n1220), .Q(n28[5]));
    nand g5542(n3588 ,n3460 ,n3476);
    dff g5543(.RN(n1), .SN(1'b1), .CK(n0), .D(n1463), .Q(n22[6]));
    nand g5544(n1934 ,n1897 ,n1911);
    not g5545(n89 ,n88);
    nand g5546(n4799 ,n4636 ,n4452);
    xnor g5547(n1821 ,n1645 ,n1755);
    or g5548(n5886 ,n5622 ,n5833);
    nand g5549(n5590 ,n5370 ,n5478);
    xnor g5550(n3779 ,n3616 ,n3640);
    nand g5551(n4216 ,n4147 ,n4201);
    not g5552(n4687 ,n4686);
    nand g5553(n5096 ,n4755 ,n5029);
    xnor g5554(n3024 ,n2972 ,n2953);
    dff g5555(.RN(n1), .SN(1'b1), .CK(n0), .D(n1449), .Q(n34[6]));
    not g5556(n158 ,n36[7]);
    nor g5557(n835 ,n560 ,n721);
    xnor g5558(n1654 ,n1635 ,n1625);
    xor g5559(n5438 ,n5201 ,n5214);
    xnor g5560(n2022 ,n2003 ,n1994);
    or g5561(n5322 ,n5185 ,n5183);
    or g5562(n4722 ,n4605 ,n4599);
    nand g5563(n1215 ,n918 ,n763);
    nand g5564(n3073 ,n3046 ,n3057);
    xnor g5565(n5154 ,n4970 ,n4612);
    xnor g5566(n4223 ,n4105 ,n4199);
    nand g5567(n4331 ,n4279 ,n4317);
    not g5568(n1570 ,n1569);
    dff g5569(.RN(n1), .SN(1'b1), .CK(n0), .D(n1367), .Q(n23[5]));
    nand g5570(n4831 ,n4448 ,n4589);
    nand g5571(n5082 ,n4713 ,n4998);
    nand g5572(n3138 ,n6564 ,n3094);
    nor g5573(n2782 ,n2636 ,n2711);
    not g5574(n64 ,n36[3]);
    xnor g5575(n5607 ,n5440 ,n5286);
    not g5576(n3274 ,n36[6]);
    or g5577(n481 ,n441 ,n464);
    xnor g5578(n3344 ,n6568 ,n6576);
    nand g5579(n4462 ,n20[4] ,n4365);
    or g5580(n4770 ,n4569 ,n4601);
    not g5581(n5628 ,n5627);
    xnor g5582(n4232 ,n4179 ,n4083);
    xnor g5583(n3215 ,n3167 ,n3169);
    dff g5584(.RN(n1), .SN(1'b1), .CK(n0), .D(n1285), .Q(n11[15]));
    or g5585(n5652 ,n5491 ,n5570);
    not g5586(n1780 ,n1779);
    nand g5587(n2173 ,n6540 ,n2127);
    xnor g5588(n2370 ,n2260 ,n2314);
    xnor g5589(n6612 ,n3365 ,n41[6]);
    nand g5590(n4041 ,n3874 ,n3983);
    xnor g5591(n3005 ,n2951 ,n2917);
    nand g5592(n910 ,n23[9] ,n715);
    nand g5593(n379 ,n219 ,n343);
    buf g5594(n13[10], n10[10]);
    not g5595(n2513 ,n2512);
    not g5596(n4783 ,n4782);
    or g5597(n251 ,n183 ,n212);
    nand g5598(n2591 ,n40[6] ,n6517);
    xnor g5599(n5876 ,n5759 ,n5541);
    or g5600(n3192 ,n3164 ,n3181);
    nand g5601(n5669 ,n5471 ,n5590);
    or g5602(n5342 ,n5280 ,n5158);
    not g5603(n2659 ,n2658);
    nor g5604(n2338 ,n2308 ,n2290);
    xor g5605(n3757 ,n3626 ,n3594);
    not g5606(n5533 ,n5532);
    nand g5607(n3812 ,n3637 ,n3729);
    not g5608(n3686 ,n3685);
    nor g5609(n2390 ,n2319 ,n2329);
    nand g5610(n2348 ,n2296 ,n2291);
    nand g5611(n1429 ,n994 ,n1187);
    xnor g5612(n3415 ,n6545 ,n6560);
    nand g5613(n1158 ,n23[9] ,n716);
    nand g5614(n4450 ,n20[7] ,n4363);
    nand g5615(n3834 ,n3686 ,n3782);
    xnor g5616(n2533 ,n2486 ,n2464);
    nor g5617(n6468 ,n6442 ,n6440);
    not g5618(n1869 ,n1852);
    nand g5619(n4810 ,n4567 ,n4590);
    nand g5620(n1663 ,n1577 ,n1651);
    xnor g5621(n6592 ,n3222 ,n3247);
    not g5622(n3555 ,n3554);
    nor g5623(n2322 ,n2269 ,n2281);
    not g5624(n5408 ,n5386);
    xnor g5625(n4916 ,n4501 ,n4573);
    nand g5626(n1127 ,n1533 ,n716);
    nand g5627(n1201 ,n603 ,n795);
    xnor g5628(n6598 ,n3407 ,n3437);
    dff g5629(.RN(n1), .SN(1'b1), .CK(n0), .D(n1358), .Q(n32[3]));
    not g5630(n5169 ,n5168);
    nand g5631(n1479 ,n825 ,n1248);
    nand g5632(n5816 ,n5682 ,n5727);
    nand g5633(n4244 ,n4185 ,n4210);
    xnor g5634(n2032 ,n2013 ,n2005);
    nor g5635(n2602 ,n2567 ,n2590);
    nor g5636(n3422 ,n3413 ,n3421);
    nor g5637(n3287 ,n3271 ,n3255);
    nand g5638(n5054 ,n4659 ,n4829);
    dff g5639(.RN(n1), .SN(1'b1), .CK(n0), .D(n1282), .Q(n1515));
    nand g5640(n3305 ,n3289 ,n3299);
    nand g5641(n5994 ,n5898 ,n5948);
    nor g5642(n330 ,n233 ,n294);
    nand g5643(n6433 ,n6296 ,n6367);
    nor g5644(n2889 ,n2768 ,n2832);
    nand g5645(n2595 ,n40[12] ,n6523);
    xnor g5646(n5213 ,n4928 ,n4458);
    nand g5647(n6420 ,n6382 ,n6349);
    not g5648(n2178 ,n2177);
    xnor g5649(n5180 ,n4937 ,n4534);
    nand g5650(n2777 ,n2671 ,n2739);
    nand g5651(n5660 ,n5550 ,n5537);
    nand g5652(n4591 ,n20[6] ,n4369);
    buf g5653(n13[13], n10[13]);
    nor g5654(n3959 ,n3901 ,n3936);
    not g5655(n6035 ,n6034);
    dff g5656(.RN(n1), .SN(1'b1), .CK(n0), .D(n1464), .Q(n22[5]));
    nand g5657(n2141 ,n6534 ,n2121);
    nand g5658(n5249 ,n5092 ,n5065);
    xnor g5659(n3212 ,n3173 ,n3156);
    nand g5660(n1408 ,n972 ,n1164);
    not g5661(n5617 ,n5616);
    dff g5662(.RN(n1), .SN(1'b1), .CK(n0), .D(n1203), .Q(n17[1]));
    nand g5663(n2732 ,n6527 ,n2624);
    nor g5664(n2992 ,n2917 ,n2952);
    nand g5665(n4128 ,n3892 ,n4056);
    dff g5666(.RN(n1), .SN(1'b1), .CK(n0), .D(n1437), .Q(n29[3]));
    not g5667(n3465 ,n37[5]);
    nand g5668(n2156 ,n6540 ,n2123);
    nor g5669(n441 ,n340 ,n397);
    nand g5670(n2111 ,n2087 ,n2102);
    not g5671(n4683 ,n4682);
    nand g5672(n4857 ,n4625 ,n4441);
    nand g5673(n5858 ,n5736 ,n5796);
    nand g5674(n3230 ,n3187 ,n3229);
    dff g5675(.RN(n1), .SN(1'b1), .CK(n0), .D(n1257), .Q(n16[5]));
    not g5676(n1649 ,n1650);
    nor g5677(n573 ,n17[4] ,n26[4]);
    nand g5678(n4308 ,n4278 ,n4290);
    nand g5679(n4452 ,n4380 ,n20[4]);
    buf g5680(n13[7], n11[7]);
    xnor g5681(n6501 ,n3050 ,n3073);
    or g5682(n4182 ,n4079 ,n4153);
    nand g5683(n5361 ,n5088 ,n5237);
    not g5684(n5604 ,n5603);
    not g5685(n292 ,n281);
    nand g5686(n6422 ,n6295 ,n6343);
    nand g5687(n1442 ,n1009 ,n1263);
    nand g5688(n3584 ,n3464 ,n3476);
    nand g5689(n3995 ,n3864 ,n3894);
    nand g5690(n2170 ,n6535 ,n2126);
    not g5691(n3974 ,n3973);
    nand g5692(n644 ,n22[6] ,n26[6]);
    nand g5693(n6072 ,n5994 ,n6048);
    nor g5694(n2726 ,n2568 ,n2631);
    xnor g5695(n4322 ,n4309 ,n4286);
    nand g5696(n4840 ,n4570 ,n4603);
    nor g5697(n6550 ,n3740 ,n3681);
    not g5698(n2236 ,n2235);
    xnor g5699(n1781 ,n1637 ,n1727);
    dff g5700(.RN(n1), .SN(1'b1), .CK(n0), .D(n1302), .Q(n11[4]));
    nand g5701(n4548 ,n21[0] ,n4388);
    nand g5702(n1280 ,n857 ,n1031);
    or g5703(n2581 ,n40[8] ,n6519);
    nand g5704(n1168 ,n5[6] ,n713);
    dff g5705(.RN(n1), .SN(1'b1), .CK(n0), .D(n1225), .Q(n27[5]));
    nand g5706(n4576 ,n20[4] ,n4369);
    nand g5707(n1273 ,n853 ,n1023);
    not g5708(n3259 ,n3258);
    nand g5709(n5022 ,n4508 ,n4847);
    nor g5710(n2644 ,n2566 ,n2593);
    nand g5711(n1260 ,n631 ,n882);
    nor g5712(n718 ,n18[2] ,n661);
    xnor g5713(n5435 ,n5196 ,n5143);
    xnor g5714(n4970 ,n4504 ,n4543);
    nor g5715(n767 ,n609 ,n720);
    xnor g5716(n5212 ,n4915 ,n4605);
    dff g5717(.RN(n1), .SN(1'b1), .CK(n0), .D(n1304), .Q(n11[2]));
    xor g5718(n3761 ,n3617 ,n3532);
    nand g5719(n4635 ,n20[2] ,n4361);
    xnor g5720(n3936 ,n3756 ,n3528);
    nand g5721(n402 ,n265 ,n359);
    dff g5722(.RN(n1), .SN(1'b1), .CK(n0), .D(n1425), .Q(n26[2]));
    nor g5723(n1973 ,n1939 ,n1950);
    nand g5724(n2846 ,n2786 ,n2760);
    xnor g5725(n683 ,n35[3] ,n31[3]);
    nor g5726(n353 ,n250 ,n330);
    nor g5727(n776 ,n598 ,n717);
    xnor g5728(n4966 ,n4548 ,n4664);
    nand g5729(n185 ,n170 ,n157);
    nand g5730(n4631 ,n21[1] ,n4386);
    not g5731(n4108 ,n4107);
    nand g5732(n5710 ,n5533 ,n5625);
    not g5733(n5804 ,n5803);
    nand g5734(n100 ,n78 ,n99);
    nand g5735(n3007 ,n2962 ,n2979);
    nor g5736(n235 ,n177 ,n174);
    or g5737(n5470 ,n5216 ,n5411);
    nand g5738(n6172 ,n6121 ,n6145);
    xnor g5739(n5431 ,n5292 ,n5134);
    nor g5740(n264 ,n195 ,n234);
    nand g5741(n5681 ,n5501 ,n5531);
    nand g5742(n1852 ,n1819 ,n1800);
    nor g5743(n3399 ,n6554 ,n39[5]);
    xnor g5744(n6584 ,n2038 ,n2048);
    xnor g5745(n5517 ,n5306 ,n5077);
    nand g5746(n5668 ,n5511 ,n5589);
    xnor g5747(n5915 ,n5823 ,n5813);
    xnor g5748(n1546 ,n32[4] ,n138);
    nand g5749(n2908 ,n2822 ,n2892);
    xnor g5750(n1801 ,n1648 ,n1744);
    not g5751(n5116 ,n5115);
    xnor g5752(n2873 ,n2708 ,n2802);
    xnor g5753(n3006 ,n2948 ,n2924);
    nand g5754(n2617 ,n2588 ,n2569);
    not g5755(n3491 ,n3484);
    nand g5756(n2258 ,n2175 ,n2219);
    nand g5757(n3710 ,n3521 ,n3589);
    not g5758(n1485 ,n1484);
    nand g5759(n5550 ,n5331 ,n5468);
    xnor g5760(n311 ,n195 ,n234);
    nand g5761(n5738 ,n5574 ,n5628);
    nand g5762(n3877 ,n3658 ,n3808);
    nand g5763(n6077 ,n5969 ,n6051);
    nand g5764(n5091 ,n4740 ,n5031);
    nand g5765(n5029 ,n4540 ,n4827);
    or g5766(n5513 ,n5404 ,n5493);
    not g5767(n174 ,n37[7]);
    nand g5768(n3701 ,n3533 ,n3581);
    nand g5769(n3844 ,n3653 ,n3797);
    xnor g5770(n3752 ,n3521 ,n3589);
    nor g5771(n2793 ,n2603 ,n2701);
    xnor g5772(n5188 ,n4943 ,n4637);
    nand g5773(n4439 ,n21[2] ,n4388);
    or g5774(n4755 ,n4463 ,n4446);
    or g5775(n4761 ,n4627 ,n4634);
    nand g5776(n1437 ,n931 ,n1211);
    nand g5777(n3633 ,n3486 ,n19[5]);
    xor g5778(n5700 ,n5571 ,n5582);
    xnor g5779(n6003 ,n5914 ,n5854);
    not g5780(n2566 ,n6529);
    nand g5781(n3703 ,n3578 ,n3540);
    nand g5782(n3725 ,n3501 ,n3591);
    xnor g5783(n4025 ,n3915 ,n3869);
    nand g5784(n1481 ,n724 ,n1200);
    dff g5785(.RN(n1), .SN(1'b1), .CK(n0), .D(n1332), .Q(n24[7]));
    nor g5786(n4650 ,n4392 ,n4404);
    nor g5787(n2136 ,n2060 ,n2124);
    nand g5788(n5077 ,n4752 ,n5028);
    not g5789(n2492 ,n2491);
    xnor g5790(n1813 ,n1761 ,n1646);
    nand g5791(n1267 ,n645 ,n877);
    nand g5792(n4033 ,n3942 ,n3986);
    nand g5793(n1014 ,n3[6] ,n557);
    or g5794(n3658 ,n3587 ,n3592);
    nand g5795(n4314 ,n4272 ,n4303);
    nand g5796(n6206 ,n6195 ,n6184);
    nand g5797(n381 ,n275 ,n354);
    xnor g5798(n2450 ,n2305 ,n2410);
    xnor g5799(n5441 ,n5157 ,n5127);
    nand g5800(n1957 ,n1914 ,n1936);
    nand g5801(n458 ,n396 ,n440);
    nor g5802(n5240 ,n5069 ,n5075);
    nand g5803(n3380 ,n3321 ,n3379);
    nand g5804(n3582 ,n3482 ,n19[3]);
    nand g5805(n5375 ,n5100 ,n5245);
    nand g5806(n1352 ,n900 ,n1105);
    xnor g5807(n5616 ,n5415 ,n5223);
    nand g5808(n6297 ,n41[13] ,n6254);
    not g5809(n2550 ,n2549);
    nand g5810(n841 ,n16[6] ,n714);
    nor g5811(n2671 ,n2568 ,n2594);
    nor g5812(n2553 ,n2520 ,n2552);
    nand g5813(n1337 ,n899 ,n1089);
    xnor g5814(n2080 ,n21[6] ,n20[6]);
    nand g5815(n3993 ,n3879 ,n3930);
    xnor g5816(n1988 ,n1956 ,n1923);
    nand g5817(n5486 ,n5140 ,n5397);
    xnor g5818(n429 ,n377 ,n344);
    not g5819(n2746 ,n2745);
    not g5820(n65 ,n64);
    xnor g5821(n1807 ,n1648 ,n1762);
    xnor g5822(n6067 ,n5997 ,n5930);
    xnor g5823(n5538 ,n5309 ,n5091);
    nor g5824(n2672 ,n2568 ,n2582);
    xor g5825(n6528 ,n3453 ,n3449);
    xnor g5826(n3917 ,n3782 ,n3685);
    xnor g5827(n3771 ,n3508 ,n3507);
    nor g5828(n3956 ,n3891 ,n3904);
    nor g5829(n2551 ,n2550 ,n2516);
    nand g5830(n1380 ,n647 ,n884);
    nand g5831(n5269 ,n5137 ,n5126);
    nand g5832(n1240 ,n1100 ,n749);
    nand g5833(n5494 ,n5256 ,n5345);
    or g5834(n5475 ,n5223 ,n5407);
    nand g5835(n4492 ,n4384 ,n20[2]);
    nand g5836(n4982 ,n4699 ,n4860);
    not g5837(n3740 ,n3727);
    nand g5838(n6440 ,n6300 ,n6371);
    not g5839(n3304 ,n3303);
    dff g5840(.RN(n1), .SN(1'b1), .CK(n0), .D(n1406), .Q(n21[1]));
    not g5841(n1913 ,n1912);
    xnor g5842(n6539 ,n3296 ,n3314);
    not g5843(n5630 ,n5629);
    or g5844(n3047 ,n3007 ,n3025);
    or g5845(n2812 ,n2781 ,n2755);
    dff g5846(.RN(n1), .SN(1'b1), .CK(n0), .D(n1402), .Q(n21[3]));
    xnor g5847(n3222 ,n3159 ,n3182);
    nand g5848(n539 ,n524 ,n535);
    not g5849(n4403 ,n4373);
    nand g5850(n526 ,n500 ,n518);
    nor g5851(n584 ,n26[1] ,n26[2]);
    nand g5852(n1254 ,n840 ,n997);
    dff g5853(.RN(n1), .SN(1'b1), .CK(n0), .D(n1423), .Q(n20[0]));
    nor g5854(n4546 ,n4414 ,n4401);
    nand g5855(n5268 ,n5136 ,n5124);
    xnor g5856(n2289 ,n2221 ,n2120);
    nand g5857(n1261 ,n845 ,n1005);
    nand g5858(n1452 ,n1128 ,n1348);
    nand g5859(n5684 ,n5491 ,n5570);
    or g5860(n728 ,n555 ,n682);
    xor g5861(n40[0] ,n38[1] ,n39[0]);
    nand g5862(n35[3] ,n6478 ,n6447);
    or g5863(n6058 ,n5969 ,n6051);
    nand g5864(n6119 ,n6053 ,n6092);
    xnor g5865(n686 ,n35[6] ,n31[6]);
    nand g5866(n3200 ,n3159 ,n3182);
    nor g5867(n1978 ,n1917 ,n1948);
    xnor g5868(n2270 ,n2119 ,n2210);
    nand g5869(n324 ,n198 ,n273);
    nand g5870(n628 ,n23[6] ,n34[6]);
    or g5871(n3041 ,n3019 ,n3023);
    nor g5872(n5666 ,n5518 ,n5544);
    nand g5873(n3608 ,n3462 ,n3485);
    nand g5874(n6321 ,n6580 ,n6247);
    nor g5875(n1676 ,n1642 ,n1651);
    nand g5876(n2963 ,n2915 ,n2921);
    nor g5877(n4046 ,n3788 ,n3992);
    nand g5878(n1389 ,n653 ,n780);
    nand g5879(n453 ,n388 ,n430);
    xnor g5880(n5874 ,n5770 ,n5810);
    nor g5881(n267 ,n242 ,n246);
    xor g5882(n5222 ,n4906 ,n4469);
    not g5883(n1192 ,n1131);
    dff g5884(.RN(n1), .SN(1'b1), .CK(n0), .D(n1352), .Q(n23[11]));
    nor g5885(n3642 ,n3492 ,n3499);
    nand g5886(n2166 ,n6538 ,n2126);
    not g5887(n50 ,n37[2]);
    nand g5888(n6264 ,n41[14] ,n6254);
    nand g5889(n964 ,n21[4] ,n714);
    nor g5890(n2404 ,n2392 ,n2364);
    xnor g5891(n5722 ,n5510 ,n5350);
    xnor g5892(n5166 ,n4879 ,n4532);
    xnor g5893(n5426 ,n5194 ,n5089);
    nor g5894(n762 ,n605 ,n723);
    xnor g5895(n3402 ,n6546 ,n6561);
    nand g5896(n651 ,n21[6] ,n30[6]);
    nand g5897(n3247 ,n3209 ,n3246);
    not g5898(n4420 ,n4419);
    or g5899(n5274 ,n5136 ,n5124);
    xnor g5900(n368 ,n320 ,n239);
    nand g5901(n2280 ,n2234 ,n2232);
    nand g5902(n3800 ,n3627 ,n3700);
    not g5903(n3283 ,n3282);
    nand g5904(n891 ,n33[5] ,n554);
    xnor g5905(n3302 ,n3285 ,n3263);
    not g5906(n3557 ,n3556);
    nand g5907(n3545 ,n3481 ,n19[1]);
    nand g5908(n6428 ,n6292 ,n6358);
    not g5909(n61 ,n60);
    nand g5910(n3293 ,n3279 ,n3261);
    dff g5911(.RN(n1), .SN(1'b1), .CK(n0), .D(n1476), .Q(n17[7]));
    nand g5912(n2446 ,n2377 ,n2422);
    nand g5913(n6392 ,n6268 ,n6319);
    nand g5914(n3598 ,n3472 ,n3476);
    xnor g5915(n5434 ,n5221 ,n5119);
    not g5916(n72 ,n36[2]);
    xnor g5917(n3891 ,n3765 ,n3530);
    nand g5918(n2167 ,n6534 ,n2126);
    nand g5919(n1198 ,n740 ,n736);
    nand g5920(n4821 ,n4638 ,n4576);
    nand g5921(n5089 ,n4720 ,n5008);
    or g5922(n1859 ,n1803 ,n1804);
    nand g5923(n5752 ,n5558 ,n5686);
    nand g5924(n3241 ,n3199 ,n3240);
    nand g5925(n3579 ,n3466 ,n3485);
    xnor g5926(n5055 ,n4583 ,n4782);
    nor g5927(n3429 ,n3393 ,n3428);
    or g5928(n4188 ,n4155 ,n4160);
    not g5929(n4392 ,n4382);
    xnor g5930(n6092 ,n6021 ,n5974);
    nor g5931(n2599 ,n2567 ,n2589);
    not g5932(n87 ,n86);
    nand g5933(n3580 ,n3481 ,n19[0]);
    not g5934(n3301 ,n3300);
    dff g5935(.RN(n1), .SN(1'b1), .CK(n0), .D(n1344), .Q(n33[9]));
    nand g5936(n5405 ,n5059 ,n5250);
    not g5937(n3568 ,n3567);
    nand g5938(n5840 ,n5748 ,n5808);
    xor g5939(n4894 ,n4527 ,n4425);
    xnor g5940(n2326 ,n2151 ,n2266);
    or g5941(n2933 ,n2855 ,n2900);
    xnor g5942(n3183 ,n3132 ,n38[7]);
    or g5943(n3046 ,n2996 ,n3022);
    or g5944(n4289 ,n4218 ,n4271);
    nand g5945(n1624 ,n1588 ,n1612);
    nand g5946(n1278 ,n635 ,n730);
    dff g5947(.RN(n1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n32[4]));
    nand g5948(n3008 ,n2964 ,n2978);
    xnor g5949(n6596 ,n3218 ,n3231);
    nand g5950(n1139 ,n33[10] ,n711);
    xnor g5951(n3897 ,n3754 ,n3620);
    nand g5952(n6394 ,n6269 ,n6320);
    nand g5953(n3252 ,n3194 ,n3251);
    xnor g5954(n1777 ,n1636 ,n1722);
    nand g5955(n4444 ,n21[1] ,n4365);
    xnor g5956(n5285 ,n4913 ,n4447);
    not g5957(n3680 ,n3681);
    xnor g5958(n425 ,n373 ,n362);
    buf g5959(n13[3], n10[3]);
    nand g5960(n2177 ,n21[7] ,n2124);
    nand g5961(n2151 ,n6533 ,n2123);
    nand g5962(n1792 ,n1646 ,n1752);
    buf g5963(n13[0], n10[0]);
    nor g5964(n2498 ,n2452 ,n2478);
    nand g5965(n1611 ,n19[6] ,n1594);
    nand g5966(n4039 ,n3873 ,n3979);
    xnor g5967(n2427 ,n2369 ,n2301);
    nand g5968(n527 ,n516 ,n510);
    xnor g5969(n5419 ,n5218 ,n5111);
    nand g5970(n1674 ,n1579 ,n1652);
    xnor g5971(n3345 ,n6574 ,n3322);
    xnor g5972(n6179 ,n6139 ,n6130);
    not g5973(n2949 ,n2948);
    nand g5974(n1491 ,n695 ,n1487);
    xnor g5975(n90 ,n73 ,n51);
    nand g5976(n700 ,n575 ,n585);
    nand g5977(n1052 ,n11[8] ,n711);
    not g5978(n125 ,n124);
    xnor g5979(n5280 ,n4917 ,n4589);
    not g5980(n151 ,n37[2]);
    nand g5981(n3539 ,n3472 ,n3486);
    nand g5982(n1255 ,n839 ,n998);
    nand g5983(n6210 ,n6189 ,n6209);
    not g5984(n4378 ,n4377);
    nor g5985(n2755 ,n2656 ,n2724);
    nand g5986(n1735 ,n1588 ,n1700);
    xnor g5987(n4153 ,n4050 ,n4056);
    nand g5988(n5740 ,n5609 ,n5689);
    xnor g5989(n4880 ,n4496 ,n4465);
    nand g5990(n4079 ,n3977 ,n4030);
    nand g5991(n6286 ,n6507 ,n6249);
    xnor g5992(n6034 ,n5959 ,n5954);
    nand g5993(n3705 ,n3516 ,n3548);
    nor g5994(n2667 ,n2568 ,n2589);
    nand g5995(n507 ,n472 ,n489);
    xor g5996(n6519 ,n6581 ,n6558);
    xnor g5997(n1967 ,n1922 ,n1919);
    xnor g5998(n2491 ,n2439 ,n2422);
    nor g5999(n2652 ,n2565 ,n2594);
    or g6000(n6111 ,n6053 ,n6092);
    nand g6001(n916 ,n1516 ,n712);
    nor g6002(n603 ,n22[6] ,n22[7]);
    xnor g6003(n5697 ,n5546 ,n5453);
    not g6004(n3444 ,n36[0]);
    not g6005(n4361 ,n4360);
    xnor g6006(n3905 ,n3751 ,n3563);
    not g6007(n5073 ,n5072);
    xor g6008(n4927 ,n4671 ,n4481);
    nand g6009(n1517 ,n108 ,n112);
    nor g6010(n2996 ,n2887 ,n2965);
    or g6011(n482 ,n447 ,n463);
    nor g6012(n2887 ,n2795 ,n2851);
    nand g6013(n5902 ,n5807 ,n5825);
    xnor g6014(n38[5] ,n2466 ,n2506);
    nand g6015(n438 ,n224 ,n419);
    xor g6016(n2328 ,n2233 ,n2272);
    nand g6017(n2590 ,n40[10] ,n6521);
    or g6018(n6162 ,n6154 ,n6113);
    nand g6019(n6106 ,n6045 ,n6071);
    xor g6020(n4882 ,n4698 ,n4580);
    or g6021(n5894 ,n5824 ,n5829);
    nor g6022(n2695 ,n2566 ,n2627);
    nand g6023(n6185 ,n6168 ,n6153);
    xor g6024(n2114 ,n2100 ,n2086);
    nand g6025(n1025 ,n1540 ,n713);
    not g6026(n5637 ,n5636);
    xor g6027(n3913 ,n3750 ,n3514);
    nand g6028(n99 ,n83 ,n98);
    not g6029(n162 ,n36[4]);
    or g6030(n3694 ,n3517 ,n3594);
    nand g6031(n1346 ,n915 ,n1095);
    nand g6032(n5943 ,n5809 ,n5897);
    nand g6033(n1300 ,n1056 ,n805);
    nand g6034(n1285 ,n1038 ,n862);
    nand g6035(n4842 ,n4497 ,n4578);
    or g6036(n4768 ,n4491 ,n4482);
    not g6037(n5175 ,n5174);
    nor g6038(n2690 ,n2568 ,n2625);
    xnor g6039(n1905 ,n1833 ,n1798);
    xnor g6040(n1819 ,n1768 ,n1645);
    nand g6041(n797 ,n26[6] ,n723);
    nand g6042(n5497 ,n5269 ,n5365);
    xnor g6043(n2918 ,n2870 ,n2739);
    xnor g6044(n3328 ,n41[15] ,n6588);
    nand g6045(n2586 ,n40[9] ,n6520);
    dff g6046(.RN(n1), .SN(1'b1), .CK(n0), .D(n1400), .Q(n27[10]));
    nand g6047(n798 ,n26[5] ,n723);
    nand g6048(n6059 ,n5882 ,n6037);
    nand g6049(n1858 ,n1803 ,n1804);
    or g6050(n4718 ,n4477 ,n4640);
    nand g6051(n217 ,n159 ,n155);
    buf g6052(n36[5] ,n1513);
    nand g6053(n2405 ,n2354 ,n2388);
    xnor g6054(n5233 ,n4957 ,n4789);
    dff g6055(.RN(n1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n31[7]));
    nand g6056(n6104 ,n6020 ,n6078);
    nand g6057(n1262 ,n847 ,n1008);
    nor g6058(n2400 ,n2332 ,n2380);
    nand g6059(n6343 ,n6547 ,n6248);
    xnor g6060(n2633 ,n6525 ,n40[14]);
    nand g6061(n4137 ,n4019 ,n4076);
    nand g6062(n2906 ,n2789 ,n2873);
    or g6063(n3660 ,n3530 ,n3537);
    nand g6064(n851 ,n16[3] ,n714);
    xnor g6065(n3401 ,n6549 ,n6564);
    dff g6066(.RN(n1), .SN(1'b1), .CK(n0), .D(n1197), .Q(n32[0]));
    xnor g6067(n6538 ,n3312 ,n3300);
    nand g6068(n5571 ,n5378 ,n5481);
    nand g6069(n5474 ,n5222 ,n5381);
    nand g6070(n5980 ,n5954 ,n5927);
    nand g6071(n5402 ,n4756 ,n5276);
    nand g6072(n131 ,n24[6] ,n130);
    xnor g6073(n684 ,n35[0] ,n31[0]);
    or g6074(n249 ,n182 ,n194);
    nand g6075(n3244 ,n3188 ,n3243);
    nor g6076(n2744 ,n2674 ,n2738);
    nand g6077(n5006 ,n4650 ,n4804);
    not g6078(n290 ,n289);
    not g6079(n5851 ,n5850);
    nand g6080(n5008 ,n4557 ,n4828);
    nor g6081(n6233 ,n41[15] ,n6589);
    nand g6082(n888 ,n33[7] ,n554);
    nand g6083(n2208 ,n2095 ,n2163);
    nand g6084(n980 ,n27[2] ,n715);
    nand g6085(n3551 ,n3476 ,n19[6]);
    nand g6086(n2227 ,n2140 ,n2191);
    nor g6087(n2745 ,n2635 ,n2690);
    nand g6088(n967 ,n27[8] ,n715);
    xnor g6089(n5596 ,n5454 ,n5209);
    or g6090(n5328 ,n5285 ,n5190);
    xnor g6091(n5955 ,n5881 ,n5850);
    nand g6092(n4986 ,n4673 ,n4801);
    nand g6093(n6373 ,n38[11] ,n6246);
    nor g6094(n2012 ,n1985 ,n1997);
    xor g6095(n5967 ,n5864 ,n5835);
    nand g6096(n1718 ,n1579 ,n1676);
    nor g6097(n3435 ,n3390 ,n3434);
    nand g6098(n4610 ,n4378 ,n20[0]);
    nand g6099(n908 ,n1545 ,n712);
    nand g6100(n720 ,n18[0] ,n662);
    nand g6101(n405 ,n339 ,n385);
    nor g6102(n5855 ,n5714 ,n5788);
    xnor g6103(n2923 ,n2868 ,n2738);
    nand g6104(n6173 ,n6143 ,n6120);
    nand g6105(n2146 ,n6536 ,n2122);
    xnor g6106(n4017 ,n3525 ,n3910);
    nand g6107(n706 ,n576 ,n568);
    nand g6108(n6313 ,n6548 ,n6248);
    not g6109(n1585 ,n36[0]);
    xnor g6110(n5194 ,n4902 ,n4453);
    nand g6111(n4818 ,n4568 ,n4453);
    not g6112(n1636 ,n1637);
    nand g6113(n1921 ,n1903 ,n1905);
    nand g6114(n2477 ,n2463 ,n2428);
    nand g6115(n3379 ,n3332 ,n3378);
    nand g6116(n4582 ,n21[2] ,n4378);
    or g6117(n487 ,n403 ,n474);
    nand g6118(n5905 ,n5812 ,n5822);
    xnor g6119(n3937 ,n3746 ,n3513);
    nand g6120(n5711 ,n5532 ,n5626);
    nor g6121(n2797 ,n2602 ,n2714);
    nand g6122(n1343 ,n942 ,n1092);
    nand g6123(n3855 ,n3665 ,n3824);
    nand g6124(n4276 ,n4238 ,n4256);
    xnor g6125(n6500 ,n3051 ,n3048);
    or g6126(n4238 ,n4154 ,n4207);
    nand g6127(n4243 ,n4192 ,n4206);
    nand g6128(n5909 ,n5738 ,n5849);
    nand g6129(n2619 ,n2585 ,n2574);
    or g6130(n4747 ,n4426 ,n4429);
    nand g6131(n5013 ,n4511 ,n4834);
    nand g6132(n1160 ,n1554 ,n716);
    xnor g6133(n91 ,n65 ,n55);
    nand g6134(n799 ,n26[4] ,n723);
    nand g6135(n5919 ,n5858 ,n5903);
    nor g6136(n6229 ,n41[7] ,n6593);
    nand g6137(n6069 ,n5992 ,n6030);
    xnor g6138(n2467 ,n2421 ,n2360);
    dff g6139(.RN(n1), .SN(1'b1), .CK(n0), .D(n1238), .Q(n33[6]));
    nand g6140(n4977 ,n4584 ,n4782);
    xnor g6141(n3050 ,n3019 ,n3023);
    nand g6142(n849 ,n1506 ,n714);
    nand g6143(n1317 ,n905 ,n1059);
    nor g6144(n2609 ,n2567 ,n2593);
    or g6145(n4876 ,n4563 ,n4440);
    nor g6146(n2802 ,n2613 ,n2716);
    nor g6147(n614 ,n33[12] ,n35[12]);
    nand g6148(n3807 ,n3699 ,n3692);
    nand g6149(n4804 ,n4619 ,n4421);
    xnor g6150(n1608 ,n1562 ,n19[6]);
    nand g6151(n4688 ,n4389 ,n20[2]);
    dff g6152(.RN(n1), .SN(1'b1), .CK(n0), .D(n1303), .Q(n11[3]));
    nand g6153(n6238 ,n41[12] ,n6592);
    nor g6154(n5346 ,n5131 ,n5164);
    not g6155(n3299 ,n3298);
    nand g6156(n3199 ,n3158 ,n3179);
    nand g6157(n5359 ,n5072 ,n5195);
    nor g6158(n3426 ,n3403 ,n3425);
    nand g6159(n1420 ,n798 ,n1176);
    xnor g6160(n704 ,n23[3] ,n16[3]);
    xnor g6161(n2911 ,n2878 ,n2858);
    xnor g6162(n3408 ,n6552 ,n39[3]);
    nand g6163(n5117 ,n4733 ,n5016);
    xnor g6164(n3355 ,n6577 ,n3353);
    not g6165(n3257 ,n3256);
    nand g6166(n399 ,n351 ,n364);
    nand g6167(n234 ,n172 ,n153);
    nand g6168(n4697 ,n21[6] ,n4369);
    or g6169(n4745 ,n4430 ,n4617);
    nor g6170(n3566 ,n3490 ,n3500);
    nand g6171(n4235 ,n4135 ,n4208);
    xnor g6172(n4341 ,n4324 ,n4319);
    nand g6173(n3699 ,n3583 ,n3596);
    nor g6174(n2519 ,n2505 ,n2493);
    nand g6175(n5889 ,n5622 ,n5833);
    xor g6176(n4896 ,n4670 ,n4464);
    or g6177(n3977 ,n3862 ,n3889);
    not g6178(n2754 ,n2753);
    nor g6179(n5466 ,n5297 ,n5408);
    nand g6180(n1374 ,n630 ,n761);
    dff g6181(.RN(n1), .SN(1'b1), .CK(n0), .D(n1316), .Q(n10[6]));
    xor g6182(n6574 ,n1781 ,n1678);
    not g6183(n4561 ,n4560);
    nor g6184(n2815 ,n2659 ,n2747);
    nand g6185(n2071 ,n20[4] ,n20[3]);
    or g6186(n5661 ,n5500 ,n5539);
    dff g6187(.RN(n1), .SN(1'b1), .CK(n0), .D(n1218), .Q(n30[0]));
    xnor g6188(n6125 ,n6053 ,n6092);
    or g6189(n5848 ,n5805 ,n5784);
    nand g6190(n3640 ,n3474 ,n3485);
    xor g6191(n1557 ,n1792 ,n1782);
    nand g6192(n1208 ,n34[6] ,n838);
    xnor g6193(n6585 ,n2031 ,n2050);
    xnor g6194(n5205 ,n4924 ,n4528);
    xor g6195(n4948 ,n4554 ,n4569);
    or g6196(n271 ,n223 ,n211);
    nand g6197(n1103 ,n1521 ,n716);
    nand g6198(n4498 ,n21[7] ,n4389);
    nand g6199(n996 ,n25[1] ,n714);
    nand g6200(n969 ,n21[1] ,n714);
    nand g6201(n1758 ,n1697 ,n1720);
    nor g6202(n3439 ,n3394 ,n3438);
    or g6203(n4709 ,n4625 ,n4441);
    xnor g6204(n1951 ,n1880 ,n1916);
    nor g6205(n2727 ,n2567 ,n2622);
    xnor g6206(n694 ,n567 ,n26[3]);
    nand g6207(n962 ,n24[3] ,n715);
    nor g6208(n2658 ,n2568 ,n2591);
    nand g6209(n3594 ,n3482 ,n19[0]);
    xnor g6210(n5423 ,n5190 ,n5285);
    xnor g6211(n5860 ,n5782 ,n5806);
    xnor g6212(n1900 ,n1848 ,n1790);
    nor g6213(n2014 ,n2004 ,n1994);
    nand g6214(n3922 ,n3829 ,n3868);
    nand g6215(n2776 ,n2674 ,n2738);
    nand g6216(n6364 ,n6544 ,n6248);
    nand g6217(n1367 ,n818 ,n1118);
    nor g6218(n5330 ,n5062 ,n5224);
    nand g6219(n3996 ,n3858 ,n3908);
    not g6220(n2997 ,n2989);
    xnor g6221(n5760 ,n5614 ,n5542);
    or g6222(n5712 ,n5512 ,n5639);
    nand g6223(n212 ,n159 ,n152);
    nor g6224(n3374 ,n3371 ,n3373);
    xnor g6225(n3896 ,n3742 ,n3607);
    nand g6226(n5679 ,n5503 ,n5513);
    nand g6227(n1476 ,n917 ,n1245);
    or g6228(n3960 ,n3938 ,n3937);
    nor g6229(n2749 ,n2655 ,n2696);
    nand g6230(n5746 ,n5506 ,n5671);
    dff g6231(.RN(n1), .SN(1'b1), .CK(n0), .D(n1469), .Q(n22[0]));
    nor g6232(n2685 ,n2568 ,n2628);
    nand g6233(n1739 ,n1582 ,n1700);
    nand g6234(n1315 ,n1167 ,n955);
    nand g6235(n6379 ,n6501 ,n6249);
    nand g6236(n899 ,n24[4] ,n715);
    nor g6237(n4525 ,n4414 ,n4408);
    nand g6238(n1334 ,n897 ,n1087);
    or g6239(n261 ,n220 ,n221);
    nand g6240(n3055 ,n3031 ,n3035);
    nand g6241(n943 ,n28[1] ,n717);
    not g6242(n4692 ,n4691);
    not g6243(n5872 ,n4359);
    nand g6244(n4456 ,n4376 ,n20[5]);
    nand g6245(n390 ,n321 ,n347);
    or g6246(n4728 ,n4462 ,n4620);
    nand g6247(n3088 ,n3034 ,n3087);
    nand g6248(n1006 ,n12[12] ,n711);
    nand g6249(n1706 ,n1586 ,n1676);
    nor g6250(n2803 ,n2604 ,n2715);
    or g6251(n2708 ,n2567 ,n2620);
    dff g6252(.RN(n1), .SN(1'b1), .CK(n0), .D(n1320), .Q(n10[4]));
    nand g6253(n395 ,n346 ,n378);
    nand g6254(n1265 ,n848 ,n1011);
    nand g6255(n822 ,n34[2] ,n717);
    nand g6256(n896 ,n24[7] ,n715);
    nand g6257(n1463 ,n1132 ,n1382);
    not g6258(n557 ,n714);
    nand g6259(n3801 ,n3634 ,n3701);
    xnor g6260(n4942 ,n4564 ,n4485);
    xnor g6261(n5436 ,n5219 ,n5109);
    nand g6262(n1398 ,n961 ,n1154);
    xor g6263(n1643 ,n1626 ,n1615);
    buf g6264(n36[7] ,n1515);
    nand g6265(n2232 ,n2147 ,n2211);
    not g6266(n231 ,n230);
    nand g6267(n6004 ,n5936 ,n5982);
    nand g6268(n3309 ,n3304 ,n3308);
    nor g6269(n2712 ,n2565 ,n2625);
    nand g6270(n2823 ,n2740 ,n2803);
    nand g6271(n4807 ,n4443 ,n4447);
    nand g6272(n5675 ,n5577 ,n5538);
    nand g6273(n1167 ,n33[13] ,n711);
    nand g6274(n4579 ,n4388 ,n20[6]);
    not g6275(n387 ,n386);
    xnor g6276(n6208 ,n6195 ,n6184);
    xnor g6277(n2929 ,n2871 ,n2771);
    nor g6278(n322 ,n231 ,n291);
    nand g6279(n4984 ,n4515 ,n4807);
    not g6280(n238 ,n237);
    nand g6281(n1687 ,n1576 ,n1651);
    not g6282(n2264 ,n2263);
    nand g6283(n6267 ,n41[12] ,n6254);
    not g6284(n54 ,n37[3]);
    nand g6285(n237 ,n169 ,n144);
    or g6286(n6163 ,n6121 ,n6145);
    nand g6287(n900 ,n23[11] ,n715);
    xnor g6288(n38[3] ,n2414 ,n2409);
    nor g6289(n6464 ,n6428 ,n6425);
    dff g6290(.RN(n1), .SN(1'b1), .CK(n0), .D(n1455), .Q(n31[4]));
    nand g6291(n975 ,n34[0] ,n717);
    nand g6292(n1048 ,n2[2] ,n713);
    nand g6293(n824 ,n23[2] ,n715);
    nand g6294(n5370 ,n5129 ,n5197);
    xor g6295(n5427 ,n5183 ,n5222);
    nand g6296(n1714 ,n1580 ,n1675);
    xor g6297(n41[15] ,n6140 ,n6221);
    xnor g6298(n38[15] ,n2508 ,n2564);
    xnor g6299(n6568 ,n5957 ,n5910);
    nand g6300(n5120 ,n4723 ,n5045);
    nand g6301(n4247 ,n4181 ,n4217);
    nand g6302(n1467 ,n939 ,n1386);
    nand g6303(n2411 ,n2350 ,n2387);
    xnor g6304(n1944 ,n1883 ,n1914);
    or g6305(n3093 ,n38[8] ,n6581);
    nand g6306(n213 ,n167 ,n146);
    not g6307(n3630 ,n3629);
    nor g6308(n5277 ,n4978 ,n5057);
    nand g6309(n987 ,n16[8] ,n714);
    nand g6310(n4260 ,n4236 ,n4246);
    nand g6311(n5027 ,n4661 ,n4821);
    nand g6312(n3638 ,n3474 ,n3476);
    nor g6313(n608 ,n33[9] ,n35[9]);
    nand g6314(n968 ,n29[6] ,n721);
    nand g6315(n1076 ,n10[4] ,n710);
    nand g6316(n4350 ,n4338 ,n4349);
    xnor g6317(n3910 ,n3770 ,n3623);
    nand g6318(n1296 ,n875 ,n1053);
    not g6319(n1587 ,n36[2]);
    dff g6320(.RN(n1), .SN(1'b1), .CK(n0), .D(n1456), .Q(n31[3]));
    nor g6321(n2563 ,n2518 ,n2562);
    xnor g6322(n1818 ,n1767 ,n1645);
    xnor g6323(n6196 ,n6173 ,n6179);
    xnor g6324(n688 ,n23[1] ,n16[1]);
    not g6325(n43 ,n42);
    nand g6326(n4220 ,n4168 ,n4188);
    nand g6327(n1080 ,n27[10] ,n718);
    nand g6328(n1185 ,n29[1] ,n724);
    nor g6329(n2675 ,n2568 ,n2584);
    xnor g6330(n3023 ,n2975 ,n2954);
    nand g6331(n5374 ,n5091 ,n5243);
    nor g6332(n1836 ,n1779 ,n1824);
    nand g6333(n6446 ,n6289 ,n6361);
    xor g6334(n40[9] ,n6602 ,n38[10]);
    nor g6335(n1949 ,n1884 ,n1927);
    nand g6336(n4129 ,n3970 ,n4065);
    xor g6337(n5862 ,n5622 ,n5816);
    nand g6338(n223 ,n172 ,n150);
    nand g6339(n1489 ,n719 ,n1483);
    xnor g6340(n4325 ,n4300 ,n4278);
    xnor g6341(n4263 ,n3975 ,n4234);
    nand g6342(n1126 ,n17[7] ,n724);
    nor g6343(n4527 ,n4394 ,n4418);
    nand g6344(n1333 ,n659 ,n738);
    nor g6345(n3031 ,n2998 ,n3011);
    not g6346(n2474 ,n2473);
    xnor g6347(n1826 ,n1645 ,n1758);
    nor g6348(n3626 ,n3496 ,n3495);
    nand g6349(n1361 ,n1115 ,n881);
    nand g6350(n5278 ,n4709 ,n5106);
    xnor g6351(n6545 ,n3331 ,n3378);
    nand g6352(n2215 ,n6538 ,n2178);
    nand g6353(n1732 ,n1586 ,n1700);
    xor g6354(n6566 ,n5595 ,n5278);
    xnor g6355(n2490 ,n2441 ,n2463);
    nand g6356(n1741 ,n1691 ,n1731);
    nand g6357(n1227 ,n982 ,n726);
    nand g6358(n1382 ,n651 ,n767);
    nand g6359(n640 ,n21[0] ,n30[0]);
    nor g6360(n5551 ,n5321 ,n5464);
    xnor g6361(n2858 ,n2773 ,n2742);
    or g6362(n6143 ,n6131 ,n6110);
    or g6363(n4237 ,n4135 ,n4208);
    nand g6364(n5547 ,n5319 ,n5463);
    xnor g6365(n5225 ,n4949 ,n4541);
    xnor g6366(n3973 ,n3755 ,n3878);
    not g6367(n3330 ,n3329);
    nand g6368(n4541 ,n20[2] ,n4374);
    nand g6369(n4994 ,n4653 ,n4825);
    nand g6370(n3713 ,n3508 ,n3507);
    xnor g6371(n6536 ,n3303 ,n3308);
    or g6372(n509 ,n466 ,n506);
    nand g6373(n6124 ,n6060 ,n6098);
    nand g6374(n6397 ,n6274 ,n6324);
    not g6375(n3468 ,n3467);
    not g6376(n4360 ,n37[7]);
    nand g6377(n1289 ,n868 ,n1043);
    not g6378(n2734 ,n2733);
    nor g6379(n116 ,n32[1] ,n114);
    or g6380(n5562 ,n5209 ,n5454);
    nor g6381(n3316 ,n3288 ,n3315);
    nor g6382(n6234 ,n41[5] ,n6595);
    nand g6383(n3110 ,n6577 ,n6554);
    nand g6384(n659 ,n19[3] ,n27[3]);
    nand g6385(n4828 ,n4639 ,n4495);
    or g6386(n2985 ,n2925 ,n2955);
    nand g6387(n3368 ,n3364 ,n3367);
    nand g6388(n1070 ,n10[10] ,n711);
    nand g6389(n5491 ,n5263 ,n5360);
    nor g6390(n4515 ,n4398 ,n4392);
    xnor g6391(n5420 ,n5283 ,n5210);
    buf g6392(n15[3], 1'b0);
    not g6393(n177 ,n161);
    nor g6394(n6495 ,n2567 ,n2631);
    nand g6395(n3204 ,n3165 ,n3180);
    nor g6396(n6247 ,n25[1] ,n6237);
    nand g6397(n1164 ,n6[0] ,n557);
    nand g6398(n872 ,n33[9] ,n712);
    dff g6399(.RN(n1), .SN(1'b1), .CK(n0), .D(n1231), .Q(n12[13]));
    nor g6400(n2663 ,n2568 ,n2592);
    xnor g6401(n3220 ,n3162 ,n3175);
    nand g6402(n4599 ,n20[2] ,n4365);
    nor g6403(n2149 ,n2114 ,n2121);
    nor g6404(n1972 ,n1925 ,n1952);
    nand g6405(n1405 ,n859 ,n1159);
    xnor g6406(n377 ,n309 ,n269);
    xnor g6407(n3223 ,n3163 ,n3176);
    xnor g6408(n374 ,n318 ,n196);
    nand g6409(n1084 ,n10[1] ,n555);
    nor g6410(n6148 ,n6129 ,n6093);
    nand g6411(n206 ,n165 ,n153);
    nand g6412(n409 ,n387 ,n371);
    nor g6413(n2353 ,n2289 ,n2287);
    or g6414(n385 ,n344 ,n337);
    nand g6415(n6307 ,n41[5] ,n6254);
    nand g6416(n4455 ,n21[2] ,n4371);
    xnor g6417(n1755 ,n1680 ,n1645);
    nand g6418(n6408 ,n6306 ,n6342);
    nor g6419(n1940 ,n1915 ,n1901);
    nand g6420(n826 ,n17[4] ,n721);
    nand g6421(n973 ,n27[5] ,n715);
    nand g6422(n3362 ,n41[5] ,n3361);
    xnor g6423(n5231 ,n4955 ,n4791);
    xnor g6424(n2118 ,n2104 ,n2086);
    xor g6425(n5759 ,n5591 ,n5629);
    not g6426(n1588 ,n1587);
    nand g6427(n6020 ,n5926 ,n5977);
    nand g6428(n5276 ,n4855 ,n5142);
    nand g6429(n3854 ,n3678 ,n3805);
    xnor g6430(n1635 ,n1592 ,n1616);
    nand g6431(n4468 ,n21[6] ,n4389);
    nand g6432(n3728 ,n3514 ,n3510);
    nand g6433(n821 ,n23[1] ,n715);
    not g6434(n3442 ,n36[1]);
    nand g6435(n4190 ,n4116 ,n4149);
    nor g6436(n2515 ,n2501 ,n2492);
    nand g6437(n4536 ,n21[4] ,n4388);
    nand g6438(n954 ,n35[12] ,n712);
    dff g6439(.RN(n1), .SN(1'b1), .CK(n0), .D(n1244), .Q(n31[2]));
    nor g6440(n2041 ,n2016 ,n2040);
    not g6441(n3476 ,n3475);
    nand g6442(n2181 ,n6538 ,n2150);
    nand g6443(n1702 ,n1577 ,n1676);
    nor g6444(n2834 ,n2702 ,n2752);
    nand g6445(n6323 ,n38[7] ,n6246);
    nand g6446(n3306 ,n3286 ,n3305);
    nand g6447(n272 ,n189 ,n191);
    xnor g6448(n6056 ,n5949 ,n6018);
    nand g6449(n1269 ,n633 ,n725);
    not g6450(n2076 ,n2075);
    nand g6451(n641 ,n21[1] ,n30[1]);
    nand g6452(n3507 ,n3462 ,n3482);
    xor g6453(n4922 ,n4519 ,n4627);
    or g6454(n5237 ,n5117 ,n5076);
    xor g6455(n1652 ,n1634 ,n1638);
    not g6456(n2266 ,n2265);
    nor g6457(n2611 ,n2567 ,n2588);
    nand g6458(n2830 ,n2737 ,n2788);
    nand g6459(n3697 ,n3608 ,n3504);
    nand g6460(n281 ,n232 ,n187);
    nand g6461(n2631 ,n2584 ,n2576);
    not g6462(n161 ,n160);
    not g6463(n2061 ,n6537);
    nand g6464(n1401 ,n965 ,n1158);
    nand g6465(n5036 ,n4535 ,n4810);
    nand g6466(n3813 ,n3613 ,n3726);
    nand g6467(n1029 ,n1542 ,n557);
    nand g6468(n3208 ,n3163 ,n3176);
    nand g6469(n5979 ,n5879 ,n5930);
    not g6470(n562 ,n17[1]);
    nor g6471(n2837 ,n2703 ,n2751);
    nand g6472(n1465 ,n935 ,n1384);
    xnor g6473(n422 ,n364 ,n350);
    nand g6474(n906 ,n1543 ,n712);
    xnor g6475(n1996 ,n1947 ,n1933);
    nand g6476(n4259 ,n4195 ,n4228);
    not g6477(n1851 ,n1844);
    xnor g6478(n1615 ,n19[3] ,n1572);
    or g6479(n4334 ,n4315 ,n4326);
    nand g6480(n3865 ,n3656 ,n3815);
    not g6481(n4389 ,n4391);
    xnor g6482(n6572 ,n6208 ,n6213);
    nand g6483(n5034 ,n4505 ,n4799);
    nand g6484(n1860 ,n1749 ,n1805);
    nand g6485(n4476 ,n4386 ,n20[2]);
    nand g6486(n3159 ,n3112 ,n3139);
    nand g6487(n1021 ,n3[4] ,n713);
    nand g6488(n1423 ,n989 ,n1178);
    nand g6489(n4861 ,n4614 ,n4444);
    nand g6490(n643 ,n31[4] ,n35[4]);
    nor g6491(n4699 ,n4394 ,n4406);
    nor g6492(n5585 ,n5369 ,n5447);
    nand g6493(n1409 ,n974 ,n1165);
    xnor g6494(n2950 ,n2857 ,n2897);
    xnor g6495(n6543 ,n3337 ,n3374);
    nor g6496(n6103 ,n6080 ,n6028);
    nand g6497(n5381 ,n5185 ,n5183);
    nand g6498(n853 ,n1503 ,n714);
    nand g6499(n4166 ,n4136 ,n4103);
    nand g6500(n2192 ,n6537 ,n2148);
    nand g6501(n6167 ,n6122 ,n6146);
    xnor g6502(n5701 ,n5585 ,n5577);
    nand g6503(n6290 ,n40[3] ,n6250);
    xnor g6504(n2312 ,n2253 ,n2119);
    nand g6505(n4044 ,n3925 ,n3981);
    nand g6506(n5140 ,n4738 ,n5043);
    nand g6507(n5925 ,n5802 ,n5875);
    nand g6508(n383 ,n279 ,n352);
    nand g6509(n1729 ,n1624 ,n1685);
    xnor g6510(n1525 ,n529 ,n540);
    nand g6511(n4474 ,n20[5] ,n4365);
    nor g6512(n6467 ,n6436 ,n6446);
    or g6513(n4134 ,n3939 ,n4063);
    nand g6514(n4820 ,n4627 ,n4634);
    dff g6515(.RN(n1), .SN(1'b1), .CK(n0), .D(n1499), .Q(n18[0]));
    nand g6516(n4872 ,n4426 ,n4429);
    not g6517(n2788 ,n2787);
    xnor g6518(n4065 ,n3947 ,n3877);
    nand g6519(n2620 ,n2592 ,n2577);
    nor g6520(n1534 ,n75 ,n105);
    nand g6521(n5803 ,n5650 ,n5705);
    nand g6522(n1701 ,n1586 ,n1649);
    xor g6523(n40[8] ,n6603 ,n38[9]);
    nand g6524(n1245 ,n28[7] ,n1191);
    nand g6525(n6404 ,n6303 ,n6332);
    xnor g6526(n5510 ,n5191 ,n5406);
    nor g6527(n2612 ,n2567 ,n2591);
    not g6528(n2527 ,n2526);
    nand g6529(n1340 ,n944 ,n1163);
    xnor g6530(n2079 ,n21[4] ,n20[4]);
    xnor g6531(n2237 ,n2154 ,n2109);
    nand g6532(n3043 ,n3007 ,n3025);
    nor g6533(n2148 ,n2116 ,n2126);
    nand g6534(n5393 ,n5279 ,n5180);
    nand g6535(n4860 ,n4628 ,n4635);
    nand g6536(n5908 ,n5733 ,n5840);
    dff g6537(.RN(n1), .SN(1'b1), .CK(n0), .D(n1390), .Q(n33[11]));
    nand g6538(n5812 ,n5684 ,n5742);
    or g6539(n5329 ,n5213 ,n5212);
    nand g6540(n35[14] ,n6458 ,n6480);
    nand g6541(n5007 ,n4538 ,n4824);
    or g6542(n2035 ,n2019 ,n2025);
    nand g6543(n844 ,n16[5] ,n714);
    nand g6544(n2175 ,n6541 ,n2126);
    nor g6545(n3373 ,n6569 ,n3372);
    not g6546(n170 ,n173);
    nand g6547(n5787 ,n5716 ,n5647);
    nand g6548(n828 ,n17[2] ,n721);
    xnor g6549(n2485 ,n2450 ,n2417);
    not g6550(n4398 ,n21[2]);
    xnor g6551(n5216 ,n4922 ,n4634);
    dff g6552(.RN(n1), .SN(1'b1), .CK(n0), .D(n1370), .Q(n23[4]));
    nand g6553(n1372 ,n656 ,n760);
    nand g6554(n2187 ,n6539 ,n2149);
    xnor g6555(n3787 ,n3565 ,n3641);
    nand g6556(n1444 ,n1015 ,n1267);
    nand g6557(n5056 ,n4704 ,n5023);
    nand g6558(n220 ,n161 ,n155);
    dff g6559(.RN(n1), .SN(1'b1), .CK(n0), .D(n1323), .Q(n34[11]));
    nor g6560(n1816 ,n1754 ,n1793);
    nand g6561(n3541 ,n3480 ,n19[4]);
    nand g6562(n4605 ,n21[4] ,n4384);
    xnor g6563(n2424 ,n2367 ,n2059);
    or g6564(n4720 ,n4639 ,n4495);
    nand g6565(n1473 ,n976 ,n1410);
    nor g6566(n4507 ,n4412 ,n4399);
    not g6567(n5569 ,n5568);
    nor g6568(n6235 ,n41[14] ,n6590);
    xnor g6569(n5972 ,n5865 ,n5855);
    nand g6570(n1323 ,n936 ,n1144);
    xnor g6571(n4013 ,n3936 ,n3901);
    nand g6572(n948 ,n21[6] ,n714);
    nand g6573(n356 ,n259 ,n325);
    nor g6574(n879 ,n570 ,n711);
    xnor g6575(n2508 ,n2475 ,n2440);
    or g6576(n5888 ,n5729 ,n5837);
    nor g6577(n2810 ,n2705 ,n2756);
    nand g6578(n1236 ,n1037 ,n732);
    nand g6579(n1673 ,n1584 ,n1652);
    or g6580(n5235 ,n5070 ,n5080);
    xnor g6581(n5192 ,n4900 ,n4428);
    xnor g6582(n3340 ,n41[13] ,n6586);
    xor g6583(n4945 ,n4690 ,n4603);
    nand g6584(n3990 ,n3901 ,n3936);
    xnor g6585(n1810 ,n1648 ,n1753);
    nand g6586(n3641 ,n3472 ,n3482);
    nand g6587(n3236 ,n3193 ,n3235);
    nor g6588(n1677 ,n1643 ,n1654);
    nand g6589(n284 ,n179 ,n228);
    xor g6590(n4920 ,n4544 ,n4473);
    xnor g6591(n3001 ,n2959 ,n2896);
    or g6592(n4712 ,n4588 ,n4626);
    nor g6593(n5454 ,n5061 ,n5330);
    nand g6594(n2176 ,n6540 ,n2121);
    nand g6595(n3849 ,n3651 ,n3822);
    nand g6596(n3021 ,n3009 ,n3012);
    xor g6597(n3774 ,n3627 ,n3575);
    nand g6598(n1709 ,n1584 ,n1677);
    nand g6599(n4481 ,n21[5] ,n4382);
    xnor g6600(n3890 ,n3741 ,n3556);
    or g6601(n3661 ,n3588 ,n3506);
    nor g6602(n3682 ,n3559 ,n3560);
    nand g6603(n4195 ,n4121 ,n4157);
    nand g6604(n1310 ,n1068 ,n954);
    xnor g6605(n5153 ,n4966 ,n4441);
    nand g6606(n1394 ,n948 ,n1150);
    dff g6607(.RN(n1), .SN(1'b1), .CK(n0), .D(n18[2]), .Q(n15[6]));
    nor g6608(n2636 ,n2566 ,n2591);
    nand g6609(n977 ,n20[6] ,n556);
    nor g6610(n3434 ,n3415 ,n3433);
    nor g6611(n3431 ,n3391 ,n3430);
    nand g6612(n4834 ,n4478 ,n4493);
    nand g6613(n4632 ,n4388 ,n20[5]);
    nor g6614(n2842 ,n2730 ,n2794);
    nand g6615(n6473 ,n6344 ,n6412);
    nand g6616(n1109 ,n32[5] ,n555);
    xnor g6617(n3895 ,n3748 ,n3628);
    nand g6618(n3516 ,n3470 ,n3480);
    nor g6619(n2407 ,n2347 ,n2384);
    dff g6620(.RN(n1), .SN(1'b1), .CK(n0), .D(n1229), .Q(n12[15]));
    xnor g6621(n5230 ,n4953 ,n4778);
    dff g6622(.RN(n1), .SN(1'b1), .CK(n0), .D(n1462), .Q(n30[2]));
    not g6623(n360 ,n359);
    nand g6624(n1364 ,n816 ,n1116);
    xnor g6625(n4015 ,n3940 ,n3907);
    xnor g6626(n4302 ,n4265 ,n4269);
    xor g6627(n3776 ,n3558 ,n3519);
    nor g6628(n2509 ,n2455 ,n2506);
    nand g6629(n5485 ,n5097 ,n5394);
    xnor g6630(n301 ,n241 ,n188);
    xnor g6631(n5303 ,n5137 ,n5145);
    nand g6632(n912 ,n23[8] ,n715);
    nor g6633(n2516 ,n2481 ,n2495);
    nand g6634(n1121 ,n31[3] ,n720);
    not g6635(n1580 ,n1589);
    nand g6636(n6270 ,n6557 ,n6251);
    not g6637(n3492 ,n3480);
    xnor g6638(n5232 ,n4959 ,n4780);
    xnor g6639(n2290 ,n2223 ,n2118);
    nand g6640(n4212 ,n4074 ,n4198);
    xnor g6641(n5304 ,n5149 ,n5071);
    not g6642(n2421 ,n2420);
    nand g6643(n3628 ,n3484 ,n19[5]);
    nor g6644(n1829 ,n1782 ,n1792);
    or g6645(n3092 ,n38[12] ,n6585);
    nand g6646(n2161 ,n6533 ,n2127);
    nand g6647(n815 ,n34[4] ,n717);
    nand g6648(n5703 ,n5586 ,n5680);
    xnor g6649(n300 ,n183 ,n212);
    not g6650(n2763 ,n2762);
    dff g6651(.RN(n1), .SN(1'b1), .CK(n0), .D(n1206), .Q(n34[4]));
    nand g6652(n192 ,n161 ,n146);
    dff g6653(.RN(n1), .SN(1'b1), .CK(n0), .D(n1460), .Q(n30[4]));
    xnor g6654(n2240 ,n2119 ,n2155);
    xnor g6655(n4879 ,n4467 ,n4575);
    nand g6656(n203 ,n165 ,n152);
    nand g6657(n6076 ,n6052 ,n6033);
    nand g6658(n5099 ,n4741 ,n5053);
    xnor g6659(n6498 ,n2974 ,n2966);
    nand g6660(n1072 ,n10[8] ,n711);
    nand g6661(n6443 ,n6307 ,n6376);
    nand g6662(n2047 ,n2046 ,n2035);
    nand g6663(n4429 ,n20[6] ,n4367);
    nand g6664(n277 ,n178 ,n215);
    nor g6665(n1497 ,n1493 ,n1486);
    nor g6666(n2410 ,n2357 ,n2385);
    nand g6667(n6120 ,n6106 ,n6096);
    nand g6668(n1469 ,n1145 ,n1388);
    nand g6669(n981 ,n20[4] ,n714);
    nand g6670(n3578 ,n3472 ,n3480);
    xor g6671(n5432 ,n5212 ,n5215);
    nand g6672(n5040 ,n4523 ,n4805);
    xor g6673(n6513 ,n6575 ,n6552);
    nand g6674(n1432 ,n996 ,n1188);
    nand g6675(n1264 ,n646 ,n879);
    nand g6676(n474 ,n407 ,n454);
    nand g6677(n1219 ,n975 ,n743);
    nand g6678(n6409 ,n6278 ,n6336);
    nand g6679(n3292 ,n3285 ,n3263);
    or g6680(n2987 ,n2956 ,n2961);
    nand g6681(n3546 ,n3460 ,n3485);
    xor g6682(n4919 ,n4693 ,n4626);
    nand g6683(n2019 ,n1982 ,n2002);
    or g6684(n6048 ,n5967 ,n6007);
    nand g6685(n3999 ,n3839 ,n3924);
    nand g6686(n6152 ,n6017 ,n6132);
    nand g6687(n898 ,n24[5] ,n715);
    xnor g6688(n4143 ,n4058 ,n4081);
    nand g6689(n3803 ,n3614 ,n3704);
    xnor g6690(n6037 ,n5963 ,n5884);
    nor g6691(n3348 ,n6575 ,n3347);
    nor g6692(n4518 ,n4398 ,n4414);
    nand g6693(n4595 ,n21[2] ,n4363);
    nand g6694(n953 ,n35[15] ,n712);
    nand g6695(n5725 ,n5488 ,n5669);
    nor g6696(n4980 ,n4613 ,n4785);
    nand g6697(n3078 ,n3055 ,n3077);
    nand g6698(n5260 ,n5133 ,n5071);
    nand g6699(n3357 ,n41[4] ,n3356);
    xnor g6700(n2301 ,n2228 ,n2120);
    xnor g6701(n3211 ,n3152 ,n3168);
    or g6702(n775 ,n720 ,n669);
    nand g6703(n242 ,n172 ,n157);
    nor g6704(n6061 ,n5966 ,n6031);
    nor g6705(n2542 ,n2512 ,n2528);
    nand g6706(n2090 ,n6537 ,n2085);
    xnor g6707(n38[6] ,n2507 ,n2534);
    nor g6708(n2662 ,n2568 ,n2590);
    xnor g6709(n2877 ,n2765 ,n2662);
    xnor g6710(n4028 ,n3917 ,n3876);
    xor g6711(n306 ,n209 ,n178);
    nand g6712(n4485 ,n21[1] ,n4373);
    nor g6713(n2028 ,n2020 ,n1993);
    or g6714(n1496 ,n1492 ,n1494);
    xnor g6715(n5199 ,n4901 ,n4961);
    nand g6716(n638 ,n33[1] ,n35[1]);
    nand g6717(n6386 ,n6265 ,n6315);
    nor g6718(n4791 ,n4647 ,n4660);
    xnor g6719(n1800 ,n1743 ,n1648);
    nand g6720(n3644 ,n3481 ,n19[7]);
    not g6721(n5549 ,n5548);
    nor g6722(n3441 ,n3396 ,n3440);
    nand g6723(n5097 ,n4731 ,n5033);
    xnor g6724(n38[8] ,n2524 ,n2548);
    nand g6725(n440 ,n405 ,n411);
    nand g6726(n3731 ,n3590 ,n3528);
    xnor g6727(n2439 ,n2411 ,n2376);
    xnor g6728(n41[6] ,n6159 ,n6157);
    xnor g6729(n3121 ,n6532 ,n6588);
    xnor g6730(n4105 ,n4008 ,n3909);
    nor g6731(n2640 ,n2566 ,n2586);
    xnor g6732(n510 ,n478 ,n467);
    nor g6733(n2468 ,n2416 ,n2448);
    nand g6734(n1063 ,n1517 ,n716);
    nand g6735(n4305 ,n4247 ,n4284);
    nand g6736(n124 ,n24[2] ,n123);
    not g6737(n2666 ,n2665);
    nand g6738(n2203 ,n2092 ,n2158);
    dff g6739(.RN(n1), .SN(1'b1), .CK(n0), .D(n1473), .Q(n27[4]));
    nor g6740(n2030 ,n1959 ,n2011);
    nand g6741(n3522 ,n3482 ,n19[7]);
    nand g6742(n3718 ,n3509 ,n3534);
    nand g6743(n6413 ,n6281 ,n6370);
    nand g6744(n5098 ,n4770 ,n4993);
    nand g6745(n5900 ,n5803 ,n5827);
    not g6746(n4082 ,n4081);
    nand g6747(n122 ,n24[1] ,n24[0]);
    nand g6748(n921 ,n34[14] ,n717);
    nand g6749(n1007 ,n31[2] ,n720);
    dff g6750(.RN(n1), .SN(1'b1), .CK(n0), .D(n1273), .Q(n1503));
    or g6751(n2825 ,n2737 ,n2788);
    nand g6752(n1033 ,n12[1] ,n711);
    nand g6753(n1169 ,n5[5] ,n713);
    nand g6754(n3253 ,n3206 ,n3252);
    nor g6755(n6481 ,n6392 ,n6471);
    not g6756(n4415 ,n4376);
    nand g6757(n5556 ,n5277 ,n5460);
    or g6758(n347 ,n322 ,n335);
    xor g6759(n6022 ,n5967 ,n5994);
    xnor g6760(n674 ,n21[3] ,n30[3]);
    xnor g6761(n6577 ,n1968 ,n1963);
    nand g6762(n3604 ,n3466 ,n3480);
    nor g6763(n593 ,n19[6] ,n27[6]);
    not g6764(n3277 ,n3276);
    nand g6765(n3576 ,n3481 ,n19[5]);
    nand g6766(n1698 ,n1580 ,n1655);
    xnor g6767(n2860 ,n2751 ,n2702);
    nand g6768(n995 ,n25[2] ,n714);
    buf g6769(n14[5], n10[5]);
    xnor g6770(n3124 ,n6577 ,n6554);
    nor g6771(n2762 ,n2647 ,n2721);
    or g6772(n3838 ,n3531 ,n3781);
    nand g6773(n1032 ,n12[2] ,n555);
    nand g6774(n4637 ,n21[5] ,n4386);
    nand g6775(n845 ,n19[1] ,n714);
    xnor g6776(n3072 ,n3036 ,n3027);
    nand g6777(n3162 ,n3118 ,n3143);
    nand g6778(n657 ,n21[5] ,n30[5]);
    nand g6779(n2878 ,n2775 ,n2819);
    nor g6780(n758 ,n619 ,n720);
    not g6781(n5282 ,n5281);
    or g6782(n3918 ,n3863 ,n3861);
    or g6783(n6200 ,n6188 ,n6194);
    nand g6784(n5145 ,n4706 ,n5025);
    buf g6785(n14[2], n11[2]);
    xnor g6786(n423 ,n359 ,n264);
    not g6787(n4363 ,n4362);
    not g6788(n384 ,n266);
    nand g6789(n1176 ,n29[6] ,n724);
    nor g6790(n5062 ,n4780 ,n4960);
    nor g6791(n2499 ,n2464 ,n2468);
    nand g6792(n6099 ,n6080 ,n6028);
    nand g6793(n6207 ,n6178 ,n6201);
    not g6794(n3263 ,n3262);
    xnor g6795(n2864 ,n2761 ,n2797);
    nor g6796(n1958 ,n1909 ,n1930);
    nand g6797(n1468 ,n1143 ,n1387);
    or g6798(n5331 ,n5201 ,n5204);
    nand g6799(n816 ,n23[7] ,n715);
    xnor g6800(n5223 ,n4931 ,n4468);
    nand g6801(n5386 ,n5193 ,n5192);
    nand g6802(n6135 ,n6124 ,n6090);
    or g6803(n4756 ,n4466 ,n4606);
    xor g6804(n1644 ,n1627 ,n1606);
    nand g6805(n5920 ,n5828 ,n5874);
    xnor g6806(n6146 ,n6086 ,n6116);
    not g6807(n175 ,n37[0]);
    xnor g6808(n5170 ,n4881 ,n4516);
    or g6809(n3094 ,n38[14] ,n6587);
    nor g6810(n1999 ,n1966 ,n1972);
    nand g6811(n5389 ,n5208 ,n5207);
    nand g6812(n3242 ,n3186 ,n3241);
    nand g6813(n5137 ,n4768 ,n5035);
    nand g6814(n637 ,n20[1] ,n28[1]);
    nand g6815(n3383 ,n3341 ,n3382);
    nor g6816(n1789 ,n1748 ,n1747);
    xnor g6817(n1522 ,n530 ,n546);
    nand g6818(n4172 ,n4073 ,n4133);
    not g6819(n1929 ,n1928);
    nor g6820(n2479 ,n2403 ,n2461);
    xnor g6821(n3004 ,n2958 ,n2928);
    nand g6822(n6153 ,n6079 ,n6128);
    nor g6823(n6452 ,n6391 ,n6404);
    dff g6824(.RN(n1), .SN(1'b1), .CK(n0), .D(n1401), .Q(n27[9]));
    xnor g6825(n5698 ,n5550 ,n5537);
    nand g6826(n216 ,n169 ,n150);
    nand g6827(n2198 ,n6536 ,n2150);
    xnor g6828(n1884 ,n1796 ,n1820);
    or g6829(n5921 ,n5828 ,n5874);
    nand g6830(n1418 ,n990 ,n1180);
    not g6831(n4414 ,n4380);
    nand g6832(n5081 ,n4708 ,n4996);
    nand g6833(n5473 ,n5294 ,n5382);
    nand g6834(n646 ,n33[10] ,n35[10]);
    nand g6835(n993 ,n19[6] ,n714);
    dff g6836(.RN(n1), .SN(1'b1), .CK(n0), .D(n1353), .Q(n32[7]));
    xor g6837(n298 ,n235 ,n194);
    buf g6838(n14[3], n11[3]);
    xnor g6839(n5913 ,n5803 ,n5858);
    nand g6840(n1303 ,n1060 ,n808);
    nand g6841(n4864 ,n4580 ,n4499);
    nand g6842(n1320 ,n1076 ,n892);
    nand g6843(n4132 ,n4044 ,n4078);
    not g6844(n3464 ,n3463);
    nand g6845(n489 ,n390 ,n469);
    not g6846(n68 ,n36[1]);
    not g6847(n3461 ,n37[6]);
    nand g6848(n6241 ,n41[4] ,n6596);
    or g6849(n533 ,n517 ,n523);
    xnor g6850(n5165 ,n4907 ,n4676);
    nor g6851(n3827 ,n3644 ,n3739);
    xnor g6852(n2947 ,n2860 ,n2899);
    not g6853(n4533 ,n4532);
    not g6854(n265 ,n264);
    xnor g6855(n3040 ,n3004 ,n2947);
    xnor g6856(n38[9] ,n2523 ,n2551);
    nand g6857(n2319 ,n2153 ,n2271);
    xnor g6858(n5764 ,n5638 ,n5524);
    xnor g6859(n2113 ,n2089 ,n2075);
    nand g6860(n5744 ,n5604 ,n5636);
    nand g6861(n5037 ,n4506 ,n4861);
    xnor g6862(n2119 ,n2102 ,n2087);
    nor g6863(n2881 ,n2796 ,n2850);
    nand g6864(n3243 ,n3201 ,n3242);
    buf g6865(n37[2] ,n1502);
    nor g6866(n4075 ,n4006 ,n4028);
    xor g6867(n2058 ,n2281 ,n2269);
    nand g6868(n5469 ,n5215 ,n5391);
    nand g6869(n5982 ,n5935 ,n5884);
    nand g6870(n6388 ,n6238 ,n6255);
    xnor g6871(n38[13] ,n2535 ,n2559);
    nand g6872(n1083 ,n27[8] ,n718);
    nand g6873(n204 ,n170 ,n146);
    nor g6874(n2397 ,n2333 ,n2381);
    nand g6875(n2629 ,n2582 ,n2581);
    dff g6876(.RN(n1), .SN(1'b1), .CK(n0), .D(n1452), .Q(n33[4]));
    nand g6877(n961 ,n27[11] ,n715);
    nand g6878(n1183 ,n29[2] ,n724);
    nor g6879(n209 ,n173 ,n176);
    nand g6880(n4633 ,n4386 ,n20[1]);
    nand g6881(n4825 ,n4477 ,n4640);
    xor g6882(n39[6] ,n38[6] ,n6612);
    buf g6883(n15[1], n15[5]);
    xnor g6884(n2013 ,n1967 ,n1951);
    nand g6885(n5685 ,n5505 ,n5556);
    nor g6886(n6449 ,n6395 ,n6393);
    xor g6887(n4359 ,n5771 ,n5579);
    xnor g6888(n5439 ,n5163 ,n5131);
    nand g6889(n1381 ,n625 ,n766);
    nand g6890(n3202 ,n3157 ,n3172);
    xnor g6891(n2308 ,n2251 ,n2119);
    dff g6892(.RN(n1), .SN(1'b1), .CK(n0), .D(n1222), .Q(n28[2]));
    or g6893(n6040 ,n5991 ,n6003);
    nand g6894(n1027 ,n12[4] ,n710);
    nor g6895(n4544 ,n4405 ,n4399);
    nand g6896(n210 ,n170 ,n153);
    nand g6897(n2189 ,n6538 ,n2148);
    xnor g6898(n671 ,n21[4] ,n30[4]);
    xor g6899(n3949 ,n3862 ,n3870);
    or g6900(n3665 ,n3601 ,n3582);
    xnor g6901(n5618 ,n5434 ,n5079);
    nor g6902(n3862 ,n3669 ,n3817);
    nand g6903(n1149 ,n23[14] ,n716);
    nor g6904(n2055 ,n2014 ,n2054);
    xnor g6905(n3412 ,n6544 ,n6559);
    nand g6906(n1854 ,n1828 ,n1806);
    nor g6907(n2798 ,n2610 ,n2710);
    nand g6908(n5813 ,n5681 ,n5709);
    or g6909(n3920 ,n3842 ,n3859);
    nand g6910(n4157 ,n4085 ,n4123);
    xnor g6911(n2874 ,n2764 ,n2769);
    nand g6912(n3722 ,n3515 ,n3600);
    nand g6913(n6421 ,n6351 ,n6348);
    nand g6914(n3146 ,n6583 ,n3101);
    nand g6915(n6332 ,n39[0] ,n6248);
    nand g6916(n5567 ,n5498 ,n5496);
endmodule
