module top (n0, n1, n6, n7, n2, n3, n8, n4, n5, n9, n10, n12, n13, n11, n14, n15, n16, n17, n18, n20, n19);
    input n0, n1, n2, n3, n4, n5;
    input [31:0] n6, n7, n8;
    output [31:0] n9, n10, n11;
    output n12, n13, n14, n15, n16, n17;
    output [7:0] n18, n19;
    output [15:0] n20;
    wire n0, n1, n2, n3, n4, n5;
    wire [31:0] n6, n7, n8;
    wire [31:0] n9, n10, n11;
    wire n12, n13, n14, n15, n16, n17;
    wire [7:0] n18, n19;
    wire [15:0] n20;
    wire [31:0] n21;
    wire [31:0] n22;
    wire [31:0] n23;
    wire [31:0] n24;
    wire [31:0] n25;
    wire [31:0] n26;
    wire [31:0] n27;
    wire [31:0] n28;
    wire [25:0] n29;
    wire [25:0] n30;
    wire [25:0] n31;
    wire [25:0] n32;
    wire [2:0] n33;
    wire [15:0] n34;
    wire [15:0] n35;
    wire [2:0] n36;
    wire [1:0] n37;
    wire n38, n39, n40, n41, n42, n43, n44, n45;
    wire n46, n47, n48, n49, n50, n51, n52, n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171, n172, n173;
    wire n174, n175, n176, n177, n178, n179, n180, n181;
    wire n182, n183, n184, n185, n186, n187, n188, n189;
    wire n190, n191, n192, n193, n194, n195, n196, n197;
    wire n198, n199, n200, n201, n202, n203, n204, n205;
    wire n206, n207, n208, n209, n210, n211, n212, n213;
    wire n214, n215, n216, n217, n218, n219, n220, n221;
    wire n222, n223, n224, n225, n226, n227, n228, n229;
    wire n230, n231, n232, n233, n234, n235, n236, n237;
    wire n238, n239, n240, n241, n242, n243, n244, n245;
    wire n246, n247, n248, n249, n250, n251, n252, n253;
    wire n254, n255, n256, n257, n258, n259, n260, n261;
    wire n262, n263, n264, n265, n266, n267, n268, n269;
    wire n270, n271, n272, n273, n274, n275, n276, n277;
    wire n278, n279, n280, n281, n282, n283, n284, n285;
    wire n286, n287, n288, n289, n290, n291, n292, n293;
    wire n294, n295, n296, n297, n298, n299, n300, n301;
    wire n302, n303, n304, n305, n306, n307, n308, n309;
    wire n310, n311, n312, n313, n314, n315, n316, n317;
    wire n318, n319, n320, n321, n322, n323, n324, n325;
    wire n326, n327, n328, n329, n330, n331, n332, n333;
    wire n334, n335, n336, n337, n338, n339, n340, n341;
    wire n342, n343, n344, n345, n346, n347, n348, n349;
    wire n350, n351, n352, n353, n354, n355, n356, n357;
    wire n358, n359, n360, n361, n362, n363, n364, n365;
    wire n366, n367, n368, n369, n370, n371, n372, n373;
    wire n374, n375, n376, n377, n378, n379, n380, n381;
    wire n382, n383, n384, n385, n386, n387, n388, n389;
    wire n390, n391, n392, n393, n394, n395, n396, n397;
    wire n398, n399, n400, n401, n402, n403, n404, n405;
    wire n406, n407, n408, n409, n410, n411, n412, n413;
    wire n414, n415, n416, n417, n418, n419, n420, n421;
    wire n422, n423, n424, n425, n426, n427, n428, n429;
    wire n430, n431, n432, n433, n434, n435, n436, n437;
    wire n438, n439, n440, n441, n442, n443, n444, n445;
    wire n446, n447, n448, n449, n450, n451, n452, n453;
    wire n454, n455, n456, n457, n458, n459, n460, n461;
    wire n462, n463, n464, n465, n466, n467, n468, n469;
    wire n470, n471, n472, n473, n474, n475, n476, n477;
    wire n478, n479, n480, n481, n482, n483, n484, n485;
    wire n486, n487, n488, n489, n490, n491, n492, n493;
    wire n494, n495, n496, n497, n498, n499, n500, n501;
    wire n502, n503, n504, n505, n506, n507, n508, n509;
    wire n510, n511, n512, n513, n514, n515, n516, n517;
    wire n518, n519, n520, n521, n522, n523, n524, n525;
    wire n526, n527, n528, n529, n530, n531, n532, n533;
    wire n534, n535, n536, n537, n538, n539, n540, n541;
    wire n542, n543, n544, n545, n546, n547, n548, n549;
    wire n550, n551, n552, n553, n554, n555, n556, n557;
    wire n558, n559, n560, n561, n562, n563, n564, n565;
    wire n566, n567, n568, n569, n570, n571, n572, n573;
    wire n574, n575, n576, n577, n578, n579, n580, n581;
    wire n582, n583, n584, n585, n586, n587, n588, n589;
    wire n590, n591, n592, n593, n594, n595, n596, n597;
    wire n598, n599, n600, n601, n602, n603, n604, n605;
    wire n606, n607, n608, n609, n610, n611, n612, n613;
    wire n614, n615, n616, n617, n618, n619, n620, n621;
    wire n622, n623, n624, n625, n626, n627, n628, n629;
    wire n630, n631, n632, n633, n634, n635, n636, n637;
    wire n638, n639, n640, n641, n642, n643, n644, n645;
    wire n646, n647, n648, n649, n650, n651, n652, n653;
    wire n654, n655, n656, n657, n658, n659, n660, n661;
    wire n662, n663, n664, n665, n666, n667, n668, n669;
    wire n670, n671, n672, n673, n674, n675, n676, n677;
    wire n678, n679, n680, n681, n682, n683, n684, n685;
    wire n686, n687, n688, n689, n690, n691, n692, n693;
    wire n694, n695, n696, n697, n698, n699, n700, n701;
    wire n702, n703, n704, n705, n706, n707, n708, n709;
    wire n710, n711, n712, n713, n714, n715, n716, n717;
    wire n718, n719, n720, n721, n722, n723, n724, n725;
    wire n726, n727, n728, n729, n730, n731, n732, n733;
    wire n734, n735, n736, n737, n738, n739, n740, n741;
    wire n742, n743, n744, n745, n746, n747, n748, n749;
    wire n750, n751, n752, n753, n754, n755, n756, n757;
    wire n758, n759, n760, n761, n762, n763, n764, n765;
    wire n766, n767, n768, n769, n770, n771, n772, n773;
    wire n774, n775, n776, n777, n778, n779, n780, n781;
    wire n782, n783, n784, n785, n786, n787, n788, n789;
    wire n790, n791, n792, n793, n794, n795, n796, n797;
    wire n798, n799, n800, n801, n802, n803, n804, n805;
    wire n806, n807, n808, n809, n810, n811, n812, n813;
    wire n814, n815, n816, n817, n818, n819, n820, n821;
    wire n822, n823, n824, n825, n826, n827, n828, n829;
    wire n830, n831, n832, n833, n834, n835, n836, n837;
    wire n838, n839, n840, n841, n842, n843, n844, n845;
    wire n846, n847, n848, n849, n850, n851, n852, n853;
    wire n854, n855, n856, n857, n858, n859, n860, n861;
    wire n862, n863, n864, n865, n866, n867, n868, n869;
    wire n870, n871, n872, n873, n874, n875, n876, n877;
    wire n878, n879, n880, n881, n882, n883, n884, n885;
    wire n886, n887, n888, n889, n890, n891, n892, n893;
    wire n894, n895, n896, n897, n898, n899, n900, n901;
    wire n902, n903, n904, n905, n906, n907, n908, n909;
    wire n910, n911, n912, n913, n914, n915, n916, n917;
    wire n918, n919, n920, n921, n922, n923, n924, n925;
    wire n926, n927, n928, n929, n930, n931, n932, n933;
    wire n934, n935, n936, n937, n938, n939, n940, n941;
    wire n942, n943, n944, n945, n946, n947, n948, n949;
    wire n950, n951, n952, n953, n954, n955, n956, n957;
    wire n958, n959, n960, n961, n962, n963, n964, n965;
    wire n966, n967, n968, n969, n970, n971, n972, n973;
    wire n974, n975, n976, n977, n978, n979, n980, n981;
    wire n982, n983, n984, n985, n986, n987, n988, n989;
    wire n990, n991, n992, n993, n994, n995, n996, n997;
    wire n998, n999, n1000, n1001, n1002, n1003, n1004, n1005;
    wire n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013;
    wire n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
    wire n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
    wire n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
    wire n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;
    wire n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053;
    wire n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061;
    wire n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069;
    wire n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077;
    wire n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085;
    wire n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093;
    wire n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101;
    wire n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109;
    wire n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117;
    wire n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125;
    wire n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133;
    wire n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141;
    wire n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149;
    wire n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157;
    wire n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165;
    wire n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173;
    wire n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181;
    wire n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189;
    wire n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197;
    wire n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205;
    wire n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
    wire n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221;
    wire n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229;
    wire n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237;
    wire n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245;
    wire n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253;
    wire n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261;
    wire n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269;
    wire n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277;
    wire n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285;
    wire n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293;
    wire n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301;
    wire n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309;
    wire n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;
    wire n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325;
    wire n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333;
    wire n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;
    wire n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349;
    wire n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;
    wire n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365;
    wire n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373;
    wire n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381;
    wire n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389;
    wire n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397;
    wire n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405;
    wire n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413;
    wire n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421;
    wire n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429;
    wire n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437;
    wire n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445;
    wire n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453;
    wire n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461;
    wire n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469;
    wire n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477;
    wire n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485;
    wire n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493;
    wire n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501;
    wire n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509;
    wire n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517;
    wire n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525;
    wire n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533;
    wire n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541;
    wire n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
    wire n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557;
    wire n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565;
    wire n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573;
    wire n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581;
    wire n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589;
    wire n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597;
    wire n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605;
    wire n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613;
    wire n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621;
    wire n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629;
    wire n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637;
    wire n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645;
    wire n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653;
    wire n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661;
    wire n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669;
    wire n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677;
    wire n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685;
    wire n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693;
    wire n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701;
    wire n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709;
    wire n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717;
    wire n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725;
    wire n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733;
    wire n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741;
    wire n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749;
    wire n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757;
    wire n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765;
    wire n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773;
    wire n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781;
    wire n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789;
    wire n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797;
    wire n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805;
    wire n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813;
    wire n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821;
    wire n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829;
    wire n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837;
    wire n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845;
    wire n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853;
    wire n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861;
    wire n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869;
    wire n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877;
    wire n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885;
    wire n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893;
    wire n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901;
    wire n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909;
    wire n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917;
    wire n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925;
    wire n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933;
    wire n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941;
    wire n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949;
    wire n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957;
    wire n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965;
    wire n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973;
    wire n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981;
    wire n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989;
    wire n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997;
    wire n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005;
    wire n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013;
    wire n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021;
    wire n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029;
    wire n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037;
    wire n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045;
    wire n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053;
    wire n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061;
    wire n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069;
    wire n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077;
    wire n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085;
    wire n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093;
    wire n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101;
    wire n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109;
    wire n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117;
    wire n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125;
    wire n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133;
    wire n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141;
    wire n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149;
    wire n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157;
    wire n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165;
    wire n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173;
    wire n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181;
    wire n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189;
    wire n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197;
    wire n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205;
    wire n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213;
    wire n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221;
    wire n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229;
    wire n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237;
    wire n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245;
    wire n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253;
    wire n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261;
    wire n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269;
    wire n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277;
    wire n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285;
    wire n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293;
    wire n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301;
    wire n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309;
    wire n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317;
    wire n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325;
    wire n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333;
    wire n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341;
    wire n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349;
    wire n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357;
    wire n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365;
    wire n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373;
    wire n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381;
    wire n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389;
    wire n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397;
    wire n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405;
    wire n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413;
    wire n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421;
    wire n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429;
    wire n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437;
    wire n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445;
    wire n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453;
    wire n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461;
    wire n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469;
    wire n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477;
    wire n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485;
    wire n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493;
    wire n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501;
    wire n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509;
    wire n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517;
    wire n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525;
    wire n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533;
    wire n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541;
    wire n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549;
    wire n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557;
    wire n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565;
    wire n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573;
    wire n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581;
    wire n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589;
    wire n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597;
    wire n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605;
    wire n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613;
    wire n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621;
    wire n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629;
    wire n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637;
    wire n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645;
    wire n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653;
    wire n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661;
    wire n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669;
    wire n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677;
    wire n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685;
    wire n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693;
    wire n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701;
    wire n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709;
    wire n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717;
    wire n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725;
    wire n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733;
    wire n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741;
    wire n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749;
    wire n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757;
    wire n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765;
    wire n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773;
    wire n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781;
    wire n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789;
    wire n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797;
    wire n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805;
    wire n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813;
    wire n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821;
    wire n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829;
    wire n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837;
    wire n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845;
    wire n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853;
    wire n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861;
    wire n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869;
    wire n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877;
    wire n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885;
    wire n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893;
    wire n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901;
    wire n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909;
    wire n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917;
    wire n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925;
    wire n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933;
    wire n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941;
    wire n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949;
    wire n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957;
    wire n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965;
    wire n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973;
    wire n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981;
    wire n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989;
    wire n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997;
    wire n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005;
    wire n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013;
    wire n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021;
    wire n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029;
    wire n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037;
    wire n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045;
    wire n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053;
    wire n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061;
    wire n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069;
    wire n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077;
    wire n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085;
    wire n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093;
    wire n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101;
    wire n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109;
    wire n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117;
    wire n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125;
    wire n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133;
    wire n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141;
    wire n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149;
    wire n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157;
    wire n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165;
    wire n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173;
    wire n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181;
    wire n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189;
    wire n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197;
    wire n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205;
    wire n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213;
    wire n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221;
    wire n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229;
    wire n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237;
    wire n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245;
    wire n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253;
    wire n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261;
    wire n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269;
    wire n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277;
    wire n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285;
    wire n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293;
    wire n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301;
    wire n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309;
    wire n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317;
    wire n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325;
    wire n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333;
    wire n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341;
    wire n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349;
    wire n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357;
    wire n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365;
    wire n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373;
    wire n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381;
    wire n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389;
    wire n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397;
    wire n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405;
    wire n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413;
    wire n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421;
    wire n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429;
    wire n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437;
    wire n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445;
    wire n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453;
    wire n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461;
    wire n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469;
    wire n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477;
    wire n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485;
    wire n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493;
    wire n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501;
    wire n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509;
    wire n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517;
    wire n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525;
    wire n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533;
    wire n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541;
    wire n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549;
    wire n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557;
    wire n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565;
    wire n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573;
    wire n3574, n3575, n3576, n3577, n3578;
    nand g0(n438 ,n3399 ,n358);
    nor g1(n461 ,n442 ,n413);
    nand g2(n2180 ,n32[21] ,n1462);
    nand g3(n1963 ,n1318 ,n1486);
    nor g4(n3076 ,n2920 ,n3034);
    dff g5(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3097), .Q(n10[22]));
    dff g6(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2010), .Q(n29[25]));
    nand g7(n2990 ,n9[25] ,n2848);
    not g8(n3220 ,n3222);
    nor g9(n1464 ,n539 ,n531);
    nor g10(n1065 ,n694 ,n1027);
    nand g11(n2287 ,n24[27] ,n1950);
    nand g12(n1293 ,n6[24] ,n530);
    nand g13(n3205 ,n3008 ,n3163);
    nand g14(n2434 ,n2191 ,n1737);
    nand g15(n1090 ,n1029 ,n1045);
    nand g16(n3199 ,n2918 ,n3049);
    nand g17(n3101 ,n2788 ,n2940);
    nand g18(n1858 ,n3513 ,n537);
    not g19(n2416 ,n2415);
    nand g20(n2187 ,n32[16] ,n1462);
    not g21(n118 ,n117);
    nor g22(n666 ,n560 ,n29[3]);
    nor g23(n3060 ,n2743 ,n3047);
    nand g24(n120 ,n23[2] ,n118);
    nor g25(n429 ,n382 ,n3401);
    not g26(n587 ,n34[1]);
    nor g27(n2911 ,n997 ,n2691);
    not g28(n2744 ,n2711);
    nand g29(n2114 ,n1428 ,n1623);
    nand g30(n2872 ,n1082 ,n2666);
    nand g31(n964 ,n792 ,n728);
    or g32(n1011 ,n984 ,n946);
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2370), .Q(n22[27]));
    nand g34(n2068 ,n1453 ,n1564);
    nand g35(n2124 ,n1433 ,n1652);
    nand g36(n2884 ,n1225 ,n2678);
    nor g37(n441 ,n373 ,n3400);
    nand g38(n2774 ,n10[31] ,n525);
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2113), .Q(n25[29]));
    or g40(n654 ,n548 ,n29[25]);
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2468), .Q(n30[16]));
    not g42(n845 ,n844);
    nand g43(n1779 ,n3445 ,n535);
    nand g44(n2809 ,n998 ,n2692);
    nand g45(n2296 ,n24[18] ,n1950);
    nor g46(n3356 ,n59 ,n61);
    nand g47(n2553 ,n1777 ,n2253);
    nor g48(n938 ,n614 ,n607);
    nor g49(n597 ,n26[31] ,n6[5]);
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2329), .Q(n30[8]));
    nand g51(n1977 ,n1336 ,n1271);
    nor g52(n397 ,n370 ,n3422);
    not g53(n193 ,n192);
    not g54(n239 ,n238);
    nor g55(n420 ,n357 ,n3432);
    nand g56(n2829 ,n1004 ,n2692);
    nand g57(n815 ,n32[2] ,n565);
    not g58(n171 ,n170);
    nand g59(n987 ,n781 ,n740);
    nand g60(n1187 ,n993 ,n1033);
    nand g61(n1260 ,n6[23] ,n530);
    nand g62(n1059 ,n92 ,n949);
    not g63(n319 ,n318);
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2406), .Q(n23[28]));
    nand g65(n492 ,n427 ,n491);
    nand g66(n2440 ,n2182 ,n1939);
    nand g67(n3032 ,n2725 ,n2763);
    nand g68(n2014 ,n1418 ,n1289);
    nand g69(n1723 ,n6[20] ,n537);
    nand g70(n2620 ,n2563 ,n2610);
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2532), .Q(n21[7]));
    nand g72(n1266 ,n6[16] ,n530);
    not g73(n833 ,n832);
    nand g74(n1660 ,n3562 ,n533);
    nor g75(n616 ,n538 ,n28[26]);
    nor g76(n1009 ,n921 ,n920);
    nor g77(n2980 ,n560 ,n2850);
    nand g78(n2036 ,n1367 ,n1276);
    nor g79(n3159 ,n2227 ,n3132);
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3139), .Q(n9[1]));
    nand g81(n1452 ,n29[25] ,n521);
    nand g82(n1531 ,n1138 ,n1153);
    nor g83(n2655 ,n2605 ,n2626);
    xnor g84(n3449 ,n332 ,n21[23]);
    nand g85(n236 ,n22[2] ,n234);
    nand g86(n2633 ,n859 ,n2610);
    nand g87(n3268 ,n23[2] ,n3222);
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2112), .Q(n25[30]));
    nand g89(n2792 ,n10[13] ,n525);
    nand g90(n1109 ,n27[1] ,n1031);
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2378), .Q(n22[20]));
    nand g92(n1798 ,n8[9] ,n536);
    nand g93(n1815 ,n8[5] ,n536);
    nand g94(n1611 ,n3493 ,n531);
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2454), .Q(n28[12]));
    xnor g96(n899 ,n6[16] ,n29[10]);
    nand g97(n2979 ,n6[10] ,n2849);
    nand g98(n1133 ,n31[24] ,n1031);
    xnor g99(n3464 ,n304 ,n21[8]);
    nand g100(n3294 ,n3221 ,n21[17]);
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n833), .Q(n20[4]));
    nor g102(n475 ,n454 ,n473);
    not g103(n151 ,n150);
    nand g104(n2041 ,n1363 ,n1304);
    nand g105(n3388 ,n3348 ,n3282);
    not g106(n2213 ,n2058);
    nand g107(n2365 ,n1544 ,n1808);
    nand g108(n2118 ,n1432 ,n1639);
    nand g109(n2129 ,n1441 ,n1668);
    nand g110(n2698 ,n7[5] ,n2642);
    nand g111(n2861 ,n25[3] ,n2696);
    nand g112(n1096 ,n1040 ,n1009);
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3190), .Q(n11[20]));
    nand g114(n1884 ,n23[27] ,n1465);
    nand g115(n965 ,n799 ,n780);
    nand g116(n704 ,n32[21] ,n555);
    not g117(n203 ,n202);
    nor g118(n64 ,n48 ,n62);
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2499), .Q(n24[30]));
    nand g120(n1456 ,n25[7] ,n1147);
    nand g121(n2105 ,n26[5] ,n1463);
    nand g122(n1683 ,n8[3] ,n532);
    nand g123(n1994 ,n30[13] ,n1463);
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2441), .Q(n32[18]));
    not g125(n552 ,n6[10]);
    nand g126(n2044 ,n1370 ,n1288);
    nand g127(n1729 ,n6[27] ,n535);
    nand g128(n2783 ,n10[22] ,n2690);
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2365), .Q(n22[31]));
    nand g130(n2168 ,n28[12] ,n1462);
    nor g131(n2607 ,n3565 ,n2600);
    nand g132(n1361 ,n29[9] ,n1147);
    nand g133(n766 ,n30[15] ,n541);
    nand g134(n3175 ,n2908 ,n3079);
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2418), .Q(n32[2]));
    nand g136(n3422 ,n3313 ,n3248);
    nand g137(n1813 ,n22[27] ,n1464);
    nor g138(n898 ,n33[2] ,n601);
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2338), .Q(n30[21]));
    or g140(n2925 ,n874 ,n2848);
    nand g141(n2559 ,n36[2] ,n2416);
    nor g142(n835 ,n587 ,n539);
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2655), .Q(n34[3]));
    nand g144(n760 ,n26[22] ,n538);
    nand g145(n756 ,n32[17] ,n549);
    nand g146(n2641 ,n2 ,n2608);
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2462), .Q(n28[19]));
    nand g148(n2316 ,n1985 ,n1722);
    nand g149(n1134 ,n27[31] ,n1031);
    or g150(n402 ,n352 ,n3437);
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2374), .Q(n22[23]));
    nand g152(n1983 ,n1342 ,n1275);
    nand g153(n1095 ,n1012 ,n1021);
    not g154(n333 ,n332);
    nor g155(n1019 ,n981 ,n956);
    nand g156(n1731 ,n6[25] ,n534);
    nand g157(n1576 ,n1106 ,n1167);
    nand g158(n2067 ,n1421 ,n1394);
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2385), .Q(n22[15]));
    nand g160(n207 ,n24[16] ,n205);
    nand g161(n2535 ,n1831 ,n2272);
    or g162(n1251 ,n22[0] ,n522);
    nand g163(n1826 ,n22[15] ,n1464);
    nand g164(n3130 ,n1401 ,n2975);
    xnor g165(n3524 ,n192 ,n24[10]);
    nand g166(n182 ,n24[4] ,n181);
    nand g167(n2782 ,n10[23] ,n525);
    nand g168(n116 ,n35[6] ,n115);
    nand g169(n1227 ,n27[14] ,n527);
    nand g170(n2262 ,n21[20] ,n1951);
    nand g171(n2096 ,n26[14] ,n1463);
    nand g172(n2315 ,n1946 ,n1698);
    nand g173(n2400 ,n1616 ,n1844);
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2334), .Q(n30[2]));
    xnor g175(n868 ,n6[14] ,n31[8]);
    nand g176(n2254 ,n21[28] ,n1951);
    nand g177(n1820 ,n22[21] ,n1464);
    nand g178(n2447 ,n2177 ,n1727);
    nand g179(n2423 ,n2200 ,n1744);
    nand g180(n62 ,n6[12] ,n61);
    nand g181(n1602 ,n3483 ,n531);
    nor g182(n1055 ,n865 ,n971);
    nor g183(n3078 ,n2911 ,n3038);
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1958), .Q(n31[19]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3182), .Q(n9[26]));
    nand g186(n3249 ,n23[31] ,n3219);
    nand g187(n2411 ,n1635 ,n1888);
    nand g188(n170 ,n23[28] ,n169);
    nor g189(n3148 ,n2317 ,n3119);
    or g190(n1147 ,n834 ,n1062);
    not g191(n2746 ,n2715);
    nor g192(n657 ,n548 ,n30[25]);
    nor g193(n2937 ,n1562 ,n2880);
    xnor g194(n3532 ,n175 ,n24[2]);
    nor g195(n502 ,n446 ,n501);
    nand g196(n910 ,n631 ,n801);
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2132), .Q(n25[12]));
    nor g198(n1248 ,n1085 ,n1095);
    nor g199(n396 ,n376 ,n3429);
    nand g200(n3295 ,n3221 ,n22[20]);
    nand g201(n1277 ,n6[13] ,n532);
    nand g202(n1483 ,n8[30] ,n530);
    nor g203(n2949 ,n1522 ,n2890);
    not g204(n221 ,n220);
    nand g205(n2490 ,n1646 ,n1897);
    nand g206(n1637 ,n3544 ,n532);
    nand g207(n1222 ,n27[18] ,n527);
    nand g208(n2309 ,n24[5] ,n1950);
    nor g209(n3067 ,n2828 ,n3025);
    not g210(n325 ,n324);
    nor g211(n605 ,n26[8] ,n6[5]);
    nand g212(n1655 ,n3558 ,n533);
    nand g213(n1654 ,n8[21] ,n533);
    nand g214(n854 ,n35[7] ,n1);
    not g215(n548 ,n6[31]);
    nand g216(n431 ,n3416 ,n362);
    not g217(n528 ,n1032);
    nand g218(n2918 ,n25[12] ,n2696);
    nand g219(n3133 ,n1577 ,n2978);
    or g220(n692 ,n562 ,n32[6]);
    nand g221(n2730 ,n11[10] ,n2641);
    nand g222(n2431 ,n2194 ,n1739);
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2038), .Q(n27[0]));
    nand g224(n1711 ,n6[9] ,n536);
    not g225(n135 ,n134);
    nand g226(n2376 ,n2105 ,n1815);
    xnor g227(n866 ,n6[15] ,n31[9]);
    not g228(n386 ,n3417);
    nand g229(n3126 ,n1395 ,n2997);
    nand g230(n1204 ,n25[25] ,n529);
    nand g231(n3436 ,n3314 ,n3246);
    or g232(n1080 ,n940 ,n1034);
    nand g233(n3216 ,n2971 ,n3154);
    nand g234(n774 ,n30[6] ,n562);
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2345), .Q(n26[25]));
    nand g236(n2904 ,n6[1] ,n2697);
    nand g237(n2341 ,n2059 ,n1759);
    nand g238(n2108 ,n26[2] ,n520);
    nand g239(n993 ,n784 ,n707);
    nand g240(n1624 ,n3481 ,n530);
    nand g241(n2097 ,n1356 ,n1295);
    nand g242(n1806 ,n3467 ,n534);
    nand g243(n1332 ,n31[8] ,n1146);
    nand g244(n1283 ,n6[15] ,n532);
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n841), .Q(n20[15]));
    nand g246(n1075 ,n933 ,n1033);
    nand g247(n2851 ,n995 ,n2692);
    nor g248(n404 ,n349 ,n3382);
    nor g249(n453 ,n405 ,n420);
    nand g250(n2066 ,n26[26] ,n1463);
    nand g251(n3238 ,n24[21] ,n3219);
    xnor g252(n3556 ,n132 ,n23[9]);
    nand g253(n3404 ,n3315 ,n3250);
    nand g254(n2469 ,n2144 ,n1918);
    nand g255(n827 ,n32[9] ,n564);
    not g256(n125 ,n124);
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2550), .Q(n21[25]));
    or g258(n885 ,n679 ,n639);
    nor g259(n3574 ,n113 ,n115);
    or g260(n2589 ,n1061 ,n2586);
    nand g261(n2327 ,n2098 ,n1721);
    nand g262(n2674 ,n7[20] ,n2642);
    nand g263(n3189 ,n2832 ,n3068);
    nor g264(n101 ,n34[5] ,n100);
    nand g265(n991 ,n816 ,n775);
    nand g266(n1967 ,n1327 ,n1264);
    not g267(n343 ,n342);
    nand g268(n2442 ,n2183 ,n1731);
    nand g269(n967 ,n735 ,n736);
    nand g270(n3193 ,n2919 ,n3076);
    nand g271(n2985 ,n9[30] ,n2848);
    nor g272(n2628 ,n835 ,n2608);
    nand g273(n2170 ,n28[10] ,n1462);
    nand g274(n326 ,n21[19] ,n325);
    dff g275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2547), .Q(n21[22]));
    nand g276(n1969 ,n1328 ,n1265);
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2579), .Q(n36[2]));
    nor g278(n65 ,n56 ,n62);
    dff g279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1981), .Q(n31[2]));
    not g280(n575 ,n31[0]);
    nand g281(n3115 ,n2802 ,n2954);
    nand g282(n745 ,n31[1] ,n563);
    dff g283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3087), .Q(n10[31]));
    nand g284(n2040 ,n798 ,n1466);
    nand g285(n2253 ,n21[29] ,n1951);
    nand g286(n768 ,n26[19] ,n538);
    nand g287(n2586 ,n886 ,n2581);
    nand g288(n3186 ,n2807 ,n3059);
    or g289(n659 ,n549 ,n29[17]);
    not g290(n103 ,n102);
    nand g291(n1193 ,n25[23] ,n529);
    nand g292(n2018 ,n1477 ,n1518);
    nand g293(n2492 ,n1644 ,n1895);
    nand g294(n3106 ,n2792 ,n2944);
    nand g295(n1195 ,n27[17] ,n1031);
    nand g296(n1480 ,n826 ,n521);
    xnor g297(n3552 ,n140 ,n23[13]);
    xnor g298(n3483 ,n268 ,n22[20]);
    nand g299(n440 ,n3387 ,n378);
    xnor g300(n3515 ,n208 ,n24[19]);
    nand g301(n204 ,n24[15] ,n203);
    or g302(n2230 ,n1619 ,n2088);
    nand g303(n146 ,n23[15] ,n145);
    nand g304(n196 ,n24[11] ,n195);
    nand g305(n3185 ,n2996 ,n3057);
    not g306(n562 ,n6[12]);
    dff g307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1964), .Q(n31[14]));
    nand g308(n912 ,n692 ,n712);
    nand g309(n2371 ,n1598 ,n1814);
    or g310(n1246 ,n965 ,n1100);
    nor g311(n483 ,n474 ,n482);
    nand g312(n1007 ,n810 ,n757);
    nand g313(n1579 ,n1184 ,n1107);
    nor g314(n473 ,n463 ,n468);
    nor g315(n514 ,n486 ,n513);
    nand g316(n1788 ,n3453 ,n534);
    dff g317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2517), .Q(n24[13]));
    nand g318(n832 ,n35[4] ,n1);
    nand g319(n2513 ,n1863 ,n2298);
    nand g320(n1949 ,n22[20] ,n1464);
    nand g321(n1139 ,n1001 ,n1033);
    nor g322(n2571 ,n1574 ,n2249);
    nand g323(n1347 ,n27[15] ,n522);
    nand g324(n2898 ,n1071 ,n2702);
    nand g325(n262 ,n22[15] ,n261);
    not g326(n199 ,n198);
    nor g327(n1465 ,n539 ,n533);
    nand g328(n266 ,n22[18] ,n264);
    dff g329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2650), .Q(n36[1]));
    nand g330(n1372 ,n29[0] ,n1147);
    nand g331(n3397 ,n3300 ,n3247);
    not g332(n247 ,n246);
    nand g333(n3089 ,n2777 ,n2929);
    nand g334(n2202 ,n28[0] ,n523);
    xnor g335(n3357 ,n6[12] ,n60);
    not g336(n353 ,n3440);
    nand g337(n2388 ,n1609 ,n1830);
    xnor g338(n3562 ,n120 ,n23[3]);
    dff g339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3091), .Q(n10[27]));
    nand g340(n2061 ,n26[27] ,n1463);
    not g341(n351 ,n3423);
    nand g342(n3279 ,n23[5] ,n3219);
    nand g343(n1476 ,n25[26] ,n521);
    nand g344(n1973 ,n1332 ,n1268);
    xnor g345(n3555 ,n134 ,n23[10]);
    nor g346(n505 ,n389 ,n504);
    nand g347(n2390 ,n1611 ,n1834);
    xnor g348(n3463 ,n306 ,n21[9]);
    nor g349(n609 ,n538 ,n28[6]);
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n838), .Q(n20[12]));
    not g351(n305 ,n304);
    nor g352(n2941 ,n1512 ,n2884);
    nand g353(n1317 ,n31[19] ,n522);
    nand g354(n2686 ,n7[9] ,n2642);
    nand g355(n1755 ,n22[25] ,n1464);
    nand g356(n1851 ,n3506 ,n537);
    not g357(n829 ,n828);
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1968), .Q(n27[25]));
    or g359(n650 ,n551 ,n30[24]);
    nand g360(n2290 ,n24[24] ,n1950);
    nand g361(n1927 ,n8[18] ,n535);
    nor g362(n2692 ,n2594 ,n2641);
    not g363(n289 ,n288);
    nor g364(n2233 ,n987 ,n1753);
    nand g365(n3257 ,n23[15] ,n3219);
    nand g366(n1402 ,n32[8] ,n1149);
    nand g367(n2369 ,n1596 ,n1812);
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3165), .Q(n9[29]));
    nor g369(n794 ,n590 ,n539);
    dff g370(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2362), .Q(n26[9]));
    nand g371(n1509 ,n1144 ,n1142);
    nand g372(n2764 ,n934 ,n2692);
    nand g373(n958 ,n724 ,n734);
    nand g374(n2472 ,n2140 ,n1915);
    dff g375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2707), .Q(n15));
    nor g376(n2659 ,n2619 ,n2649);
    nand g377(n747 ,n31[21] ,n555);
    nand g378(n2004 ,n1383 ,n1586);
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3177), .Q(n11[4]));
    nand g380(n119 ,n23[17] ,n23[16]);
    nor g381(n498 ,n406 ,n497);
    not g382(n581 ,n27[20]);
    dff g383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3090), .Q(n10[29]));
    nand g384(n2366 ,n1594 ,n1810);
    dff g385(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n858), .Q(n19[4]));
    not g386(n129 ,n128);
    xnor g387(n3557 ,n130 ,n23[8]);
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2543), .Q(n21[18]));
    nor g389(n2661 ,n2613 ,n2645);
    nand g390(n956 ,n795 ,n758);
    nand g391(n1929 ,n8[16] ,n534);
    nor g392(n489 ,n432 ,n488);
    nor g393(n112 ,n105 ,n111);
    nor g394(n3163 ,n2231 ,n3137);
    nor g395(n1015 ,n982 ,n959);
    nand g396(n1662 ,n3564 ,n533);
    dff g397(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2442), .Q(n32[19]));
    nand g398(n811 ,n28[20] ,n6[5]);
    or g399(n672 ,n541 ,n30[15]);
    dff g400(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2358), .Q(n26[14]));
    xnor g401(n3501 ,n233 ,n22[2]);
    or g402(n633 ,n551 ,n32[24]);
    nor g403(n624 ,n538 ,n28[1]);
    nand g404(n2056 ,n26[29] ,n1463);
    nor g405(n2860 ,n580 ,n2693);
    dff g406(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2449), .Q(n32[24]));
    nand g407(n773 ,n32[4] ,n552);
    nand g408(n1225 ,n27[16] ,n527);
    not g409(n582 ,n25[17]);
    not g410(n229 ,n228);
    dff g411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3199), .Q(n11[12]));
    nand g412(n1330 ,n31[9] ,n1146);
    nand g413(n1795 ,n3459 ,n534);
    nand g414(n2055 ,n1378 ,n1455);
    not g415(n2210 ,n2053);
    nand g416(n2895 ,n1104 ,n2698);
    nand g417(n3194 ,n2910 ,n3078);
    nand g418(n2681 ,n7[13] ,n2642);
    nand g419(n3168 ,n2810 ,n3060);
    dff g420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2663), .Q(n35[2]));
    nand g421(n81 ,n6[23] ,n76);
    dff g422(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2708), .Q(n14));
    nand g423(n1367 ,n29[6] ,n521);
    xnor g424(n3561 ,n122 ,n23[4]);
    nand g425(n1238 ,n999 ,n1033);
    nor g426(n2622 ,n841 ,n2608);
    nand g427(n1639 ,n8[24] ,n532);
    nand g428(n2143 ,n28[26] ,n523);
    nand g429(n2971 ,n6[18] ,n2849);
    xnor g430(n3355 ,n6[10] ,n58);
    dff g431(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3089), .Q(n10[28]));
    dff g432(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2115), .Q(n25[27]));
    nand g433(n2460 ,n2159 ,n1928);
    nand g434(n1898 ,n23[13] ,n1465);
    nand g435(n3172 ,n2841 ,n3071);
    nand g436(n3021 ,n2817 ,n2760);
    xnor g437(n3451 ,n328 ,n21[21]);
    nand g438(n3263 ,n24[1] ,n3219);
    nand g439(n2961 ,n6[28] ,n2849);
    dff g440(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n835), .Q(n20[9]));
    nand g441(n208 ,n24[18] ,n206);
    nor g442(n1024 ,n953 ,n917);
    not g443(n858 ,n857);
    nand g444(n2885 ,n1206 ,n2679);
    not g445(n2215 ,n2078);
    nand g446(n1299 ,n6[24] ,n532);
    nor g447(n59 ,n6[11] ,n57);
    nand g448(n1679 ,n8[7] ,n532);
    nand g449(n2350 ,n2080 ,n1767);
    or g450(n881 ,n673 ,n674);
    dff g451(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2546), .Q(n21[21]));
    nand g452(n232 ,n24[30] ,n231);
    nand g453(n1668 ,n8[15] ,n532);
    not g454(n2691 ,n2692);
    nand g455(n2054 ,n26[30] ,n520);
    nand g456(n1913 ,n8[30] ,n535);
    nand g457(n1312 ,n31[22] ,n1146);
    nand g458(n3124 ,n1390 ,n2968);
    or g459(n394 ,n350 ,n3438);
    nand g460(n415 ,n3412 ,n388);
    nand g461(n3389 ,n3349 ,n3284);
    nand g462(n2987 ,n9[28] ,n2848);
    nand g463(n1549 ,n1137 ,n1216);
    nor g464(n3153 ,n2220 ,n3124);
    nand g465(n1796 ,n3460 ,n534);
    nand g466(n2840 ,n25[18] ,n2696);
    xor g467(n863 ,n6[20] ,n30[14]);
    dff g468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2352), .Q(n26[19]));
    dff g469(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2391), .Q(n22[9]));
    nand g470(n2354 ,n2089 ,n1770);
    nand g471(n2049 ,n1372 ,n1278);
    or g472(n1146 ,n856 ,n1062);
    nand g473(n1460 ,n31[0] ,n522);
    nor g474(n1242 ,n1098 ,n1088);
    not g475(n565 ,n6[8]);
    nand g476(n1736 ,n6[20] ,n534);
    not g477(n355 ,n3426);
    nand g478(n1627 ,n8[25] ,n533);
    nand g479(n1061 ,n896 ,n899);
    or g480(n669 ,n544 ,n32[5]);
    nand g481(n192 ,n24[9] ,n191);
    not g482(n187 ,n186);
    nand g483(n403 ,n3379 ,n384);
    nand g484(n1420 ,n29[13] ,n1147);
    nand g485(n946 ,n696 ,n791);
    dff g486(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2553), .Q(n21[29]));
    nand g487(n1271 ,n6[11] ,n530);
    nand g488(n49 ,n6[7] ,n43);
    dff g489(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2342), .Q(n26[27]));
    nor g490(n2769 ,n929 ,n2691);
    nand g491(n2334 ,n2006 ,n1704);
    nand g492(n268 ,n22[19] ,n267);
    nand g493(n1180 ,n29[25] ,n1032);
    nand g494(n1321 ,n31[16] ,n522);
    nand g495(n1324 ,n31[14] ,n1146);
    nor g496(n942 ,n610 ,n596);
    not g497(n157 ,n156);
    nand g498(n2153 ,n28[21] ,n523);
    nand g499(n1351 ,n29[24] ,n1147);
    nand g500(n3229 ,n24[16] ,n3222);
    nand g501(n162 ,n23[24] ,n161);
    dff g502(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n840), .Q(n20[14]));
    nand g503(n1541 ,n8[0] ,n531);
    nor g504(n510 ,n399 ,n509);
    nand g505(n3040 ,n2733 ,n2907);
    dff g506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3213), .Q(n9[28]));
    nor g507(n592 ,n26[10] ,n6[5]);
    nand g508(n814 ,n28[16] ,n6[5]);
    nor g509(n652 ,n556 ,n29[19]);
    not g510(n313 ,n312);
    nand g511(n1976 ,n1335 ,n1270);
    nand g512(n2123 ,n1434 ,n1657);
    nand g513(n1062 ,n4 ,n945);
    nand g514(n751 ,n30[16] ,n546);
    nor g515(n482 ,n478 ,n477);
    nand g516(n3405 ,n3316 ,n3252);
    nand g517(n3336 ,n3221 ,n22[3]);
    nand g518(n2192 ,n32[12] ,n1462);
    nand g519(n1254 ,n6[31] ,n530);
    nand g520(n2796 ,n10[9] ,n525);
    not g521(n251 ,n250);
    nand g522(n1527 ,n8[5] ,n530);
    nand g523(n2179 ,n28[7] ,n1462);
    dff g524(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n839), .Q(n20[13]));
    nor g525(n148 ,n119 ,n146);
    nand g526(n1993 ,n30[15] ,n1463);
    nand g527(n1586 ,n8[13] ,n530);
    nand g528(n1168 ,n27[8] ,n1031);
    nand g529(n1350 ,n25[4] ,n1147);
    nand g530(n410 ,n3410 ,n385);
    nor g531(n3048 ,n2759 ,n3020);
    nand g532(n2263 ,n21[19] ,n1951);
    nand g533(n2021 ,n1362 ,n1585);
    nor g534(n2945 ,n1517 ,n2888);
    nand g535(n1389 ,n32[16] ,n1149);
    nand g536(n3102 ,n2789 ,n2941);
    nand g537(n2184 ,n32[18] ,n1462);
    nand g538(n1699 ,n6[30] ,n536);
    nand g539(n310 ,n21[10] ,n309);
    nand g540(n2996 ,n9[19] ,n2848);
    nand g541(n3230 ,n24[10] ,n3219);
    nor g542(n679 ,n561 ,n31[7]);
    nand g543(n788 ,n30[4] ,n552);
    nor g544(n1028 ,n876 ,n918);
    nand g545(n818 ,n28[23] ,n6[5]);
    nor g546(n3158 ,n2226 ,n3130);
    nand g547(n1231 ,n27[26] ,n1031);
    nand g548(n1264 ,n6[18] ,n530);
    dff g549(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3216), .Q(n9[18]));
    nand g550(n1556 ,n1141 ,n1235);
    nand g551(n450 ,n3389 ,n368);
    nor g552(n622 ,n538 ,n28[4]);
    not g553(n997 ,n996);
    nand g554(n2000 ,n1386 ,n1521);
    nand g555(n1421 ,n32[13] ,n1149);
    dff g556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n718), .Q(n19[7]));
    nor g557(n2588 ,n2585 ,n2238);
    nand g558(n2008 ,n30[1] ,n520);
    nand g559(n1744 ,n6[12] ,n534);
    nand g560(n1155 ,n31[13] ,n527);
    or g561(n869 ,n666 ,n634);
    nand g562(n2854 ,n994 ,n2692);
    nor g563(n2624 ,n839 ,n2608);
    nand g564(n1670 ,n8[14] ,n532);
    nand g565(n1159 ,n29[10] ,n1032);
    nand g566(n1577 ,n30[5] ,n1150);
    dff g567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3207), .Q(n9[14]));
    not g568(n524 ,n2690);
    nand g569(n2483 ,n1655 ,n1904);
    nand g570(n117 ,n23[1] ,n23[0]);
    dff g571(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2371), .Q(n22[26]));
    dff g572(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2469), .Q(n28[25]));
    nand g573(n2183 ,n32[19] ,n523);
    dff g574(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2356), .Q(n26[13]));
    nand g575(n2491 ,n1645 ,n1896);
    nand g576(n265 ,n22[16] ,n263);
    nand g577(n2775 ,n10[30] ,n2690);
    nand g578(n320 ,n21[15] ,n319);
    dff g579(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2138), .Q(n25[8]));
    nand g580(n2188 ,n32[15] ,n1462);
    nand g581(n1447 ,n25[11] ,n521);
    nand g582(n734 ,n29[2] ,n565);
    nand g583(n2372 ,n1599 ,n1755);
    not g584(n331 ,n330);
    nand g585(n3009 ,n9[6] ,n2848);
    xnor g586(n3558 ,n128 ,n23[7]);
    nor g587(n640 ,n544 ,n31[5]);
    xnor g588(n3472 ,n290 ,n22[31]);
    nor g589(n595 ,n26[14] ,n6[5]);
    or g590(n676 ,n545 ,n31[18]);
    nand g591(n1216 ,n29[20] ,n1032);
    nand g592(n754 ,n26[18] ,n538);
    dff g593(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3115), .Q(n10[3]));
    nand g594(n2048 ,n30[20] ,n1463);
    not g595(n853 ,n852);
    nand g596(n1566 ,n30[11] ,n1150);
    dff g597(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2535), .Q(n21[10]));
    dff g598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3103), .Q(n10[15]));
    nand g599(n1529 ,n1166 ,n1163);
    dff g600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2097), .Q(n29[17]));
    not g601(n173 ,n172);
    nand g602(n1665 ,n8[17] ,n533);
    nand g603(n750 ,n31[24] ,n551);
    nand g604(n1107 ,n25[22] ,n1032);
    nand g605(n1524 ,n1190 ,n1176);
    nand g606(n1632 ,n3539 ,n532);
    nand g607(n1933 ,n8[12] ,n534);
    xnor g608(n3361 ,n6[16] ,n69);
    or g609(n2225 ,n1571 ,n2075);
    xnor g610(n3444 ,n342 ,n21[28]);
    nand g611(n1177 ,n31[2] ,n527);
    nand g612(n2629 ,n842 ,n2609);
    nand g613(n3326 ,n3221 ,n21[2]);
    nand g614(n2361 ,n2119 ,n1791);
    dff g615(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2537), .Q(n21[12]));
    dff g616(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1963), .Q(n27[27]));
    nand g617(n1535 ,n1120 ,n1124);
    nand g618(n1221 ,n27[11] ,n527);
    nand g619(n1582 ,n30[3] ,n1150);
    nand g620(n1821 ,n1310 ,n1294);
    nand g621(n2479 ,n1660 ,n1908);
    nand g622(n2119 ,n26[10] ,n1463);
    nand g623(n968 ,n749 ,n748);
    nand g624(n2481 ,n1658 ,n1906);
    nand g625(n58 ,n6[9] ,n54);
    nand g626(n1640 ,n3546 ,n532);
    nor g627(n673 ,n562 ,n31[6]);
    nand g628(n1590 ,n1182 ,n1181);
    nand g629(n1757 ,n8[30] ,n537);
    not g630(n362 ,n3384);
    nand g631(n1786 ,n3451 ,n534);
    dff g632(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2538), .Q(n21[13]));
    nand g633(n736 ,n31[12] ,n543);
    nand g634(n456 ,n424 ,n425);
    nand g635(n1828 ,n22[14] ,n1464);
    nand g636(n2117 ,n1430 ,n1627);
    nor g637(n446 ,n378 ,n3387);
    nand g638(n114 ,n35[5] ,n112);
    nand g639(n2240 ,n1251 ,n1846);
    nor g640(n840 ,n586 ,n539);
    nand g641(n1428 ,n25[28] ,n1147);
    dff g642(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1974), .Q(n31[7]));
    nand g643(n258 ,n22[13] ,n257);
    nand g644(n1525 ,n30[24] ,n1150);
    nand g645(n3417 ,n3293 ,n3228);
    nor g646(n3578 ,n108 ,n106);
    nand g647(n1768 ,n8[19] ,n536);
    nand g648(n2340 ,n2056 ,n1758);
    nand g649(n256 ,n22[12] ,n255);
    nand g650(n775 ,n26[0] ,n538);
    nand g651(n1807 ,n3471 ,n534);
    nand g652(n2322 ,n1991 ,n1709);
    not g653(n137 ,n136);
    xnor g654(n874 ,n6[5] ,n33[2]);
    nand g655(n2592 ,n1247 ,n2590);
    nand g656(n2554 ,n1779 ,n2255);
    nand g657(n3433 ,n3327 ,n3260);
    dff g658(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2116), .Q(n25[26]));
    nand g659(n3204 ,n3003 ,n3159);
    nor g660(n2963 ,n557 ,n2850);
    xnor g661(n3542 ,n158 ,n23[23]);
    nand g662(n1937 ,n8[8] ,n534);
    nand g663(n3132 ,n1343 ,n2977);
    nand g664(n2435 ,n2189 ,n1736);
    nand g665(n2252 ,n21[30] ,n1951);
    nand g666(n2530 ,n1806 ,n2277);
    nand g667(n1812 ,n22[28] ,n1464);
    nand g668(n1891 ,n23[20] ,n1465);
    nand g669(n1399 ,n3361 ,n1148);
    nand g670(n1608 ,n3489 ,n531);
    dff g671(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2507), .Q(n24[22]));
    nand g672(n2305 ,n24[9] ,n1950);
    nand g673(n3296 ,n3221 ,n21[18]);
    nand g674(n1915 ,n8[28] ,n535);
    nand g675(n2675 ,n7[19] ,n2642);
    dff g676(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2033), .Q(n27[3]));
    nand g677(n980 ,n698 ,n779);
    nand g678(n2404 ,n1628 ,n1881);
    nand g679(n324 ,n21[18] ,n322);
    nand g680(n2276 ,n21[6] ,n1951);
    nand g681(n3036 ,n2916 ,n2917);
    nand g682(n2137 ,n1451 ,n1675);
    nand g683(n1122 ,n29[2] ,n1032);
    nand g684(n1936 ,n8[9] ,n535);
    nand g685(n3129 ,n1570 ,n3000);
    nand g686(n1722 ,n6[31] ,n536);
    nand g687(n2489 ,n1647 ,n1898);
    not g688(n924 ,n925);
    nor g689(n3150 ,n2218 ,n3122);
    or g690(n656 ,n542 ,n30[13]);
    nand g691(n280 ,n22[25] ,n279);
    nand g692(n817 ,n28[11] ,n6[5]);
    nand g693(n3264 ,n24[2] ,n3219);
    nand g694(n1682 ,n8[4] ,n533);
    nand g695(n1896 ,n23[15] ,n1465);
    nand g696(n1431 ,n25[23] ,n1147);
    nand g697(n2917 ,n25[11] ,n2696);
    nor g698(n2664 ,n2616 ,n2648);
    nand g699(n2300 ,n24[14] ,n1950);
    nor g700(n646 ,n546 ,n30[16]);
    nand g701(n1226 ,n25[12] ,n529);
    nor g702(n683 ,n555 ,n29[21]);
    nand g703(n1959 ,n1319 ,n1293);
    nand g704(n2098 ,n30[10] ,n1463);
    nand g705(n511 ,n401 ,n510);
    nand g706(n2278 ,n21[4] ,n1951);
    nand g707(n1500 ,n1220 ,n1080);
    nor g708(n713 ,n576 ,n6[11]);
    nor g709(n653 ,n540 ,n29[0]);
    nand g710(n2355 ,n2092 ,n1771);
    not g711(n66 ,n65);
    nand g712(n2452 ,n2170 ,n1935);
    nand g713(n2833 ,n25[20] ,n2696);
    xnor g714(n3572 ,n35[7] ,n116);
    nand g715(n104 ,n34[6] ,n103);
    nand g716(n1207 ,n25[27] ,n529);
    or g717(n1244 ,n1090 ,n1089);
    nand g718(n3146 ,n2762 ,n3072);
    nand g719(n970 ,n636 ,n710);
    nand g720(n2245 ,n1676 ,n2211);
    nand g721(n126 ,n23[5] ,n125);
    or g722(n873 ,n664 ,n667);
    not g723(n329 ,n328);
    or g724(n651 ,n562 ,n29[6]);
    nand g725(n3203 ,n3005 ,n3161);
    nor g726(n3082 ,n2753 ,n3043);
    nor g727(n602 ,n26[15] ,n6[5]);
    nor g728(n3364 ,n71 ,n73);
    nor g729(n1048 ,n889 ,n976);
    nor g730(n593 ,n26[27] ,n6[5]);
    nand g731(n2992 ,n9[23] ,n2848);
    nor g732(n433 ,n369 ,n3407);
    nand g733(n2181 ,n32[20] ,n523);
    nand g734(n999 ,n814 ,n767);
    dff g735(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3211), .Q(n9[21]));
    dff g736(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3194), .Q(n11[9]));
    dff g737(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2367), .Q(n22[29]));
    nand g738(n1760 ,n8[27] ,n537);
    nor g739(n678 ,n557 ,n32[20]);
    nand g740(n2496 ,n1805 ,n2280);
    nand g741(n792 ,n31[23] ,n553);
    dff g742(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2651), .Q(n34[6]));
    nor g743(n939 ,n616 ,n598);
    nand g744(n1561 ,n1101 ,n1217);
    nand g745(n2640 ,n852 ,n2610);
    nand g746(n1721 ,n6[16] ,n537);
    nand g747(n3392 ,n3291 ,n3227);
    nand g748(n2324 ,n1993 ,n1702);
    nand g749(n2908 ,n27[8] ,n2694);
    nand g750(n1403 ,n3358 ,n1148);
    nand g751(n3206 ,n3009 ,n3164);
    buf g752(n18[5], 1'b0);
    xnor g753(n896 ,n6[29] ,n29[23]);
    nand g754(n793 ,n32[16] ,n546);
    nand g755(n1659 ,n3561 ,n533);
    nor g756(n94 ,n34[1] ,n34[0]);
    nor g757(n3052 ,n2576 ,n2959);
    nand g758(n1769 ,n8[18] ,n536);
    nand g759(n1157 ,n31[11] ,n527);
    nand g760(n308 ,n21[9] ,n307);
    not g761(n283 ,n282);
    nand g762(n2079 ,n32[1] ,n523);
    dff g763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2524), .Q(n24[5]));
    not g764(n529 ,n528);
    nand g765(n2720 ,n11[20] ,n2641);
    nand g766(n1889 ,n23[22] ,n1465);
    nand g767(n2427 ,n2193 ,n1943);
    nand g768(n3403 ,n3312 ,n3281);
    xnor g769(n3546 ,n150 ,n23[19]);
    nand g770(n2877 ,n1188 ,n2671);
    not g771(n554 ,n6[17]);
    nand g772(n290 ,n22[30] ,n289);
    nor g773(n509 ,n397 ,n508);
    nor g774(n2931 ,n1688 ,n2874);
    nand g775(n708 ,n32[13] ,n542);
    dff g776(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3191), .Q(n11[19]));
    nand g777(n2793 ,n10[12] ,n2690);
    nand g778(n1803 ,n3468 ,n534);
    nand g779(n1885 ,n23[26] ,n1465);
    nand g780(n2721 ,n11[19] ,n2641);
    nor g781(n391 ,n368 ,n3389);
    nand g782(n1358 ,n27[5] ,n1146);
    nand g783(n1871 ,n3525 ,n536);
    nand g784(n3118 ,n2805 ,n2957);
    nand g785(n1158 ,n25[24] ,n1032);
    nand g786(n1052 ,n887 ,n904);
    nand g787(n1802 ,n8[7] ,n536);
    dff g788(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2330), .Q(n30[7]));
    nand g789(n2090 ,n1414 ,n1413);
    nand g790(n1121 ,n27[28] ,n527);
    nand g791(n3006 ,n9[9] ,n2848);
    nand g792(n1161 ,n1003 ,n1033);
    xor g793(n3564 ,n23[1] ,n23[0]);
    nand g794(n2821 ,n27[24] ,n2694);
    dff g795(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2555), .Q(n21[30]));
    nand g796(n1537 ,n1109 ,n1068);
    dff g797(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n853), .Q(n20[6]));
    nand g798(n2011 ,n1439 ,n1677);
    nor g799(n2651 ,n2602 ,n2623);
    nand g800(n1106 ,n31[6] ,n1031);
    dff g801(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2409), .Q(n23[25]));
    nand g802(n42 ,n6[6] ,n6[5]);
    nand g803(n1713 ,n6[26] ,n537);
    nor g804(n414 ,n384 ,n3379);
    nand g805(n1209 ,n25[11] ,n1032);
    nand g806(n2391 ,n1663 ,n1835);
    nand g807(n3138 ,n1416 ,n2983);
    dff g808(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3198), .Q(n11[27]));
    nand g809(n727 ,n31[5] ,n544);
    nand g810(n1581 ,n1154 ,n1171);
    nand g811(n2598 ,n937 ,n2595);
    nand g812(n2182 ,n28[6] ,n523);
    nand g813(n2430 ,n2196 ,n1740);
    nand g814(n1475 ,n29[20] ,n1147);
    dff g815(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2036), .Q(n29[6]));
    nand g816(n1213 ,n31[12] ,n527);
    nand g817(n1816 ,n22[24] ,n1464);
    nand g818(n316 ,n21[13] ,n315);
    nand g819(n1902 ,n23[9] ,n1465);
    dff g820(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2476), .Q(n28[31]));
    dff g821(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2533), .Q(n21[8]));
    nand g822(n2197 ,n32[9] ,n1462);
    nand g823(n1144 ,n31[16] ,n527);
    nand g824(n3254 ,n24[13] ,n3222);
    not g825(n2214 ,n2067);
    nand g826(n3402 ,n3310 ,n3245);
    nand g827(n2791 ,n10[14] ,n2690);
    nor g828(n513 ,n479 ,n512);
    dff g829(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3173), .Q(n11[16]));
    dff g830(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2041), .Q(n29[3]));
    nand g831(n1919 ,n8[24] ,n535);
    nand g832(n2532 ,n1801 ,n2275);
    nand g833(n294 ,n21[2] ,n292);
    nand g834(n916 ,n691 ,n773);
    not g835(n54 ,n53);
    nand g836(n3437 ,n3333 ,n3258);
    nand g837(n3246 ,n23[27] ,n3219);
    nand g838(n2458 ,n1987 ,n1718);
    not g839(n1033 ,n1034);
    nand g840(n2665 ,n7[29] ,n2642);
    nand g841(n318 ,n21[14] ,n317);
    nand g842(n2302 ,n24[12] ,n1950);
    dff g843(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2465), .Q(n28[22]));
    nand g844(n2799 ,n10[6] ,n2690);
    xnor g845(n3466 ,n300 ,n21[6]);
    nand g846(n1473 ,n3373 ,n1148);
    nand g847(n1868 ,n22[17] ,n1464);
    dff g848(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3195), .Q(n11[7]));
    nand g849(n2159 ,n28[17] ,n523);
    nor g850(n2935 ,n1579 ,n2878);
    dff g851(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2505), .Q(n24[24]));
    nand g852(n2540 ,n1793 ,n2267);
    dff g853(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1980), .Q(n31[3]));
    nand g854(n2051 ,n26[31] ,n1463);
    nor g855(n490 ,n404 ,n489);
    xnor g856(n897 ,n6[11] ,n29[5]);
    nand g857(n1256 ,n6[28] ,n530);
    xnor g858(n3526 ,n188 ,n24[8]);
    nor g859(n455 ,n390 ,n433);
    nand g860(n786 ,n28[21] ,n6[5]);
    nor g861(n671 ,n550 ,n29[22]);
    dff g862(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2028), .Q(n29[13]));
    dff g863(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2149), .Q(n25[1]));
    not g864(n549 ,n6[23]);
    nor g865(n3080 ,n2906 ,n3040);
    xnor g866(n3575 ,n35[4] ,n111);
    nand g867(n1647 ,n3552 ,n533);
    nand g868(n1573 ,n1102 ,n1164);
    or g869(n702 ,n550 ,n30[22]);
    not g870(n339 ,n338);
    nand g871(n3107 ,n2793 ,n2945);
    nand g872(n1939 ,n8[6] ,n534);
    nand g873(n2531 ,n1819 ,n2276);
    nand g874(n954 ,n756 ,n759);
    nand g875(n3228 ,n23[8] ,n3219);
    nand g876(n911 ,n630 ,n800);
    nand g877(n2332 ,n2026 ,n1717);
    nand g878(n2919 ,n25[13] ,n2696);
    nand g879(n1621 ,n8[18] ,n531);
    nand g880(n1388 ,n3367 ,n1148);
    nand g881(n959 ,n739 ,n714);
    nand g882(n2257 ,n21[25] ,n1951);
    not g883(n121 ,n120);
    dff g884(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2117), .Q(n25[25]));
    nand g885(n2100 ,n26[11] ,n520);
    dff g886(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2049), .Q(n29[0]));
    or g887(n688 ,n541 ,n32[15]);
    nand g888(n2110 ,n26[0] ,n1463);
    nand g889(n1191 ,n29[3] ,n529);
    dff g890(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2316), .Q(n30[25]));
    or g891(n630 ,n556 ,n32[19]);
    nand g892(n2318 ,n1986 ,n1699);
    nand g893(n2425 ,n2199 ,n1743);
    nand g894(n2422 ,n2202 ,n1945);
    dff g895(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2336), .Q(n26[30]));
    nand g896(n336 ,n21[24] ,n335);
    nand g897(n2761 ,n938 ,n2692);
    nand g898(n3276 ,n24[8] ,n3219);
    nand g899(n1228 ,n29[21] ,n1032);
    nand g900(n2666 ,n7[28] ,n2642);
    nand g901(n2196 ,n32[10] ,n1462);
    dff g902(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2401), .Q(n22[1]));
    dff g903(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2118), .Q(n25[24]));
    nand g904(n2842 ,n27[17] ,n2694);
    nand g905(n2733 ,n11[7] ,n2641);
    dff g906(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2380), .Q(n22[18]));
    nand g907(n3213 ,n2987 ,n3149);
    nand g908(n3091 ,n2778 ,n2930);
    nand g909(n2005 ,n30[3] ,n520);
    nand g910(n1360 ,n27[11] ,n1146);
    nand g911(n1175 ,n1004 ,n1033);
    nor g912(n3149 ,n2217 ,n3121);
    nand g913(n1887 ,n23[24] ,n1465);
    nand g914(n1912 ,n8[31] ,n535);
    nand g915(n1311 ,n31[23] ,n522);
    nand g916(n1540 ,n1132 ,n1180);
    nand g917(n2428 ,n2197 ,n1741);
    nand g918(n1578 ,n1169 ,n1145);
    or g919(n2229 ,n1581 ,n2083);
    nand g920(n2037 ,n1344 ,n1286);
    nand g921(n3025 ,n2718 ,n2827);
    dff g922(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3192), .Q(n11[15]));
    nor g923(n1035 ,n539 ,n926);
    dff g924(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2430), .Q(n32[10]));
    nand g925(n2238 ,n1754 ,n1242);
    nand g926(n2966 ,n6[23] ,n2849);
    nand g927(n1370 ,n29[2] ,n521);
    xnor g928(n3573 ,n35[6] ,n114);
    nand g929(n3328 ,n3220 ,n21[3]);
    nand g930(n2409 ,n1633 ,n1886);
    nand g931(n2019 ,n1354 ,n1301);
    nand g932(n2839 ,n1001 ,n2692);
    nand g933(n3300 ,n3220 ,n21[20]);
    not g934(n307 ,n306);
    nand g935(n1630 ,n3537 ,n532);
    nand g936(n3285 ,n23[19] ,n3219);
    nand g937(n2707 ,n1197 ,n2643);
    nand g938(n507 ,n393 ,n506);
    dff g939(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3205), .Q(n9[7]));
    nand g940(n1817 ,n22[23] ,n1464);
    nand g941(n458 ,n409 ,n408);
    nand g942(n2546 ,n1786 ,n2261);
    nand g943(n1705 ,n6[14] ,n536);
    nand g944(n238 ,n22[3] ,n237);
    nor g945(n2759 ,n940 ,n2691);
    nor g946(n927 ,n624 ,n606);
    nand g947(n2871 ,n1074 ,n2665);
    nor g948(n3051 ,n2769 ,n3041);
    not g949(n2747 ,n2716);
    nand g950(n1322 ,n31[15] ,n1146);
    nand g951(n142 ,n23[13] ,n141);
    nand g952(n2543 ,n1789 ,n2264);
    nand g953(n1235 ,n29[17] ,n1032);
    not g954(n572 ,n34[4]);
    nand g955(n755 ,n31[13] ,n542);
    nand g956(n2503 ,n1853 ,n2288);
    nand g957(n764 ,n30[0] ,n540);
    nor g958(n3351 ,n43 ,n41);
    dff g959(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2660), .Q(n35[5]));
    xnor g960(n3476 ,n282 ,n22[27]);
    nand g961(n1717 ,n6[10] ,n537);
    nand g962(n1071 ,n928 ,n1033);
    nand g963(n2293 ,n24[21] ,n1950);
    dff g964(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2520), .Q(n24[9]));
    nand g965(n1823 ,n22[19] ,n1464);
    dff g966(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2420), .Q(n32[4]));
    xnor g967(n3494 ,n248 ,n22[9]);
    not g968(n147 ,n146);
    nor g969(n664 ,n565 ,n30[2]);
    nand g970(n1532 ,n8[3] ,n530);
    nand g971(n1194 ,n27[10] ,n527);
    dff g972(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2419), .Q(n32[3]));
    nand g973(n2017 ,n1475 ,n1303);
    not g974(n279 ,n278);
    nand g975(n746 ,n31[22] ,n550);
    nand g976(n136 ,n23[10] ,n135);
    nand g977(n178 ,n24[2] ,n176);
    nand g978(n408 ,n3394 ,n355);
    dff g979(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3094), .Q(n10[24]));
    nand g980(n488 ,n418 ,n484);
    xnor g981(n3539 ,n164 ,n23[26]);
    dff g982(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n796), .Q(n33[1]));
    nor g983(n2948 ,n1526 ,n2891);
    nand g984(n2894 ,n1066 ,n2689);
    nand g985(n3243 ,n23[12] ,n3222);
    dff g986(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2339), .Q(n30[20]));
    nand g987(n3047 ,n2808 ,n2809);
    nand g988(n2514 ,n1864 ,n2299);
    nand g989(n2169 ,n28[11] ,n523);
    nand g990(n2673 ,n7[21] ,n2642);
    nor g991(n3055 ,n2574 ,n2964);
    dff g992(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2037), .Q(n29[5]));
    nand g993(n1404 ,n3357 ,n1148);
    nand g994(n2381 ,n1606 ,n1868);
    nor g995(n838 ,n572 ,n539);
    dff g996(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2496), .Q(n21[2]));
    nand g997(n2563 ,n925 ,n2415);
    nand g998(n948 ,n625 ,n741);
    dff g999(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2773), .Q(n13));
    nand g1000(n2401 ,n1617 ,n1845);
    nand g1001(n1384 ,n3368 ,n1148);
    nand g1002(n270 ,n22[20] ,n269);
    nand g1003(n3007 ,n9[8] ,n2848);
    nor g1004(n2601 ,n3571 ,n2600);
    nand g1005(n1862 ,n3517 ,n536);
    or g1006(n1020 ,n716 ,n898);
    nor g1007(n663 ,n565 ,n29[2]);
    nor g1008(n2922 ,n577 ,n2695);
    nand g1009(n2763 ,n935 ,n2692);
    nand g1010(n3034 ,n2727 ,n2765);
    dff g1011(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n855), .Q(n20[7]));
    dff g1012(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2325), .Q(n30[14]));
    not g1013(n526 ,n1031);
    nor g1014(n3374 ,n85 ,n87);
    or g1015(n2227 ,n1576 ,n2081);
    nand g1016(n132 ,n23[8] ,n131);
    nand g1017(n823 ,n92 ,n1);
    not g1018(n2755 ,n2739);
    nand g1019(n1118 ,n1000 ,n1033);
    nand g1020(n1002 ,n811 ,n762);
    xnor g1021(n904 ,n6[13] ,n32[7]);
    nand g1022(n3320 ,n3221 ,n21[30]);
    xor g1023(n3362 ,n6[17] ,n65);
    xnor g1024(n3481 ,n272 ,n22[22]);
    nor g1025(n945 ,n717 ,n719);
    dff g1026(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1972), .Q(n27[24]));
    nand g1027(n1362 ,n27[17] ,n522);
    nand g1028(n1829 ,n22[13] ,n1464);
    dff g1029(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2461), .Q(n28[18]));
    nand g1030(n1279 ,n6[7] ,n532);
    nand g1031(n2306 ,n24[8] ,n1950);
    nand g1032(n2386 ,n1608 ,n1828);
    nand g1033(n3345 ,n3221 ,n22[5]);
    xnor g1034(n3551 ,n142 ,n23[14]);
    nand g1035(n172 ,n23[29] ,n171);
    dff g1036(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2490), .Q(n23[14]));
    nor g1037(n684 ,n550 ,n31[22]);
    nand g1038(n1056 ,n866 ,n892);
    nand g1039(n2010 ,n1452 ,n1302);
    nor g1040(n596 ,n26[29] ,n6[5]);
    or g1041(n631 ,n561 ,n29[7]);
    nand g1042(n2265 ,n21[17] ,n1951);
    nand g1043(n220 ,n24[24] ,n219);
    nand g1044(n2190 ,n28[4] ,n523);
    not g1045(n2648 ,n2637);
    nand g1046(n426 ,n3438 ,n350);
    nand g1047(n3120 ,n2568 ,n2986);
    nand g1048(n1724 ,n6[13] ,n537);
    nand g1049(n809 ,n28[30] ,n6[5]);
    nand g1050(n1741 ,n6[15] ,n534);
    nand g1051(n2175 ,n32[24] ,n1462);
    nand g1052(n1850 ,n3505 ,n537);
    nand g1053(n2085 ,n26[18] ,n520);
    nand g1054(n2519 ,n1870 ,n2304);
    not g1055(n271 ,n270);
    nor g1056(n1013 ,n968 ,n967);
    not g1057(n588 ,n34[7]);
    nand g1058(n782 ,n30[9] ,n564);
    dff g1059(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2528), .Q(n24[1]));
    nand g1060(n1601 ,n3482 ,n531);
    nand g1061(n2845 ,n25[16] ,n2696);
    nand g1062(n2887 ,n1075 ,n2681);
    dff g1063(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n794), .Q(n33[0]));
    nor g1064(n3072 ,n2843 ,n3030);
    nand g1065(n2321 ,n1990 ,n1710);
    nand g1066(n1555 ,n30[17] ,n1150);
    nand g1067(n1749 ,n6[7] ,n535);
    nor g1068(n2595 ,n2594 ,n2591);
    nor g1069(n1149 ,n538 ,n1034);
    nor g1070(n497 ,n436 ,n496);
    nand g1071(n1289 ,n6[28] ,n533);
    nand g1072(n1210 ,n998 ,n1033);
    not g1073(n2212 ,n2057);
    nand g1074(n2865 ,n25[1] ,n2696);
    nand g1075(n1297 ,n6[19] ,n533);
    nor g1076(n1040 ,n863 ,n922);
    or g1077(n2573 ,n1554 ,n2247);
    nand g1078(n2902 ,n6[3] ,n2697);
    nand g1079(n2773 ,n785 ,n2690);
    nand g1080(n3439 ,n3346 ,n3286);
    nor g1081(n944 ,n622 ,n703);
    dff g1082(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2327), .Q(n30[10]));
    nand g1083(n2035 ,n1345 ,n1536);
    nand g1084(n2539 ,n1794 ,n2268);
    dff g1085(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2027), .Q(n27[4]));
    nand g1086(n740 ,n29[9] ,n564);
    nand g1087(n2444 ,n2180 ,n1729);
    nor g1088(n1022 ,n961 ,n980);
    or g1089(n929 ,n609 ,n603);
    nand g1090(n1966 ,n1323 ,n1487);
    or g1091(n932 ,n619 ,n604);
    nand g1092(n200 ,n24[13] ,n199);
    nand g1093(n1596 ,n3475 ,n531);
    nand g1094(n1409 ,n29[12] ,n1147);
    dff g1095(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2508), .Q(n24[21]));
    nand g1096(n1625 ,n8[27] ,n533);
    nand g1097(n3105 ,n2796 ,n2947);
    nand g1098(n1162 ,n31[9] ,n1031);
    dff g1099(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2459), .Q(n28[16]));
    nand g1100(n3191 ,n2839 ,n3070);
    not g1101(n578 ,n25[22]);
    nor g1102(n674 ,n542 ,n31[13]);
    dff g1103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2552), .Q(n21[28]));
    nand g1104(n1709 ,n6[23] ,n536);
    not g1105(n2209 ,n2050);
    nand g1106(n2132 ,n1445 ,n1672);
    nand g1107(n1424 ,n3354 ,n1148);
    nand g1108(n3188 ,n2829 ,n3067);
    nand g1109(n1684 ,n8[2] ,n532);
    not g1110(n3221 ,n3222);
    nand g1111(n3258 ,n23[28] ,n3222);
    nand g1112(n3329 ,n3220 ,n21[4]);
    nand g1113(n2879 ,n1156 ,n2673);
    nand g1114(n3273 ,n23[18] ,n3219);
    nand g1115(n1583 ,n1174 ,n1191);
    nand g1116(n1259 ,n6[25] ,n531);
    nand g1117(n1610 ,n3492 ,n530);
    or g1118(n686 ,n543 ,n29[12]);
    nand g1119(n2271 ,n21[11] ,n1951);
    xnor g1120(n3521 ,n198 ,n24[13]);
    dff g1121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3107), .Q(n10[12]));
    nand g1122(n767 ,n26[16] ,n538);
    nand g1123(n2685 ,n7[10] ,n2642);
    nand g1124(n3020 ,n2713 ,n2815);
    nand g1125(n1830 ,n22[12] ,n1464);
    nand g1126(n757 ,n26[24] ,n538);
    not g1127(n590 ,n36[0]);
    not g1128(n110 ,n109);
    nand g1129(n1849 ,n3504 ,n537);
    dff g1130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3168), .Q(n11[30]));
    nand g1131(n2043 ,n1457 ,n1494);
    dff g1132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3101), .Q(n10[17]));
    or g1133(n2582 ,n901 ,n2566);
    not g1134(n357 ,n3400);
    nand g1135(n1140 ,n31[18] ,n1031);
    or g1136(n687 ,n563 ,n30[1]);
    nand g1137(n2712 ,n11[28] ,n2641);
    nand g1138(n2998 ,n9[17] ,n2848);
    nand g1139(n1506 ,n1185 ,n1161);
    nor g1140(n2947 ,n1524 ,n2892);
    nand g1141(n2558 ,n36[1] ,n2416);
    nand g1142(n3100 ,n2787 ,n2939);
    nand g1143(n1089 ,n1010 ,n1015);
    dff g1144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1979), .Q(n31[4]));
    nand g1145(n3016 ,n2709 ,n2756);
    or g1146(n690 ,n553 ,n32[23]);
    nand g1147(n102 ,n34[5] ,n100);
    nand g1148(n1131 ,n25[0] ,n1032);
    nand g1149(n2643 ,n3 ,n2608);
    nand g1150(n753 ,n31[10] ,n547);
    nand g1151(n765 ,n32[24] ,n551);
    nor g1152(n2942 ,n1513 ,n2885);
    nand g1153(n2360 ,n2100 ,n1784);
    dff g1154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3109), .Q(n10[10]));
    nand g1155(n2798 ,n10[7] ,n525);
    dff g1156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1976), .Q(n31[6]));
    nand g1157(n1777 ,n3443 ,n535);
    dff g1158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2240), .Q(n22[0]));
    xnor g1159(n891 ,n6[7] ,n32[1]);
    xnor g1160(n3376 ,n6[31] ,n88);
    nand g1161(n2160 ,n30[14] ,n520);
    nand g1162(n3262 ,n23[16] ,n3219);
    nand g1163(n2689 ,n7[6] ,n2642);
    nand g1164(n2785 ,n10[20] ,n2690);
    xnor g1165(n3566 ,n34[6] ,n102);
    nand g1166(n70 ,n6[17] ,n65);
    nand g1167(n2500 ,n1852 ,n2287);
    nand g1168(n712 ,n32[19] ,n556);
    nand g1169(n2846 ,n27[16] ,n2694);
    nand g1170(n2242 ,n1525 ,n2208);
    nand g1171(n1198 ,n25[10] ,n529);
    nand g1172(n1739 ,n6[17] ,n534);
    nand g1173(n1771 ,n8[16] ,n536);
    dff g1174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2658), .Q(n35[7]));
    nor g1175(n1466 ,n945 ,n1148);
    nand g1176(n3286 ,n23[30] ,n3219);
    nand g1177(n1346 ,n3374 ,n1148);
    nand g1178(n1725 ,n6[31] ,n534);
    nand g1179(n2367 ,n1595 ,n1811);
    or g1180(n629 ,n565 ,n31[2]);
    not g1181(n527 ,n526);
    dff g1182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n849), .Q(n20[3]));
    dff g1183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1999), .Q(n29[7]));
    nand g1184(n2320 ,n1989 ,n1716);
    not g1185(n215 ,n214);
    nand g1186(n2740 ,n11[21] ,n2641);
    nand g1187(n1436 ,n32[7] ,n1149);
    nand g1188(n857 ,n17 ,n1);
    nor g1189(n442 ,n355 ,n3394);
    nand g1190(n467 ,n438 ,n437);
    nand g1191(n1708 ,n6[6] ,n537);
    nand g1192(n1079 ,n930 ,n1033);
    nand g1193(n2178 ,n32[22] ,n1462);
    nand g1194(n2874 ,n1070 ,n2668);
    or g1195(n3166 ,n2976 ,n3131);
    nor g1196(n3085 ,n2755 ,n3046);
    not g1197(n297 ,n296);
    nand g1198(n3225 ,n23[7] ,n3219);
    nand g1199(n1397 ,n32[11] ,n1149);
    nand g1200(n3396 ,n3299 ,n3235);
    not g1201(n243 ,n242);
    dff g1202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3144), .Q(n11[25]));
    xor g1203(n3368 ,n6[23] ,n76);
    nor g1204(n598 ,n26[26] ,n6[5]);
    or g1205(n665 ,n554 ,n29[11]);
    nand g1206(n1616 ,n3501 ,n531);
    nand g1207(n1163 ,n25[6] ,n529);
    nand g1208(n2900 ,n1103 ,n2704);
    nand g1209(n2449 ,n2175 ,n1726);
    dff g1210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2047), .Q(n29[1]));
    nand g1211(n1510 ,n1202 ,n1223);
    dff g1212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2488), .Q(n23[12]));
    not g1213(n237 ,n236);
    nand g1214(n1747 ,n6[9] ,n534);
    nand g1215(n1710 ,n6[24] ,n537);
    xnor g1216(n3447 ,n336 ,n21[25]);
    nand g1217(n2191 ,n32[13] ,n523);
    nand g1218(n2989 ,n9[26] ,n2848);
    nand g1219(n3196 ,n2861 ,n3084);
    nor g1220(n390 ,n353 ,n3408);
    nor g1221(n3064 ,n2746 ,n3022);
    nand g1222(n1589 ,n30[0] ,n1150);
    nand g1223(n1223 ,n25[19] ,n529);
    nand g1224(n2547 ,n1785 ,n2260);
    nor g1225(n1031 ,n856 ,n924);
    nand g1226(n186 ,n24[6] ,n185);
    not g1227(n381 ,n3425);
    xnor g1228(n3570 ,n34[2] ,n95);
    not g1229(n349 ,n3414);
    nand g1230(n2802 ,n10[3] ,n525);
    nand g1231(n819 ,n28[9] ,n6[5]);
    nand g1232(n2637 ,n846 ,n2610);
    nand g1233(n2858 ,n27[4] ,n2694);
    nand g1234(n2993 ,n9[22] ,n2848);
    nand g1235(n2015 ,n1471 ,n1281);
    not g1236(n571 ,n25[28]);
    nand g1237(n2527 ,n1878 ,n2312);
    nand g1238(n2152 ,n1472 ,n1686);
    xnor g1239(n3480 ,n274 ,n22[23]);
    or g1240(n719 ,n33[0] ,n33[2]);
    dff g1241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2087), .Q(n27[5]));
    nand g1242(n2770 ,n944 ,n2692);
    nand g1243(n1043 ,n908 ,n923);
    not g1244(n131 ,n130);
    nand g1245(n2958 ,n6[31] ,n2849);
    nand g1246(n1268 ,n6[14] ,n531);
    nand g1247(n2125 ,n1437 ,n1664);
    nand g1248(n3265 ,n23[1] ,n3219);
    nor g1249(n2906 ,n570 ,n2695);
    nand g1250(n1548 ,n1136 ,n1228);
    nand g1251(n721 ,n26[30] ,n538);
    nand g1252(n3135 ,n2570 ,n3006);
    not g1253(n2745 ,n2714);
    nand g1254(n2454 ,n2168 ,n1933);
    nand g1255(n2261 ,n21[21] ,n1951);
    nor g1256(n2581 ,n2565 ,n2237);
    nand g1257(n852 ,n35[6] ,n1);
    nand g1258(n1468 ,n25[3] ,n521);
    nand g1259(n2378 ,n1602 ,n1949);
    or g1260(n2218 ,n1556 ,n2060);
    nand g1261(n2029 ,n1409 ,n1305);
    dff g1262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2498), .Q(n24[31]));
    nand g1263(n2311 ,n24[3] ,n1950);
    not g1264(n523 ,n535);
    nand g1265(n346 ,n21[29] ,n345);
    nand g1266(n3013 ,n9[3] ,n2848);
    nand g1267(n1727 ,n6[29] ,n534);
    nand g1268(n812 ,n28[19] ,n6[5]);
    nand g1269(n2284 ,n24[30] ,n1950);
    nand g1270(n1875 ,n3529 ,n536);
    nand g1271(n46 ,n6[10] ,n6[9]);
    dff g1272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2477), .Q(n23[1]));
    nand g1273(n758 ,n32[6] ,n562);
    nand g1274(n2523 ,n1874 ,n2308);
    nand g1275(n2070 ,n1397 ,n1396);
    xnor g1276(n3455 ,n323 ,n21[17]);
    nand g1277(n2370 ,n1597 ,n1813);
    dff g1278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1977), .Q(n31[5]));
    nand g1279(n2672 ,n7[22] ,n2642);
    xnor g1280(n3541 ,n160 ,n23[24]);
    nand g1281(n1917 ,n8[26] ,n535);
    not g1282(n287 ,n286);
    dff g1283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2315), .Q(n32[0]));
    nand g1284(n1692 ,n30[4] ,n1150);
    dff g1285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2125), .Q(n25[18]));
    dff g1286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2639), .Q(n17));
    dff g1287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2664), .Q(n35[1]));
    nand g1288(n1411 ,n32[2] ,n1149);
    nand g1289(n3119 ,n1539 ,n2958);
    not g1290(n384 ,n3411);
    nand g1291(n971 ,n755 ,n753);
    xnor g1292(n888 ,n6[31] ,n31[25]);
    nand g1293(n2521 ,n1872 ,n2306);
    dff g1294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3193), .Q(n11[13]));
    nand g1295(n2817 ,n25[26] ,n2696);
    or g1296(n870 ,n626 ,n678);
    nand g1297(n799 ,n30[20] ,n557);
    nand g1298(n3252 ,n24[28] ,n3219);
    xnor g1299(n3487 ,n262 ,n22[16]);
    nand g1300(n3383 ,n3334 ,n3271);
    nand g1301(n2362 ,n2101 ,n1798);
    nor g1302(n1241 ,n1059 ,n1087);
    nand g1303(n2635 ,n848 ,n2610);
    nand g1304(n1716 ,n6[25] ,n536);
    not g1305(n2632 ,n2625);
    nand g1306(n1280 ,n6[30] ,n532);
    dff g1307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3146), .Q(n11[17]));
    nand g1308(n478 ,n419 ,n472);
    nor g1309(n1083 ,n881 ,n1060);
    nand g1310(n2737 ,n11[3] ,n2641);
    nand g1311(n1514 ,n1227 ,n1229);
    nand g1312(n2072 ,n1387 ,n1621);
    nand g1313(n2807 ,n27[31] ,n2694);
    or g1314(n2219 ,n1509 ,n2062);
    nor g1315(n2590 ,n1093 ,n2587);
    nand g1316(n2995 ,n9[20] ,n2848);
    nand g1317(n1513 ,n1219 ,n1078);
    nand g1318(n1357 ,n29[15] ,n521);
    nor g1319(n448 ,n360 ,n3398);
    nand g1320(n2484 ,n1653 ,n1903);
    nand g1321(n2551 ,n1780 ,n2256);
    nand g1322(n1955 ,n1313 ,n1484);
    nand g1323(n1810 ,n22[30] ,n1464);
    nand g1324(n1341 ,n27[21] ,n522);
    dff g1325(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2422), .Q(n28[0]));
    nand g1326(n332 ,n21[22] ,n331);
    nand g1327(n1922 ,n8[22] ,n535);
    nand g1328(n1217 ,n29[14] ,n1032);
    nand g1329(n1615 ,n3499 ,n531);
    nand g1330(n3313 ,n3220 ,n22[13]);
    nand g1331(n741 ,n30[2] ,n565);
    nand g1332(n2268 ,n21[14] ,n1951);
    dff g1333(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2421), .Q(n32[5]));
    dff g1334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n831), .Q(n19[5]));
    nand g1335(n328 ,n21[20] ,n327);
    nand g1336(n1501 ,n1115 ,n1118);
    nand g1337(n128 ,n23[6] ,n127);
    nor g1338(n3061 ,n2744 ,n3018);
    dff g1339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2544), .Q(n21[19]));
    nand g1340(n3235 ,n24[19] ,n3219);
    dff g1341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3204), .Q(n9[12]));
    nand g1342(n714 ,n29[0] ,n540);
    xnor g1343(n3508 ,n222 ,n24[26]);
    nand g1344(n1261 ,n6[22] ,n530);
    nor g1345(n2654 ,n2604 ,n2630);
    nor g1346(n623 ,n538 ,n28[2]);
    nand g1347(n69 ,n6[15] ,n64);
    nand g1348(n1857 ,n3512 ,n537);
    dff g1349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2341), .Q(n26[28]));
    nand g1350(n1141 ,n31[17] ,n1031);
    nand g1351(n2890 ,n1076 ,n2685);
    nand g1352(n1084 ,n1020 ,n1025);
    nand g1353(n1338 ,n27[22] ,n1146);
    nand g1354(n1479 ,n824 ,n522);
    nand g1355(n2121 ,n1423 ,n1650);
    nand g1356(n111 ,n35[3] ,n110);
    nand g1357(n1894 ,n23[17] ,n1465);
    nand g1358(n3245 ,n24[25] ,n3219);
    nand g1359(n1819 ,n3466 ,n535);
    nand g1360(n1808 ,n22[31] ,n1464);
    dff g1361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1948), .Q(n31[25]));
    nand g1362(n963 ,n729 ,n745);
    nand g1363(n2076 ,n26[21] ,n1463);
    nand g1364(n1620 ,n8[30] ,n533);
    nand g1365(n1287 ,n6[10] ,n533);
    dff g1366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2410), .Q(n23[24]));
    dff g1367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2453), .Q(n28[11]));
    nand g1368(n2149 ,n1470 ,n1685);
    nor g1369(n612 ,n538 ,n28[28]);
    dff g1370(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2319), .Q(n30[23]));
    dff g1371(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2657), .Q(n34[1]));
    nand g1372(n1352 ,n29[23] ,n521);
    nor g1373(n1017 ,n894 ,n915);
    nand g1374(n2364 ,n2102 ,n1799);
    nand g1375(n1986 ,n30[24] ,n520);
    nand g1376(n2395 ,n1614 ,n1839);
    nand g1377(n1375 ,n3372 ,n1148);
    nand g1378(n1988 ,n30[21] ,n1463);
    nand g1379(n1005 ,n818 ,n778);
    nand g1380(n947 ,n628 ,n738);
    nand g1381(n771 ,n26[5] ,n538);
    xnor g1382(n3458 ,n316 ,n21[14]);
    nand g1383(n1865 ,n3520 ,n536);
    dff g1384(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2424), .Q(n28[1]));
    nand g1385(n1382 ,n32[18] ,n1149);
    nand g1386(n2144 ,n28[25] ,n1462);
    nand g1387(n1183 ,n27[23] ,n527);
    nand g1388(n2348 ,n2073 ,n1765);
    nand g1389(n2891 ,n1239 ,n2687);
    dff g1390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2013), .Q(n29[23]));
    dff g1391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2540), .Q(n21[15]));
    nand g1392(n1867 ,n3522 ,n536);
    dff g1393(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n843), .Q(n20[8]));
    nand g1394(n2349 ,n2076 ,n1766);
    not g1395(n387 ,n3401);
    nor g1396(n950 ,n538 ,n732);
    dff g1397(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2350), .Q(n26[20]));
    or g1398(n649 ,n549 ,n31[17]);
    nand g1399(n2758 ,n941 ,n2692);
    nand g1400(n2356 ,n2095 ,n1781);
    nor g1401(n474 ,n462 ,n467);
    nand g1402(n2352 ,n2207 ,n1768);
    nand g1403(n2522 ,n1873 ,n2307);
    nand g1404(n3169 ,n2812 ,n3061);
    nand g1405(n2136 ,n28[30] ,n1462);
    nand g1406(n2883 ,n1108 ,n2677);
    not g1407(n567 ,n27[13]);
    nand g1408(n717 ,n33[1] ,n1);
    dff g1409(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2493), .Q(n23[17]));
    nor g1410(n836 ,n591 ,n539);
    nand g1411(n1957 ,n1316 ,n1485);
    nand g1412(n2006 ,n30[2] ,n1463);
    nand g1413(n1956 ,n1315 ,n1258);
    nand g1414(n1536 ,n8[2] ,n530);
    nand g1415(n278 ,n22[24] ,n277);
    nand g1416(n1078 ,n935 ,n1033);
    xnor g1417(n3479 ,n276 ,n22[24]);
    xnor g1418(n3363 ,n6[18] ,n70);
    nand g1419(n3378 ,n3342 ,n3263);
    nand g1420(n1906 ,n23[5] ,n1465);
    nor g1421(n436 ,n372 ,n3417);
    nand g1422(n2711 ,n11[29] ,n2641);
    xnor g1423(n3482 ,n270 ,n22[21]);
    nand g1424(n3339 ,n3220 ,n22[4]);
    or g1425(n2574 ,n1552 ,n2246);
    nand g1426(n1622 ,n8[29] ,n533);
    nand g1427(n2881 ,n1139 ,n2675);
    nand g1428(n3434 ,n3344 ,n3278);
    nand g1429(n2013 ,n1352 ,n1298);
    nand g1430(n1427 ,n25[29] ,n521);
    nand g1431(n3239 ,n24[22] ,n3222);
    nand g1432(n1004 ,n822 ,n760);
    nand g1433(n226 ,n24[27] ,n225);
    nand g1434(n2916 ,n27[11] ,n2694);
    nand g1435(n1869 ,n3523 ,n537);
    xnor g1436(n3486 ,n265 ,n22[17]);
    not g1437(n1467 ,n1466);
    nand g1438(n3418 ,n3297 ,n3233);
    xnor g1439(n3550 ,n144 ,n23[15]);
    nor g1440(n2658 ,n2617 ,n2632);
    nand g1441(n250 ,n22[9] ,n249);
    nand g1442(n1508 ,n1133 ,n1123);
    nand g1443(n2419 ,n2205 ,n1747);
    nand g1444(n1178 ,n31[1] ,n527);
    nand g1445(n1863 ,n3518 ,n536);
    nand g1446(n3104 ,n2791 ,n2943);
    nand g1447(n2756 ,n943 ,n2692);
    nor g1448(n1030 ,n966 ,n978);
    nand g1449(n995 ,n820 ,n744);
    nand g1450(n1776 ,n3442 ,n535);
    nor g1451(n2965 ,n545 ,n2850);
    nand g1452(n3429 ,n3295 ,n3226);
    not g1453(n176 ,n175);
    nand g1454(n1112 ,n29[23] ,n1032);
    dff g1455(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3102), .Q(n10[16]));
    nand g1456(n2512 ,n1804 ,n2279);
    xnor g1457(n3540 ,n162 ,n23[25]);
    nand g1458(n1854 ,n3509 ,n537);
    nand g1459(n282 ,n22[26] ,n281);
    nand g1460(n2269 ,n21[13] ,n1951);
    nand g1461(n744 ,n26[7] ,n538);
    nor g1462(n1023 ,n972 ,n986);
    not g1463(n561 ,n6[13]);
    nand g1464(n3210 ,n2995 ,n3152);
    nand g1465(n2288 ,n24[26] ,n1950);
    nand g1466(n1197 ,n15 ,n1035);
    nand g1467(n1712 ,n6[18] ,n537);
    nand g1468(n981 ,n680 ,n807);
    dff g1469(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2661), .Q(n35[4]));
    nand g1470(n1658 ,n3560 ,n533);
    nand g1471(n1626 ,n8[26] ,n532);
    nand g1472(n3385 ,n3338 ,n3276);
    nand g1473(n1192 ,n25[20] ,n529);
    nand g1474(n1521 ,n8[14] ,n530);
    nand g1475(n1188 ,n1005 ,n1033);
    nand g1476(n1767 ,n8[20] ,n536);
    xnor g1477(n3448 ,n334 ,n21[24]);
    not g1478(n38 ,n6[28]);
    nand g1479(n3097 ,n2783 ,n2935);
    nand g1480(n1762 ,n8[25] ,n536);
    nand g1481(n856 ,n6[5] ,n37[0]);
    nand g1482(n2081 ,n1575 ,n1404);
    nand g1483(n1471 ,n29[21] ,n521);
    not g1484(n564 ,n6[15]);
    nor g1485(n3075 ,n2922 ,n3033);
    nand g1486(n1239 ,n25[8] ,n1032);
    dff g1487(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2439), .Q(n32[17]));
    nand g1488(n2042 ,n1368 ,n1478);
    nand g1489(n2905 ,n6[0] ,n2697);
    nand g1490(n1948 ,n1308 ,n1254);
    nand g1491(n1454 ,n25[8] ,n1147);
    xor g1492(n3360 ,n6[15] ,n64);
    nor g1493(n3063 ,n2745 ,n3021);
    nand g1494(n1484 ,n8[29] ,n531);
    nor g1495(n487 ,n460 ,n485);
    dff g1496(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2742), .Q(n34[0]));
    nand g1497(n846 ,n35[1] ,n1);
    nand g1498(n1730 ,n6[26] ,n534);
    nand g1499(n3181 ,n2988 ,n3053);
    dff g1500(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2398), .Q(n22[3]));
    nand g1501(n1980 ,n1339 ,n1273);
    not g1502(n2608 ,n2609);
    nor g1503(n2867 ,n992 ,n2691);
    nor g1504(n879 ,n662 ,n683);
    xnor g1505(n908 ,n6[29] ,n30[23]);
    dff g1506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2483), .Q(n23[7]));
    xnor g1507(n3563 ,n117 ,n23[2]);
    nand g1508(n1236 ,n27[13] ,n527);
    nor g1509(n1018 ,n911 ,n975);
    nand g1510(n986 ,n705 ,n774);
    dff g1511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2395), .Q(n22[6]));
    dff g1512(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2486), .Q(n23[10]));
    dff g1513(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2497), .Q(n21[1]));
    dff g1514(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2386), .Q(n22[14]));
    nand g1515(n1872 ,n3526 ,n537);
    nand g1516(n1706 ,n6[12] ,n536);
    dff g1517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2124), .Q(n25[19]));
    nand g1518(n2508 ,n1858 ,n2293);
    nand g1519(n1799 ,n8[8] ,n537);
    dff g1520(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1955), .Q(n27[29]));
    nand g1521(n2020 ,n1442 ,n1299);
    nand g1522(n2507 ,n1857 ,n2292);
    nand g1523(n1593 ,n3488 ,n531);
    nand g1524(n1704 ,n6[8] ,n537);
    nand g1525(n982 ,n659 ,n730);
    nand g1526(n3425 ,n3325 ,n3262);
    not g1527(n169 ,n168);
    nand g1528(n724 ,n29[17] ,n549);
    nand g1529(n2374 ,n1591 ,n1817);
    xnor g1530(n3465 ,n302 ,n21[7]);
    nor g1531(n3050 ,n2767 ,n3037);
    nand g1532(n1814 ,n22[26] ,n1464);
    not g1533(n2751 ,n2732);
    nand g1534(n1886 ,n23[25] ,n1465);
    nand g1535(n1487 ,n8[26] ,n531);
    not g1536(n584 ,n36[1]);
    nand g1537(n2045 ,n1353 ,n1369);
    nand g1538(n1940 ,n8[5] ,n535);
    nand g1539(n1450 ,n25[10] ,n1147);
    nand g1540(n1791 ,n8[10] ,n536);
    nand g1541(n2319 ,n2128 ,n1719);
    or g1542(n691 ,n555 ,n32[21]);
    dff g1543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3179), .Q(n11[1]));
    dff g1544(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2539), .Q(n21[14]));
    dff g1545(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2375), .Q(n22[22]));
    nand g1546(n212 ,n24[20] ,n211);
    nand g1547(n1861 ,n3516 ,n537);
    nand g1548(n445 ,n3408 ,n353);
    nand g1549(n1523 ,n8[6] ,n530);
    nand g1550(n2668 ,n7[26] ,n2642);
    dff g1551(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2363), .Q(n26[6]));
    nand g1552(n508 ,n395 ,n507);
    dff g1553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3174), .Q(n11[11]));
    nor g1554(n444 ,n377 ,n3397);
    not g1555(n532 ,n521);
    dff g1556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3186), .Q(n11[31]));
    xnor g1557(n3529 ,n182 ,n24[5]);
    or g1558(n2226 ,n1573 ,n2077);
    nand g1559(n2565 ,n1022 ,n2233);
    nand g1560(n3416 ,n3290 ,n3225);
    nand g1561(n3096 ,n2782 ,n2934);
    dff g1562(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2541), .Q(n21[16]));
    nand g1563(n1574 ,n1165 ,n1196);
    or g1564(n2228 ,n1578 ,n2082);
    nand g1565(n1335 ,n31[6] ,n522);
    nand g1566(n1633 ,n3540 ,n532);
    dff g1567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3113), .Q(n10[5]));
    dff g1568(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n797), .Q(n33[2]));
    nand g1569(n3331 ,n3221 ,n22[17]);
    nand g1570(n748 ,n31[15] ,n541);
    not g1571(n189 ,n188);
    nand g1572(n2200 ,n32[6] ,n1462);
    nand g1573(n2610 ,n1 ,n2597);
    nand g1574(n1417 ,n3351 ,n1148);
    nand g1575(n3330 ,n3221 ,n22[2]);
    nand g1576(n2394 ,n1613 ,n1838);
    dff g1577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2333), .Q(n30[3]));
    nand g1578(n340 ,n21[26] ,n339);
    nor g1579(n2239 ,n964 ,n1697);
    nand g1580(n3173 ,n2846 ,n3073);
    nand g1581(n184 ,n24[5] ,n183);
    nor g1582(n3567 ,n101 ,n103);
    nand g1583(n1272 ,n6[10] ,n531);
    nor g1584(n2970 ,n542 ,n2850);
    nand g1585(n447 ,n3420 ,n359);
    nand g1586(n2875 ,n1201 ,n2669);
    nor g1587(n1021 ,n973 ,n913);
    not g1588(n2216 ,n2086);
    buf g1589(n18[6], 1'b0);
    nand g1590(n1971 ,n1330 ,n1267);
    not g1591(n544 ,n6[11]);
    nand g1592(n2342 ,n2061 ,n1760);
    nand g1593(n1811 ,n22[29] ,n1464);
    nand g1594(n3302 ,n3220 ,n22[29]);
    nor g1595(n3062 ,n2814 ,n3019);
    nand g1596(n3043 ,n2857 ,n2770);
    or g1597(n1695 ,n21[0] ,n523);
    nand g1598(n2016 ,n1474 ,n1515);
    nand g1599(n2329 ,n2001 ,n1705);
    or g1600(n1696 ,n24[0] ,n520);
    nand g1601(n3174 ,n2915 ,n3077);
    xnor g1602(n3510 ,n218 ,n24[24]);
    dff g1603(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2346), .Q(n26[24]));
    nand g1604(n293 ,n21[17] ,n21[16]);
    nand g1605(n107 ,n35[1] ,n35[0]);
    nand g1606(n2560 ,n1696 ,n2314);
    not g1607(n551 ,n6[30]);
    dff g1608(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2389), .Q(n22[11]));
    nand g1609(n1365 ,n29[7] ,n521);
    not g1610(n1006 ,n1005);
    nand g1611(n2009 ,n30[0] ,n1463);
    nand g1612(n2151 ,n1459 ,n1681);
    nand g1613(n1685 ,n8[1] ,n533);
    nor g1614(n3057 ,n2572 ,n2970);
    nand g1615(n2145 ,n28[24] ,n1462);
    nand g1616(n2705 ,n2611 ,n2638);
    nand g1617(n1255 ,n6[29] ,n530);
    nand g1618(n2138 ,n1454 ,n1678);
    dff g1619(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3196), .Q(n11[3]));
    nand g1620(n466 ,n421 ,n428);
    nor g1621(n477 ,n466 ,n471);
    not g1622(n2631 ,n2620);
    nand g1623(n1270 ,n6[12] ,n531);
    nand g1624(n1278 ,n6[6] ,n532);
    nor g1625(n392 ,n358 ,n3399);
    nand g1626(n2859 ,n993 ,n2692);
    nand g1627(n2146 ,n1446 ,n1667);
    dff g1628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2458), .Q(n30[22]));
    nor g1629(n41 ,n6[6] ,n6[5]);
    nand g1630(n1407 ,n32[5] ,n1149);
    nand g1631(n1603 ,n3556 ,n532);
    nand g1632(n3275 ,n23[4] ,n3222);
    dff g1633(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1995), .Q(n27[16]));
    nand g1634(n3236 ,n23[21] ,n3219);
    nor g1635(n493 ,n417 ,n492);
    nand g1636(n3266 ,n24[29] ,n3222);
    dff g1637(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3118), .Q(n10[0]));
    nor g1638(n405 ,n387 ,n3433);
    nor g1639(n934 ,n617 ,n595);
    nor g1640(n677 ,n546 ,n31[16]);
    dff g1641(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2423), .Q(n32[6]));
    nand g1642(n300 ,n21[5] ,n299);
    nand g1643(n2091 ,n1589 ,n1417);
    nand g1644(n2436 ,n2188 ,n1735);
    not g1645(n576 ,n32[5]);
    nor g1646(n57 ,n46 ,n53);
    nand g1647(n2323 ,n2008 ,n1707);
    nand g1648(n1433 ,n25[19] ,n1147);
    or g1649(n883 ,n644 ,n641);
    nand g1650(n1103 ,n991 ,n1033);
    nand g1651(n2977 ,n6[12] ,n2849);
    nand g1652(n3045 ,n2862 ,n2771);
    nand g1653(n1715 ,n6[15] ,n537);
    or g1654(n1076 ,n931 ,n1034);
    nand g1655(n1240 ,n27[29] ,n1031);
    nor g1656(n1016 ,n6[5] ,n962);
    nand g1657(n1205 ,n25[31] ,n1032);
    nand g1658(n1855 ,n3510 ,n537);
    nand g1659(n3012 ,n9[0] ,n2848);
    dff g1660(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2487), .Q(n23[11]));
    dff g1661(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2577), .Q(n24[17]));
    nand g1662(n2555 ,n1776 ,n2252);
    not g1663(n115 ,n114);
    dff g1664(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3093), .Q(n10[25]));
    nor g1665(n2928 ,n1498 ,n2871);
    nand g1666(n1848 ,n8[0] ,n537);
    nand g1667(n3202 ,n3004 ,n3160);
    nand g1668(n2140 ,n28[28] ,n1462);
    not g1669(n364 ,n3416);
    nand g1670(n401 ,n3423 ,n354);
    nand g1671(n2433 ,n2190 ,n1941);
    nand g1672(n222 ,n24[25] ,n221);
    nand g1673(n3217 ,n2966 ,n3150);
    dff g1674(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2372), .Q(n22[25]));
    nand g1675(n1897 ,n23[14] ,n1465);
    nand g1676(n2819 ,n25[25] ,n2696);
    nor g1677(n430 ,n383 ,n3383);
    nand g1678(n2562 ,n926 ,n2415);
    nand g1679(n3381 ,n3329 ,n3269);
    nand g1680(n2474 ,n2139 ,n1914);
    dff g1681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2484), .Q(n23[8]));
    nand g1682(n334 ,n21[23] ,n333);
    nand g1683(n1599 ,n3478 ,n531);
    nand g1684(n1314 ,n31[21] ,n522);
    nor g1685(n837 ,n573 ,n539);
    buf g1686(n18[1], 1'b0);
    dff g1687(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2393), .Q(n26[2]));
    dff g1688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2475), .Q(n28[30]));
    nand g1689(n2824 ,n25[23] ,n2696);
    nand g1690(n1681 ,n8[5] ,n532);
    nand g1691(n1408 ,n3355 ,n1148);
    nand g1692(n1652 ,n8[19] ,n533);
    nand g1693(n3293 ,n3220 ,n22[8]);
    dff g1694(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2474), .Q(n28[29]));
    dff g1695(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2452), .Q(n28[10]));
    dff g1696(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2478), .Q(n23[2]));
    nand g1697(n3087 ,n2774 ,n2926);
    nand g1698(n801 ,n29[14] ,n559);
    dff g1699(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2530), .Q(n21[5]));
    nand g1700(n1485 ,n8[28] ,n531);
    nand g1701(n3419 ,n3301 ,n3237);
    nand g1702(n1432 ,n25[24] ,n1147);
    not g1703(n341 ,n340);
    nand g1704(n140 ,n23[12] ,n139);
    not g1705(n269 ,n268);
    not g1706(n61 ,n60);
    dff g1707(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n860), .Q(n20[5]));
    dff g1708(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2326), .Q(n30[13]));
    nand g1709(n3137 ,n1587 ,n2982);
    nand g1710(n3110 ,n2797 ,n2948);
    nand g1711(n2577 ,n1862 ,n2297);
    nand g1712(n1614 ,n3497 ,n530);
    nand g1713(n1391 ,n32[15] ,n1149);
    xnor g1714(n3453 ,n324 ,n21[19]);
    dff g1715(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2016), .Q(n27[8]));
    nand g1716(n2550 ,n1923 ,n2257);
    nand g1717(n1345 ,n27[2] ,n1146);
    not g1718(n317 ,n316);
    not g1719(n855 ,n854);
    nor g1720(n2831 ,n583 ,n2695);
    dff g1721(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2417), .Q(n32[1]));
    or g1722(n1063 ,n1057 ,n1056);
    nand g1723(n2473 ,n1998 ,n1703);
    nand g1724(n1507 ,n8[11] ,n530);
    nand g1725(n2470 ,n2143 ,n1917);
    nand g1726(n1526 ,n1168 ,n1079);
    xnor g1727(n903 ,n6[9] ,n30[3]);
    nand g1728(n3190 ,n2835 ,n3069);
    nand g1729(n2650 ,n2558 ,n2631);
    nor g1730(n494 ,n430 ,n493);
    nor g1731(n435 ,n356 ,n3402);
    nand g1732(n2455 ,n2166 ,n1932);
    dff g1733(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1954), .Q(n31[21]));
    nand g1734(n2446 ,n2179 ,n1938);
    nand g1735(n1387 ,n27[18] ,n1146);
    dff g1736(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2364), .Q(n26[8]));
    or g1737(n1051 ,n912 ,n906);
    nand g1738(n2310 ,n24[4] ,n1950);
    nand g1739(n2697 ,n1466 ,n2643);
    nor g1740(n68 ,n44 ,n66);
    not g1741(n382 ,n3433);
    nand g1742(n1847 ,n3503 ,n537);
    nand g1743(n500 ,n440 ,n499);
    nand g1744(n99 ,n34[3] ,n98);
    nand g1745(n3407 ,n3320 ,n3256);
    dff g1746(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3112), .Q(n10[6]));
    nor g1747(n3571 ,n96 ,n94);
    nand g1748(n1543 ,n30[7] ,n1150);
    nand g1749(n957 ,n742 ,n751);
    nand g1750(n1544 ,n3472 ,n530);
    not g1751(n577 ,n25[14]);
    nand g1752(n134 ,n23[9] ,n133);
    nor g1753(n3053 ,n2569 ,n2962);
    nand g1754(n1781 ,n8[13] ,n536);
    nand g1755(n2776 ,n10[29] ,n525);
    or g1756(n2572 ,n1563 ,n2248);
    nor g1757(n2653 ,n2603 ,n2624);
    nand g1758(n2046 ,n30[12] ,n1463);
    nand g1759(n1733 ,n6[23] ,n535);
    nand g1760(n2399 ,n2109 ,n1841);
    nand g1761(n2835 ,n1002 ,n2692);
    dff g1762(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2137), .Q(n25[9]));
    dff g1763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2368), .Q(n26[7]));
    nand g1764(n2923 ,n27[14] ,n2694);
    nand g1765(n202 ,n24[14] ,n201);
    not g1766(n133 ,n132);
    nand g1767(n3290 ,n3221 ,n22[7]);
    dff g1768(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2443), .Q(n32[20]));
    nand g1769(n3247 ,n24[20] ,n3219);
    dff g1770(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2413), .Q(n23[21]));
    nand g1771(n3195 ,n2851 ,n3080);
    nand g1772(n2739 ,n11[1] ,n2641);
    nor g1773(n637 ,n540 ,n32[0]);
    nand g1774(n274 ,n22[22] ,n273);
    dff g1775(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2337), .Q(n26[31]));
    nand g1776(n2727 ,n11[13] ,n2641);
    nand g1777(n348 ,n21[30] ,n347);
    nand g1778(n2078 ,n1436 ,n1403);
    nand g1779(n152 ,n23[19] ,n151);
    nand g1780(n1522 ,n1194 ,n1198);
    dff g1781(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2519), .Q(n24[10]));
    nand g1782(n3281 ,n24[26] ,n3219);
    xnor g1783(n3474 ,n286 ,n22[29]);
    nand g1784(n1785 ,n3450 ,n534);
    nor g1785(n84 ,n38 ,n83);
    not g1786(n385 ,n3378);
    not g1787(n245 ,n244);
    xnor g1788(n3493 ,n250 ,n22[10]);
    nand g1789(n2368 ,n2103 ,n1802);
    dff g1790(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2433), .Q(n28[4]));
    nand g1791(n1773 ,n8[14] ,n536);
    nand g1792(n1284 ,n6[14] ,n532);
    nand g1793(n2201 ,n28[1] ,n1462);
    nand g1794(n3122 ,n1555 ,n2992);
    nand g1795(n780 ,n30[13] ,n542);
    xnor g1796(n3373 ,n6[28] ,n83);
    nand g1797(n2337 ,n2051 ,n1756);
    nand g1798(n3197 ,n2868 ,n3083);
    dff g1799(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3208), .Q(n9[16]));
    nand g1800(n2494 ,n1641 ,n1893);
    nand g1801(n2438 ,n2186 ,n1940);
    nand g1802(n3231 ,n24[17] ,n3222);
    nand g1803(n3103 ,n2790 ,n2942);
    nor g1804(n481 ,n414 ,n476);
    nand g1805(n3305 ,n3221 ,n21[22]);
    nand g1806(n1070 ,n939 ,n1033);
    nand g1807(n1224 ,n29[12] ,n529);
    nand g1808(n2039 ,n1435 ,n1287);
    nand g1809(n1629 ,n3536 ,n532);
    nand g1810(n1520 ,n1212 ,n1172);
    dff g1811(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2392), .Q(n22[8]));
    nand g1812(n3033 ,n2726 ,n2923);
    not g1813(n541 ,n6[21]);
    nor g1814(n634 ,n559 ,n29[14]);
    nand g1815(n2142 ,n28[27] ,n1462);
    nand g1816(n2448 ,n2176 ,n1937);
    dff g1817(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2172), .Q(n90));
    nand g1818(n1553 ,n30[18] ,n1150);
    nand g1819(n710 ,n29[6] ,n562);
    nand g1820(n2241 ,n1250 ,n1911);
    not g1821(n225 ,n224);
    nand g1822(n2505 ,n1855 ,n2290);
    nand g1823(n790 ,n32[11] ,n554);
    nand g1824(n2387 ,n1592 ,n1829);
    dff g1825(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3185), .Q(n9[19]));
    nand g1826(n2304 ,n24[10] ,n1950);
    not g1827(n555 ,n6[27]);
    nand g1828(n2762 ,n936 ,n2692);
    dff g1829(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2114), .Q(n25[28]));
    nand g1830(n56 ,n6[15] ,n52);
    nand g1831(n803 ,n30[1] ,n563);
    nand g1832(n2351 ,n2003 ,n1714);
    nand g1833(n1325 ,n31[13] ,n522);
    dff g1834(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2400), .Q(n22[2]));
    nand g1835(n785 ,n13 ,n1);
    nand g1836(n2463 ,n2154 ,n1925);
    nand g1837(n1308 ,n31[25] ,n522);
    dff g1838(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2039), .Q(n29[4]));
    dff g1839(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2134), .Q(n25[10]));
    dff g1840(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3170), .Q(n11[26]));
    dff g1841(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2171), .Q(n92));
    dff g1842(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1693), .Q(n31[23]));
    nor g1843(n642 ,n545 ,n32[18]);
    nand g1844(n1707 ,n6[7] ,n536);
    nand g1845(n1656 ,n3559 ,n533);
    dff g1846(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3110), .Q(n10[8]));
    dff g1847(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1973), .Q(n31[8]));
    nand g1848(n2398 ,n1551 ,n1843);
    or g1849(n716 ,n33[0] ,n33[1]);
    nand g1850(n2347 ,n2071 ,n1764);
    nand g1851(n1334 ,n31[7] ,n1146);
    nand g1852(n975 ,n632 ,n815);
    nand g1853(n1954 ,n1314 ,n1257);
    nor g1854(n2612 ,n3574 ,n2598);
    nand g1855(n1190 ,n27[9] ,n527);
    xnor g1856(n3462 ,n308 ,n21[10]);
    xnor g1857(n861 ,n545 ,n29[18]);
    nand g1858(n1974 ,n1334 ,n1269);
    nand g1859(n2520 ,n1871 ,n2305);
    nand g1860(n1069 ,n936 ,n1033);
    dff g1861(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3172), .Q(n11[18]));
    nor g1862(n685 ,n549 ,n32[17]);
    dff g1863(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2011), .Q(n27[9]));
    nand g1864(n166 ,n23[26] ,n165);
    not g1865(n253 ,n252);
    nand g1866(n2161 ,n28[16] ,n1462);
    not g1867(n263 ,n262);
    nand g1868(n2052 ,n1374 ,n1545);
    nand g1869(n424 ,n3393 ,n381);
    not g1870(n550 ,n6[28]);
    or g1871(n469 ,n460 ,n457);
    xnor g1872(n3492 ,n252 ,n22[11]);
    nand g1873(n1435 ,n29[4] ,n521);
    or g1874(n1697 ,n963 ,n1252);
    buf g1875(n19[2], 1'b0);
    nand g1876(n1326 ,n27[25] ,n1146);
    nand g1877(n2994 ,n9[21] ,n2848);
    nand g1878(n2101 ,n26[9] ,n520);
    nand g1879(n1119 ,n29[9] ,n1032);
    nand g1880(n2889 ,n1221 ,n2684);
    dff g1881(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3099), .Q(n10[19]));
    or g1882(n940 ,n613 ,n593);
    nor g1883(n655 ,n552 ,n30[4]);
    nand g1884(n2618 ,n34[0] ,n2599);
    nand g1885(n499 ,n439 ,n498);
    not g1886(n536 ,n520);
    nand g1887(n972 ,n687 ,n787);
    nor g1888(n610 ,n538 ,n28[29]);
    or g1889(n877 ,n653 ,n652);
    or g1890(n2222 ,n1565 ,n2068);
    dff g1891(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2025), .Q(n29[14]));
    nor g1892(n2959 ,n551 ,n2850);
    nand g1893(n1642 ,n8[23] ,n532);
    nand g1894(n3270 ,n23[17] ,n3222);
    nand g1895(n2537 ,n1796 ,n2270);
    or g1896(n1463 ,n6[5] ,n1152);
    nand g1897(n3001 ,n9[14] ,n2848);
    nand g1898(n834 ,n37[0] ,n538);
    dff g1899(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3096), .Q(n10[23]));
    nor g1900(n839 ,n589 ,n539);
    nand g1901(n3015 ,n9[1] ,n2848);
    nand g1902(n1740 ,n6[16] ,n535);
    nor g1903(n2814 ,n571 ,n2695);
    not g1904(n2645 ,n2634);
    nand g1905(n711 ,n31[3] ,n560);
    nand g1906(n2882 ,n1222 ,n2676);
    nand g1907(n2033 ,n1366 ,n1532);
    nand g1908(n491 ,n422 ,n490);
    nand g1909(n2157 ,n1350 ,n1682);
    nand g1910(n149 ,n23[16] ,n147);
    nand g1911(n1995 ,n1377 ,n1689);
    nand g1912(n3309 ,n3220 ,n22[12]);
    nand g1913(n1182 ,n31[0] ,n527);
    nand g1914(n989 ,n672 ,n726);
    dff g1915(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2155), .Q(n27[10]));
    or g1916(n2587 ,n1050 ,n2580);
    nand g1917(n2841 ,n27[18] ,n2694);
    not g1918(n301 ,n300);
    dff g1919(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1953), .Q(n31[22]));
    dff g1920(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2491), .Q(n23[15]));
    nand g1921(n3027 ,n2720 ,n2833);
    nand g1922(n2511 ,n1861 ,n2296);
    nand g1923(n1145 ,n29[5] ,n1032);
    nand g1924(n705 ,n30[24] ,n551);
    not g1925(n585 ,n36[2]);
    xnor g1926(n3536 ,n170 ,n23[29]);
    nand g1927(n48 ,n6[14] ,n6[13]);
    nand g1928(n921 ,n661 ,n783);
    nand g1929(n2818 ,n27[26] ,n2694);
    nand g1930(n3251 ,n23[14] ,n3222);
    or g1931(n681 ,n543 ,n31[12]);
    nand g1932(n1503 ,n1158 ,n1160);
    dff g1933(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3145), .Q(n11[28]));
    nand g1934(n2109 ,n26[1] ,n520);
    nand g1935(n2397 ,n1615 ,n1842);
    not g1936(n553 ,n6[29]);
    nor g1937(n594 ,n26[13] ,n6[5]);
    nand g1938(n1930 ,n8[15] ,n534);
    nand g1939(n1135 ,n29[22] ,n1032);
    nand g1940(n1528 ,n1126 ,n1117);
    dff g1941(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2121), .Q(n25[22]));
    nor g1942(n893 ,n695 ,n697);
    nand g1943(n1385 ,n32[17] ,n1149);
    nor g1944(n618 ,n538 ,n28[13]);
    nand g1945(n3311 ,n3221 ,n22[22]);
    nand g1946(n2461 ,n2158 ,n1927);
    nand g1947(n802 ,n29[16] ,n546);
    dff g1948(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3183), .Q(n9[25]));
    not g1949(n139 ,n138);
    not g1950(n2849 ,n2850);
    nand g1951(n1120 ,n27[2] ,n1031);
    dff g1952(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2526), .Q(n24[3]));
    nand g1953(n2380 ,n1605 ,n1824);
    nand g1954(n44 ,n6[18] ,n6[17]);
    dff g1955(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3197), .Q(n11[0]));
    nand g1956(n3272 ,n23[3] ,n3222);
    nand g1957(n154 ,n23[20] ,n153);
    nand g1958(n1899 ,n23[12] ,n1465);
    nand g1959(n2870 ,n1210 ,n2682);
    dff g1960(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2366), .Q(n22[30]));
    nand g1961(n1900 ,n23[11] ,n1465);
    nand g1962(n3237 ,n23[10] ,n3222);
    xnor g1963(n886 ,n6[30] ,n29[24]);
    nand g1964(n1947 ,n1481 ,n1580);
    or g1965(n647 ,n563 ,n31[1]);
    nand g1966(n2544 ,n1788 ,n2263);
    nand g1967(n1111 ,n29[15] ,n1032);
    not g1968(n249 ,n248);
    nand g1969(n1676 ,n30[20] ,n1150);
    nand g1970(n1313 ,n27[29] ,n1146);
    xnor g1971(n923 ,n6[16] ,n30[10]);
    dff g1972(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2344), .Q(n30[12]));
    nand g1973(n2148 ,n28[23] ,n523);
    buf g1974(n19[0], 1'b0);
    nand g1975(n1923 ,n3447 ,n535);
    nor g1976(n1092 ,n1046 ,n1011);
    nand g1977(n246 ,n22[7] ,n245);
    dff g1978(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2084), .Q(n31[0]));
    nand g1979(n1077 ,n934 ,n1033);
    not g1980(n459 ,n458);
    not g1981(n3219 ,n3221);
    nand g1982(n216 ,n24[22] ,n215);
    not g1983(n360 ,n3430);
    nand g1984(n1413 ,n3352 ,n1148);
    nand g1985(n1953 ,n1312 ,n1256);
    nand g1986(n1189 ,n29[1] ,n1032);
    nor g1987(n463 ,n435 ,n429);
    nand g1988(n2896 ,n1067 ,n2700);
    buf g1989(n18[0], 1'b0);
    nand g1990(n1689 ,n8[16] ,n531);
    dff g1991(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2383), .Q(n22[16]));
    nand g1992(n3192 ,n2924 ,n3074);
    or g1993(n632 ,n560 ,n32[3]);
    nand g1994(n1641 ,n3547 ,n532);
    xnor g1995(n3359 ,n6[14] ,n67);
    nand g1996(n3011 ,n9[4] ,n2848);
    nand g1997(n2679 ,n7[15] ,n2642);
    nand g1998(n1864 ,n3519 ,n537);
    nand g1999(n1438 ,n25[17] ,n1147);
    dff g2000(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2369), .Q(n22[28]));
    nand g2001(n2738 ,n11[2] ,n2641);
    nand g2002(n1530 ,n8[4] ,n530);
    xnor g2003(n890 ,n6[20] ,n31[14]);
    nand g2004(n1551 ,n3500 ,n530);
    nand g2005(n1288 ,n6[8] ,n532);
    nor g2006(n2660 ,n2612 ,n2644);
    dff g2007(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2152), .Q(n25[0]));
    nand g2008(n2343 ,n2066 ,n1761);
    or g2009(n2591 ,n2588 ,n2584);
    not g2010(n321 ,n320);
    nand g2011(n1837 ,n22[8] ,n1464);
    nand g2012(n3327 ,n3220 ,n22[24]);
    nand g2013(n1942 ,n8[3] ,n534);
    nand g2014(n2420 ,n2204 ,n1746);
    nand g2015(n3321 ,n3221 ,n22[15]);
    nor g2016(n77 ,n55 ,n74);
    nand g2017(n1068 ,n927 ,n1033);
    not g2018(n543 ,n6[18]);
    nand g2019(n1598 ,n3477 ,n531);
    xnor g2020(n3507 ,n224 ,n24[27]);
    nor g2021(n619 ,n538 ,n28[12]);
    nand g2022(n1545 ,n30[22] ,n1150);
    nand g2023(n1085 ,n1054 ,n1017);
    not g2024(n537 ,n1463);
    nor g2025(n406 ,n386 ,n3385);
    nand g2026(n451 ,n3436 ,n371);
    nand g2027(n468 ,n416 ,n411);
    dff g2028(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2450), .Q(n32[25]));
    dff g2029(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n829), .Q(n19[6]));
    nand g2030(n2074 ,n1568 ,n1399);
    not g2031(n347 ,n346);
    nand g2032(n3093 ,n2780 ,n2932);
    nand g2033(n2272 ,n21[10] ,n1951);
    nand g2034(n2134 ,n1450 ,n1674);
    nand g2035(n177 ,n24[17] ,n24[16]);
    nand g2036(n411 ,n3402 ,n356);
    nand g2037(n2873 ,n1207 ,n2667);
    nand g2038(n1878 ,n3532 ,n537);
    dff g2039(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3143), .Q(n9[2]));
    nand g2040(n2335 ,n2009 ,n1708);
    nand g2041(n2826 ,n27[23] ,n2694);
    nand g2042(n2464 ,n2153 ,n1924);
    nand g2043(n421 ,n3428 ,n365);
    nand g2044(n1339 ,n31[3] ,n1146);
    not g2045(n359 ,n3388);
    nand g2046(n1651 ,n3555 ,n533);
    nand g2047(n2025 ,n1379 ,n1290);
    nand g2048(n288 ,n22[29] ,n287);
    nand g2049(n2709 ,n11[31] ,n2641);
    nand g2050(n769 ,n26[9] ,n538);
    not g2051(n547 ,n6[16]);
    nand g2052(n1478 ,n3376 ,n1148);
    nand g2053(n707 ,n26[3] ,n538);
    nand g2054(n1455 ,n3371 ,n1148);
    nor g2055(n797 ,n585 ,n539);
    nand g2056(n83 ,n6[27] ,n80);
    nor g2057(n621 ,n538 ,n28[8]);
    nand g2058(n2625 ,n854 ,n2610);
    nand g2059(n2001 ,n30[8] ,n520);
    nand g2060(n124 ,n23[4] ,n123);
    nand g2061(n1844 ,n22[2] ,n1464);
    nand g2062(n1743 ,n6[13] ,n535);
    nand g2063(n3223 ,n23[26] ,n3222);
    dff g2064(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2167), .Q(n25[2]));
    nand g2065(n1987 ,n30[22] ,n1463);
    nand g2066(n2557 ,n36[0] ,n2416);
    nand g2067(n1064 ,n629 ,n1053);
    nand g2068(n2456 ,n2165 ,n1931);
    nand g2069(n2408 ,n1632 ,n1885);
    nor g2070(n1045 ,n877 ,n985);
    nand g2071(n434 ,n3384 ,n364);
    not g2072(n2754 ,n2738);
    nand g2073(n1495 ,n1205 ,n1072);
    nand g2074(n1612 ,n3495 ,n530);
    nand g2075(n2267 ,n21[15] ,n1951);
    nand g2076(n1392 ,n3365 ,n1148);
    dff g2077(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3105), .Q(n10[9]));
    nand g2078(n1412 ,n3353 ,n1148);
    nand g2079(n2407 ,n1631 ,n1884);
    dff g2080(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1997), .Q(n27[12]));
    not g2081(n992 ,n991);
    nand g2082(n1914 ,n8[29] ,n535);
    not g2083(n185 ,n184);
    nor g2084(n2662 ,n2614 ,n2646);
    nand g2085(n1199 ,n14 ,n1035);
    nand g2086(n2984 ,n9[31] ,n2848);
    nand g2087(n1989 ,n30[19] ,n520);
    nand g2088(n961 ,n743 ,n776);
    nand g2089(n3259 ,n24[31] ,n3222);
    or g2090(n1245 ,n1042 ,n1097);
    nor g2091(n925 ,n828 ,n720);
    dff g2092(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2146), .Q(n27[19]));
    nand g2093(n1728 ,n6[28] ,n534);
    nand g2094(n3123 ,n1388 ,n2967);
    nand g2095(n2082 ,n1407 ,n1406);
    dff g2096(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1821), .Q(n31[24]));
    nand g2097(n1784 ,n8[11] ,n536);
    nand g2098(n214 ,n24[21] ,n213);
    nand g2099(n3121 ,n1473 ,n2961);
    nand g2100(n1519 ,n1209 ,n1211);
    nand g2101(n3308 ,n3220 ,n21[24]);
    nand g2102(n1571 ,n1162 ,n1119);
    nor g2103(n2603 ,n3567 ,n2600);
    nor g2104(n643 ,n557 ,n29[20]);
    nand g2105(n2095 ,n26[13] ,n520);
    dff g2106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1965), .Q(n31[13]));
    dff g2107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2407), .Q(n23[27]));
    dff g2108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3175), .Q(n11[8]));
    nand g2109(n2515 ,n1865 ,n2300);
    nand g2110(n1337 ,n31[4] ,n1146);
    nand g2111(n2504 ,n1854 ,n2289);
    nor g2112(n2626 ,n837 ,n2608);
    not g2113(n2695 ,n2696);
    nand g2114(n1206 ,n27[15] ,n1031);
    dff g2115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2021), .Q(n27[17]));
    not g2116(n141 ,n140);
    nand g2117(n2784 ,n10[21] ,n525);
    nand g2118(n2636 ,n850 ,n2610);
    not g2119(n108 ,n107);
    dff g2120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2438), .Q(n28[5]));
    nand g2121(n1737 ,n6[19] ,n535);
    nand g2122(n3141 ,n2901 ,n3011);
    dff g2123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3214), .Q(n9[31]));
    nand g2124(n122 ,n23[3] ,n121);
    nand g2125(n1617 ,n3502 ,n530);
    nand g2126(n1748 ,n6[8] ,n535);
    nand g2127(n2023 ,n1357 ,n1292);
    nand g2128(n2377 ,n1601 ,n1820);
    nand g2129(n3386 ,n3340 ,n3277);
    dff g2130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2460), .Q(n28[17]));
    nor g2131(n3151 ,n2219 ,n3123);
    nand g2132(n2382 ,n2106 ,n1822);
    not g2133(n556 ,n6[25]);
    nand g2134(n45 ,n6[22] ,n6[21]);
    nand g2135(n3256 ,n24[30] ,n3222);
    nand g2136(n1323 ,n27[26] ,n522);
    nand g2137(n2189 ,n32[14] ,n1462);
    xnor g2138(n3470 ,n291 ,n21[2]);
    nand g2139(n1100 ,n766 ,n1023);
    nand g2140(n1702 ,n6[21] ,n536);
    nand g2141(n395 ,n3391 ,n351);
    nand g2142(n298 ,n21[4] ,n297);
    nand g2143(n2103 ,n26[7] ,n520);
    nand g2144(n3250 ,n24[27] ,n3222);
    dff g2145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2425), .Q(n32[7]));
    nand g2146(n2714 ,n11[26] ,n2641);
    nand g2147(n2437 ,n2187 ,n1734);
    nand g2148(n1664 ,n8[18] ,n532);
    nand g2149(n1797 ,n3461 ,n534);
    nand g2150(n1903 ,n23[8] ,n1465);
    nand g2151(n2204 ,n32[4] ,n1462);
    or g2152(n3165 ,n2960 ,n3120);
    nand g2153(n1824 ,n22[18] ,n1464);
    nand g2154(n1636 ,n3543 ,n532);
    nand g2155(n1542 ,n30[23] ,n1150);
    nand g2156(n2273 ,n21[9] ,n1951);
    nand g2157(n1970 ,n1329 ,n1266);
    xor g2158(n864 ,n6[28] ,n32[22]);
    nor g2159(n2614 ,n3576 ,n2598);
    nand g2160(n1445 ,n25[12] ,n521);
    nand g2161(n1474 ,n27[8] ,n522);
    nand g2162(n3004 ,n9[11] ,n2848);
    nand g2163(n1380 ,n3370 ,n1148);
    dff g2164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3147), .Q(n11[14]));
    nand g2165(n1918 ,n8[25] ,n535);
    nor g2166(n603 ,n26[6] ,n6[5]);
    xor g2167(n901 ,n6[17] ,n30[11]);
    nand g2168(n464 ,n426 ,n423);
    not g2169(n358 ,n3431);
    nand g2170(n3420 ,n3306 ,n3240);
    dff g2171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3188), .Q(n11[22]));
    nand g2172(n1457 ,n27[1] ,n1146);
    nor g2173(n2605 ,n3569 ,n2600);
    nand g2174(n1735 ,n6[21] ,n535);
    nor g2175(n3071 ,n2748 ,n3029);
    nand g2176(n3019 ,n2712 ,n2813);
    xnor g2177(n3548 ,n149 ,n23[17]);
    nand g2178(n1114 ,n25[1] ,n1032);
    xnor g2179(n3512 ,n214 ,n24[22]);
    dff g2180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2503), .Q(n24[26]));
    nand g2181(n1115 ,n25[18] ,n529);
    dff g2182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3141), .Q(n9[4]));
    nand g2183(n816 ,n28[0] ,n6[5]);
    nand g2184(n3413 ,n3339 ,n3275);
    nor g2185(n3070 ,n2838 ,n3028);
    nand g2186(n825 ,n90 ,n1);
    nand g2187(n1329 ,n31[10] ,n522);
    not g2188(n277 ,n276);
    nand g2189(n3315 ,n3220 ,n21[27]);
    nand g2190(n1619 ,n1177 ,n1122);
    nor g2191(n2848 ,n925 ,n2697);
    nand g2192(n2375 ,n1624 ,n1818);
    nor g2193(n2623 ,n840 ,n2608);
    nand g2194(n2089 ,n26[17] ,n520);
    dff g2195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2322), .Q(n30[17]));
    nand g2196(n1907 ,n23[4] ,n1465);
    nand g2197(n3232 ,n24[18] ,n3219);
    nand g2198(n1606 ,n3486 ,n530);
    nand g2199(n807 ,n32[18] ,n545);
    nor g2200(n1150 ,n6[5] ,n1034);
    xnor g2201(n3553 ,n138 ,n23[12]);
    dff g2202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2545), .Q(n21[20]));
    nand g2203(n2158 ,n28[18] ,n1462);
    nand g2204(n425 ,n3392 ,n374);
    nand g2205(n1958 ,n1317 ,n1259);
    nand g2206(n1355 ,n27[6] ,n522);
    nand g2207(n1406 ,n3356 ,n1148);
    not g2208(n197 ,n196);
    or g2209(n400 ,n371 ,n3436);
    nor g2210(n732 ,n575 ,n6[6]);
    nor g2211(n407 ,n367 ,n3409);
    nand g2212(n2027 ,n1359 ,n1530);
    nand g2213(n1451 ,n25[9] ,n521);
    nand g2214(n3288 ,n3220 ,n22[19]);
    nand g2215(n323 ,n21[16] ,n321);
    nand g2216(n338 ,n21[25] ,n337);
    dff g2217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1983), .Q(n31[1]));
    nand g2218(n1832 ,n22[11] ,n1464);
    nand g2219(n2516 ,n1869 ,n2303);
    not g2220(n586 ,n34[6]);
    nand g2221(n1418 ,n29[22] ,n1147);
    nand g2222(n2345 ,n2063 ,n1762);
    nand g2223(n2195 ,n28[3] ,n1462);
    dff g2224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2489), .Q(n23[13]));
    nand g2225(n1462 ,n6[5] ,n1151);
    nand g2226(n2868 ,n25[0] ,n2696);
    xnor g2227(n3517 ,n207 ,n24[17]);
    nand g2228(n1166 ,n27[6] ,n1031);
    xnor g2229(n3514 ,n210 ,n24[20]);
    nand g2230(n953 ,n704 ,n793);
    nand g2231(n2024 ,n1355 ,n1523);
    nor g2232(n1038 ,n875 ,n948);
    xnor g2233(n902 ,n6[24] ,n30[18]);
    not g2234(n201 ,n200);
    or g2235(n1752 ,n990 ,n1245);
    nand g2236(n1646 ,n3551 ,n532);
    nand g2237(n1925 ,n8[20] ,n535);
    nand g2238(n1673 ,n8[11] ,n532);
    dff g2239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2020), .Q(n29[18]));
    not g2240(n583 ,n25[21]);
    nand g2241(n2107 ,n26[3] ,n1463);
    dff g2242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2554), .Q(n21[27]));
    not g2243(n93 ,n34[4]);
    nand g2244(n1050 ,n888 ,n890);
    nand g2245(n3267 ,n24[3] ,n3219);
    nor g2246(n3157 ,n2225 ,n3129);
    xnor g2247(n3353 ,n6[8] ,n49);
    nand g2248(n3039 ,n2909 ,n2768);
    nand g2249(n1126 ,n25[7] ,n529);
    nand g2250(n2162 ,n1468 ,n1683);
    xnor g2251(n3478 ,n278 ,n22[25]);
    nand g2252(n1675 ,n8[9] ,n533);
    nand g2253(n2193 ,n28[2] ,n523);
    nand g2254(n2405 ,n1629 ,n1882);
    nand g2255(n2392 ,n1612 ,n1837);
    nand g2256(n2073 ,n26[22] ,n1463);
    or g2257(n680 ,n546 ,n32[16]);
    nand g2258(n2480 ,n1659 ,n1907);
    nand g2259(n1490 ,n8[23] ,n531);
    dff g2260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2044), .Q(n29[2]));
    nand g2261(n2026 ,n30[4] ,n520);
    nor g2262(n76 ,n45 ,n74);
    xor g2263(n3471 ,n21[1] ,n21[0]);
    dff g2264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2556), .Q(n21[31]));
    xnor g2265(n3554 ,n136 ,n23[11]);
    nand g2266(n1025 ,n951 ,n867);
    nor g2267(n322 ,n293 ,n320);
    nor g2268(n697 ,n541 ,n31[15]);
    nor g2269(n599 ,n26[28] ,n6[5]);
    nor g2270(n2950 ,n1528 ,n2893);
    not g2271(n370 ,n3390);
    nand g2272(n1046 ,n880 ,n879);
    nand g2273(n3399 ,n3305 ,n3239);
    nand g2274(n2728 ,n11[12] ,n2641);
    or g2275(n675 ,n561 ,n30[7]);
    dff g2276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2509), .Q(n24[20]));
    nand g2277(n1366 ,n27[3] ,n522);
    nand g2278(n2259 ,n21[23] ,n1951);
    nor g2279(n930 ,n621 ,n605);
    nand g2280(n1560 ,n30[14] ,n1150);
    nand g2281(n2525 ,n1876 ,n2310);
    nand g2282(n418 ,n3380 ,n379);
    xor g2283(n906 ,n6[18] ,n32[12]);
    not g2284(n860 ,n859);
    nand g2285(n2112 ,n1426 ,n1620);
    dff g2286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2479), .Q(n23[3]));
    nand g2287(n2510 ,n1860 ,n2295);
    not g2288(n155 ,n154);
    nand g2289(n2130 ,n1443 ,n1670);
    nand g2290(n67 ,n6[13] ,n63);
    not g2291(n1152 ,n1151);
    nor g2292(n2960 ,n553 ,n2850);
    nand g2293(n3343 ,n3220 ,n21[10]);
    nand g2294(n3227 ,n24[15] ,n3222);
    not g2295(n143 ,n142);
    nand g2296(n3176 ,n2856 ,n3081);
    dff g2297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2328), .Q(n30[9]));
    nand g2298(n2804 ,n10[1] ,n2690);
    nor g2299(n645 ,n541 ,n29[15]);
    not g2300(n376 ,n3397);
    nand g2301(n2823 ,n25[24] ,n2696);
    nand g2302(n1342 ,n31[1] ,n522);
    nor g2303(n3154 ,n2222 ,n3126);
    nand g2304(n2810 ,n27[30] ,n2694);
    dff g2305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3106), .Q(n10[13]));
    dff g2306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2332), .Q(n30[4]));
    dff g2307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1961), .Q(n31[16]));
    nand g2308(n302 ,n21[6] ,n301);
    nand g2309(n1395 ,n3363 ,n1148);
    xnor g2310(n3568 ,n34[4] ,n99);
    dff g2311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2377), .Q(n22[21]));
    nand g2312(n1648 ,n3553 ,n532);
    nand g2313(n2476 ,n2135 ,n1912);
    nand g2314(n730 ,n29[8] ,n558);
    not g2315(n591 ,n34[2]);
    dff g2316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2335), .Q(n30[0]));
    dff g2317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2405), .Q(n23[29]));
    nand g2318(n3140 ,n2905 ,n3012);
    nand g2319(n503 ,n447 ,n502);
    xnor g2320(n3509 ,n220 ,n24[25]);
    nand g2321(n1172 ,n25[30] ,n529);
    nand g2322(n3178 ,n2864 ,n3086);
    nand g2323(n1434 ,n25[20] ,n521);
    nand g2324(n457 ,n402 ,n400);
    nor g2325(n3156 ,n2224 ,n3128);
    nand g2326(n1088 ,n1049 ,n1038);
    nand g2327(n913 ,n693 ,n706);
    nand g2328(n3316 ,n3220 ,n21[28]);
    nand g2329(n230 ,n24[29] ,n229);
    nand g2330(n2579 ,n1062 ,n2559);
    nand g2331(n2465 ,n2150 ,n1922);
    nand g2332(n2275 ,n21[7] ,n1951);
    or g2333(n2583 ,n1052 ,n2567);
    nand g2334(n1999 ,n1365 ,n1277);
    nand g2335(n1215 ,n25[16] ,n529);
    or g2336(n416 ,n366 ,n3435);
    nand g2337(n2495 ,n1640 ,n1892);
    xnor g2338(n3468 ,n296 ,n21[4]);
    dff g2339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2133), .Q(n25[11]));
    nand g2340(n1422 ,n25[21] ,n521);
    dff g2341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2029), .Q(n29[12]));
    nand g2342(n1138 ,n27[5] ,n1031);
    nand g2343(n2493 ,n1643 ,n1894);
    not g2344(n2211 ,n2055);
    nand g2345(n1943 ,n8[2] ,n535);
    nand g2346(n2528 ,n1879 ,n2313);
    nor g2347(n1037 ,n883 ,n909);
    dff g2348(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2434), .Q(n32[13]));
    nand g2349(n1443 ,n25[14] ,n1147);
    nand g2350(n1276 ,n6[12] ,n532);
    nand g2351(n2886 ,n1077 ,n2680);
    nand g2352(n2292 ,n24[22] ,n1950);
    nand g2353(n233 ,n22[1] ,n22[0]);
    nand g2354(n2080 ,n26[20] ,n1463);
    nand g2355(n3029 ,n2840 ,n2837);
    not g2356(n368 ,n3421);
    nand g2357(n1419 ,n27[10] ,n522);
    nand g2358(n2678 ,n7[16] ,n2642);
    not g2359(n379 ,n3412);
    nand g2360(n2541 ,n1792 ,n2266);
    nand g2361(n1472 ,n25[0] ,n521);
    nand g2362(n1097 ,n900 ,n1016);
    nand g2363(n2876 ,n1170 ,n2670);
    nand g2364(n3284 ,n24[12] ,n3219);
    or g2365(n2217 ,n1546 ,n2052);
    nand g2366(n978 ,n649 ,n711);
    dff g2367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1960), .Q(n31[17]));
    not g2368(n545 ,n6[24]);
    nor g2369(n615 ,n538 ,n28[17]);
    nand g2370(n1298 ,n6[29] ,n533);
    nand g2371(n2485 ,n1603 ,n1902);
    nand g2372(n3024 ,n2717 ,n2824);
    nand g2373(n2059 ,n26[28] ,n520);
    nor g2374(n2236 ,n989 ,n1752);
    nand g2375(n706 ,n32[3] ,n560);
    nand g2376(n3391 ,n3289 ,n3224);
    nand g2377(n974 ,n688 ,n827);
    nor g2378(n3054 ,n2575 ,n2963);
    nand g2379(n3092 ,n2779 ,n2931);
    nor g2380(n2956 ,n1537 ,n2899);
    dff g2381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2482), .Q(n23[6]));
    or g2382(n1066 ,n929 ,n1034);
    nand g2383(n3023 ,n2821 ,n2822);
    or g2384(n2576 ,n1508 ,n2242);
    nand g2385(n1766 ,n8[21] ,n536);
    nand g2386(n2501 ,n1850 ,n2285);
    nand g2387(n1718 ,n6[28] ,n537);
    nand g2388(n2246 ,n1550 ,n2212);
    nand g2389(n850 ,n35[2] ,n1);
    not g2390(n161 ,n160);
    nand g2391(n1756 ,n8[31] ,n536);
    nand g2392(n800 ,n32[14] ,n559);
    dff g2393(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2403), .Q(n23[31]));
    xnor g2394(n3475 ,n284 ,n22[28]);
    nand g2395(n848 ,n35[3] ,n1);
    nand g2396(n2913 ,n25[9] ,n2696);
    nand g2397(n2811 ,n27[29] ,n2694);
    nand g2398(n3292 ,n3221 ,n21[16]);
    xnor g2399(n3565 ,n34[7] ,n104);
    nand g2400(n314 ,n21[12] ,n313);
    nand g2401(n738 ,n30[21] ,n555);
    nand g2402(n1901 ,n23[10] ,n1465);
    not g2403(n540 ,n6[6]);
    nand g2404(n820 ,n28[7] ,n6[5]);
    nand g2405(n486 ,n452 ,n483);
    dff g2406(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2436), .Q(n32[15]));
    nor g2407(n626 ,n542 ,n32[13]);
    nand g2408(n3427 ,n3341 ,n3273);
    nand g2409(n3147 ,n2764 ,n3075);
    nor g2410(n515 ,n468 ,n514);
    nand g2411(n3098 ,n2785 ,n2937);
    nand g2412(n1497 ,n1110 ,n1112);
    nor g2413(n71 ,n6[19] ,n68);
    nand g2414(n1738 ,n6[18] ,n535);
    nand g2415(n1588 ,n1178 ,n1189);
    dff g2416(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2481), .Q(n23[5]));
    dff g2417(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3180), .Q(n9[30]));
    nand g2418(n3307 ,n3220 ,n21[23]);
    nand g2419(n1130 ,n31[10] ,n527);
    nor g2420(n3049 ,n2766 ,n3035);
    nand g2421(n2258 ,n21[24] ,n1951);
    not g2422(n538 ,n6[5]);
    nand g2423(n1234 ,n31[22] ,n1031);
    not g2424(n211 ,n210);
    nand g2425(n3182 ,n2989 ,n3054);
    nor g2426(n606 ,n26[1] ,n6[5]);
    nand g2427(n2086 ,n1482 ,n1424);
    nand g2428(n2901 ,n6[4] ,n2697);
    nand g2429(n1910 ,n23[1] ,n1465);
    nand g2430(n1774 ,n8[12] ,n536);
    dff g2431(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2348), .Q(n26[22]));
    xnor g2432(n3523 ,n194 ,n24[11]);
    nand g2433(n1171 ,n29[4] ,n529);
    nand g2434(n2336 ,n2054 ,n1757);
    nand g2435(n2424 ,n2201 ,n1944);
    nand g2436(n422 ,n3413 ,n380);
    nand g2437(n1383 ,n27[13] ,n522);
    nand g2438(n454 ,n451 ,n449);
    nand g2439(n806 ,n32[8] ,n558);
    dff g2440(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3218), .Q(n9[8]));
    nor g2441(n3162 ,n2230 ,n3136);
    not g2442(n337 ,n336);
    not g2443(n352 ,n3405);
    nand g2444(n3291 ,n3221 ,n21[15]);
    not g2445(n2752 ,n2735);
    xnor g2446(n3443 ,n344 ,n21[29]);
    nand g2447(n1793 ,n3457 ,n534);
    not g2448(n227 ,n226);
    nand g2449(n1502 ,n1204 ,n1073);
    nor g2450(n699 ,n564 ,n32[9]);
    nand g2451(n1992 ,n30[16] ,n520);
    nand g2452(n2383 ,n1607 ,n1825);
    nand g2453(n1775 ,n3441 ,n534);
    or g2454(n876 ,n635 ,n657);
    nand g2455(n3041 ,n2734 ,n2852);
    nand g2456(n248 ,n22[8] ,n247);
    dff g2457(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2511), .Q(n24[18]));
    not g2458(n181 ,n180);
    nand g2459(n3430 ,n3303 ,n3236);
    not g2460(n531 ,n1146);
    nor g2461(n936 ,n615 ,n600);
    dff g2462(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1996), .Q(n27[15]));
    nand g2463(n1328 ,n31[11] ,n1146);
    nand g2464(n3111 ,n2798 ,n2950);
    nand g2465(n2897 ,n1187 ,n2701);
    dff g2466(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2472), .Q(n28[28]));
    or g2467(n696 ,n564 ,n29[9]);
    nand g2468(n1356 ,n29[17] ,n1147);
    nor g2469(n2920 ,n567 ,n2693);
    nand g2470(n952 ,n89 ,n668);
    nand g2471(n47 ,n6[26] ,n6[25]);
    or g2472(n419 ,n365 ,n3428);
    dff g2473(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3104), .Q(n10[14]));
    dff g2474(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2022), .Q(n29[16]));
    nand g2475(n3180 ,n2985 ,n3052);
    nand g2476(n2088 ,n1584 ,n1412);
    nand g2477(n1396 ,n3362 ,n1148);
    nand g2478(n1946 ,n32[0] ,n1462);
    nand g2479(n1336 ,n31[5] ,n1146);
    xor g2480(n3502 ,n22[1] ,n22[0]);
    nand g2481(n1998 ,n30[11] ,n520);
    nand g2482(n3240 ,n23[11] ,n3219);
    xnor g2483(n3461 ,n310 ,n21[11]);
    nand g2484(n1613 ,n3496 ,n530);
    nand g2485(n2888 ,n1081 ,n2683);
    nand g2486(n919 ,n656 ,n782);
    nand g2487(n726 ,n30[22] ,n550);
    nand g2488(n2676 ,n7[18] ,n2642);
    nand g2489(n3322 ,n3221 ,n21[31]);
    nand g2490(n779 ,n29[12] ,n543);
    dff g2491(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2662), .Q(n35[3]));
    or g2492(n2585 ,n1043 ,n2582);
    nand g2493(n242 ,n22[5] ,n241);
    not g2494(n2750 ,n2729);
    dff g2495(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3167), .Q(n9[9]));
    dff g2496(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1959), .Q(n31[18]));
    nand g2497(n2432 ,n2192 ,n1738);
    nor g2498(n1029 ,n861 ,n970);
    nand g2499(n1534 ,n1125 ,n1186);
    nand g2500(n1978 ,n1338 ,n1491);
    nand g2501(n2677 ,n7[17] ,n2642);
    nand g2502(n1203 ,n29[18] ,n529);
    nand g2503(n3338 ,n3220 ,n21[8]);
    nor g2504(n949 ,n538 ,n713);
    nand g2505(n983 ,n665 ,n802);
    not g2506(n234 ,n233);
    nand g2507(n1700 ,n6[27] ,n536);
    xnor g2508(n3513 ,n212 ,n24[21]);
    xnor g2509(n3519 ,n202 ,n24[15]);
    dff g2510(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1969), .Q(n31[11]));
    dff g2511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n847), .Q(n20[1]));
    nand g2512(n2301 ,n24[13] ,n1950);
    nand g2513(n1086 ,n1039 ,n1018);
    nand g2514(n1269 ,n6[13] ,n530);
    or g2515(n661 ,n562 ,n30[6]);
    nand g2516(n2863 ,n27[1] ,n2694);
    nand g2517(n1546 ,n1234 ,n1135);
    nand g2518(n1232 ,n27[7] ,n527);
    nand g2519(n82 ,n6[25] ,n77);
    nand g2520(n1102 ,n31[8] ,n1031);
    nand g2521(n2864 ,n27[2] ,n2694);
    nand g2522(n1000 ,n813 ,n754);
    nand g2523(n2426 ,n2198 ,n1742);
    nand g2524(n1001 ,n812 ,n768);
    nand g2525(n3287 ,n3220 ,n21[13]);
    dff g2526(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3217), .Q(n9[23]));
    nand g2527(n144 ,n23[14] ,n143);
    nand g2528(n2331 ,n2002 ,n1706);
    nand g2529(n2794 ,n10[11] ,n525);
    nand g2530(n783 ,n30[7] ,n561);
    nand g2531(n1416 ,n32[0] ,n1149);
    dff g2532(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2447), .Q(n32[23]));
    nand g2533(n1968 ,n1326 ,n1488);
    nand g2534(n1759 ,n8[28] ,n537);
    dff g2535(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1984), .Q(n27[20]));
    nor g2536(n2602 ,n3566 ,n2600);
    not g2537(n573 ,n34[3]);
    nand g2538(n917 ,n633 ,n806);
    xnor g2539(n3534 ,n174 ,n23[31]);
    nand g2540(n1253 ,n27[20] ,n1146);
    nand g2541(n2286 ,n24[28] ,n1950);
    dff g2542(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2411), .Q(n23[23]));
    nand g2543(n2808 ,n25[30] ,n2696);
    xnor g2544(n3442 ,n346 ,n21[30]);
    nor g2545(n412 ,n385 ,n3410);
    dff g2546(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2512), .Q(n21[3]));
    nand g2547(n1290 ,n6[20] ,n533);
    dff g2548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2510), .Q(n24[19]));
    nand g2549(n3038 ,n2731 ,n2913);
    nand g2550(n2312 ,n24[2] ,n1950);
    nand g2551(n3134 ,n1692 ,n2979);
    nand g2552(n512 ,n459 ,n511);
    xor g2553(n3372 ,n6[27] ,n80);
    nand g2554(n1782 ,n3448 ,n534);
    nand g2555(n2566 ,n1028 ,n2236);
    nor g2556(n417 ,n361 ,n3415);
    nand g2557(n2638 ,n844 ,n2610);
    nand g2558(n276 ,n22[23] ,n275);
    nand g2559(n1295 ,n6[23] ,n533);
    nand g2560(n2735 ,n11[5] ,n2641);
    nand g2561(n2803 ,n10[2] ,n2690);
    nand g2562(n1881 ,n23[30] ,n1465);
    dff g2563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2388), .Q(n22[12]));
    not g2564(n354 ,n3391);
    nor g2565(n2953 ,n1533 ,n2896);
    nand g2566(n2488 ,n1648 ,n1899);
    dff g2567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n851), .Q(n20[2]));
    nand g2568(n955 ,n708 ,n790);
    not g2569(n533 ,n1147);
    nand g2570(n1605 ,n3485 ,n531);
    nand g2571(n1082 ,n941 ,n1033);
    nand g2572(n437 ,n3398 ,n360);
    nand g2573(n1302 ,n6[31] ,n533);
    nand g2574(n2910 ,n27[9] ,n2694);
    nand g2575(n1732 ,n6[24] ,n534);
    or g2576(n871 ,n637 ,n689);
    nand g2577(n1072 ,n943 ,n1033);
    nand g2578(n3003 ,n9[12] ,n2848);
    nand g2579(n2198 ,n32[8] ,n523);
    dff g2580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3200), .Q(n11[10]));
    nor g2581(n106 ,n35[1] ,n35[0]);
    nand g2582(n3317 ,n3221 ,n22[14]);
    nor g2583(n471 ,n461 ,n458);
    nand g2584(n966 ,n747 ,n777);
    nand g2585(n2022 ,n1405 ,n1282);
    dff g2586(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n845), .Q(n20[0]));
    nand g2587(n342 ,n21[27] ,n341);
    nand g2588(n3008 ,n9[7] ,n2848);
    nand g2589(n3398 ,n3304 ,n3238);
    nand g2590(n3312 ,n3220 ,n21[26]);
    nand g2591(n2084 ,n1460 ,n1300);
    nand g2592(n749 ,n31[16] ,n546);
    nand g2593(n1905 ,n23[6] ,n1465);
    dff g2594(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2131), .Q(n25[13]));
    nand g2595(n1275 ,n6[7] ,n531);
    nand g2596(n2972 ,n6[17] ,n2849);
    xnor g2597(n3504 ,n230 ,n24[30]);
    nand g2598(n1680 ,n8[6] ,n533);
    nor g2599(n608 ,n538 ,n28[15]);
    nand g2600(n2057 ,n1448 ,n1380);
    nand g2601(n3349 ,n3221 ,n21[12]);
    xnor g2602(n3488 ,n260 ,n22[15]);
    not g2603(n535 ,n1462);
    nand g2604(n2850 ,n716 ,n2697);
    dff g2605(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2435), .Q(n32[14]));
    nor g2606(n1058 ,n862 ,n919);
    nand g2607(n2771 ,n928 ,n2692);
    nand g2608(n3274 ,n24[7] ,n3222);
    nor g2609(n2570 ,n1583 ,n2250);
    nand g2610(n2389 ,n1610 ,n1832);
    nand g2611(n3018 ,n2811 ,n2757);
    nor g2612(n264 ,n235 ,n262);
    nand g2613(n2634 ,n832 ,n2610);
    nand g2614(n1377 ,n27[16] ,n522);
    nand g2615(n1057 ,n868 ,n893);
    not g2616(n356 ,n3434);
    not g2617(n831 ,n830);
    dff g2618(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2536), .Q(n21[11]));
    nand g2619(n312 ,n21[11] ,n311);
    nor g2620(n3160 ,n2228 ,n3133);
    xnor g2621(n895 ,n556 ,n31[19]);
    nand g2622(n2486 ,n1651 ,n1901);
    nor g2623(n2657 ,n2601 ,n2628);
    dff g2624(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2455), .Q(n28[13]));
    nand g2625(n2594 ,n2593 ,n2589);
    nand g2626(n3346 ,n3220 ,n22[30]);
    nand g2627(n1879 ,n3533 ,n537);
    dff g2628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2012), .Q(n29[24]));
    not g2629(n257 ,n256);
    not g2630(n50 ,n49);
    nand g2631(n1764 ,n8[23] ,n536);
    nand g2632(n2234 ,n1694 ,n1248);
    nand g2633(n260 ,n22[14] ,n259);
    xnor g2634(n3549 ,n146 ,n23[16]);
    dff g2635(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2654), .Q(n34[4]));
    nand g2636(n2708 ,n1199 ,n2641);
    nand g2637(n1300 ,n6[6] ,n531);
    nand g2638(n1074 ,n942 ,n1033);
    or g2639(n1027 ,n871 ,n916);
    nand g2640(n272 ,n22[21] ,n271);
    not g2641(n361 ,n3383);
    nand g2642(n2379 ,n1604 ,n1823);
    nand g2643(n2285 ,n24[29] ,n1950);
    not g2644(n374 ,n3424);
    nand g2645(n1363 ,n29[3] ,n1147);
    nor g2646(n2943 ,n1514 ,n2886);
    nand g2647(n1493 ,n8[20] ,n530);
    nand g2648(n1164 ,n29[8] ,n529);
    nand g2649(n1516 ,n1236 ,n1237);
    nand g2650(n1801 ,n3465 ,n534);
    dff g2651(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3206), .Q(n9[6]));
    xnor g2652(n3497 ,n242 ,n22[6]);
    xor g2653(n3370 ,n6[25] ,n77);
    nand g2654(n3242 ,n24[23] ,n3219);
    nand g2655(n810 ,n28[24] ,n6[5]);
    dff g2656(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2130), .Q(n25[14]));
    xnor g2657(n3505 ,n228 ,n24[29]);
    nand g2658(n1505 ,n8[12] ,n530);
    nand g2659(n1373 ,n27[0] ,n1146);
    nand g2660(n2003 ,n30[5] ,n520);
    nand g2661(n1368 ,n32[25] ,n1149);
    nand g2662(n2133 ,n1447 ,n1673);
    nor g2663(n3086 ,n2754 ,n3045);
    nand g2664(n1258 ,n6[26] ,n530);
    nand g2665(n2308 ,n24[6] ,n1950);
    nand g2666(n2986 ,n9[29] ,n2848);
    dff g2667(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3184), .Q(n9[24]));
    nor g2668(n3068 ,n2831 ,n3026);
    or g2669(n2317 ,n1540 ,n2042);
    nand g2670(n1442 ,n29[18] ,n1147);
    nand g2671(n2914 ,n25[10] ,n2696);
    dff g2672(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3092), .Q(n10[26]));
    nand g2673(n2457 ,n2164 ,n1930);
    nand g2674(n1517 ,n1230 ,n1226);
    nand g2675(n1804 ,n3469 ,n535);
    nand g2676(n3298 ,n3221 ,n22[26]);
    nand g2677(n3432 ,n3319 ,n3253);
    nand g2678(n915 ,n669 ,n765);
    nand g2679(n2790 ,n10[15] ,n525);
    nand g2680(n2855 ,n25[5] ,n2696);
    nand g2681(n2536 ,n1797 ,n2271);
    not g2682(n259 ,n258);
    dff g2683(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2340), .Q(n26[29]));
    nand g2684(n2393 ,n2108 ,n1836);
    nor g2685(n2235 ,n1051 ,n1751);
    nand g2686(n1105 ,n27[0] ,n1031);
    xnor g2687(n3530 ,n180 ,n24[4]);
    not g2688(n383 ,n3415);
    nand g2689(n826 ,n89 ,n1);
    nand g2690(n2506 ,n1856 ,n2291);
    nor g2691(n462 ,n448 ,n444);
    not g2692(n365 ,n3396);
    dff g2693(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2473), .Q(n30[11]));
    nand g2694(n2477 ,n1662 ,n1910);
    nand g2695(n1935 ,n8[10] ,n535);
    nand g2696(n2734 ,n11[6] ,n2641);
    nor g2697(n2825 ,n1006 ,n2691);
    nand g2698(n1645 ,n3550 ,n532);
    nor g2699(n480 ,n457 ,n475);
    nand g2700(n2797 ,n10[8] ,n2690);
    nand g2701(n1498 ,n1240 ,n1113);
    dff g2702(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2525), .Q(n24[4]));
    nand g2703(n1926 ,n8[19] ,n534);
    nand g2704(n1883 ,n23[28] ,n1465);
    nand g2705(n1333 ,n27[23] ,n522);
    nand g2706(n1877 ,n3531 ,n537);
    nand g2707(n2282 ,n21[0] ,n1951);
    nor g2708(n689 ,n554 ,n32[11]);
    nand g2709(n1809 ,n8[6] ,n536);
    buf g2710(n19[3], 1'b0);
    nor g2711(n638 ,n559 ,n32[14]);
    nand g2712(n3090 ,n2776 ,n2928);
    nor g2713(n2936 ,n1506 ,n2879);
    nor g2714(n2767 ,n931 ,n2691);
    dff g2715(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3169), .Q(n11[29]));
    xnor g2716(n3477 ,n280 ,n22[26]);
    nor g2717(n796 ,n584 ,n539);
    nand g2718(n1975 ,n1333 ,n1490);
    nand g2719(n1301 ,n6[25] ,n533);
    nand g2720(n1575 ,n30[6] ,n1150);
    nand g2721(n973 ,n690 ,n770);
    dff g2722(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2523), .Q(n24[6]));
    nand g2723(n2671 ,n7[23] ,n2642);
    nand g2724(n3017 ,n2719 ,n2866);
    nand g2725(n1184 ,n27[22] ,n1031);
    nand g2726(n2725 ,n11[15] ,n2641);
    nand g2727(n795 ,n32[15] ,n541);
    xnor g2728(n3538 ,n166 ,n23[27]);
    nand g2729(n1569 ,n1130 ,n1159);
    nand g2730(n198 ,n24[12] ,n197);
    dff g2731(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2408), .Q(n23[26]));
    nand g2732(n2639 ,n857 ,n2610);
    nand g2733(n2113 ,n1427 ,n1622);
    nand g2734(n1371 ,n29[1] ,n521);
    dff g2735(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3203), .Q(n9[10]));
    nand g2736(n2475 ,n2136 ,n1913);
    nor g2737(n2951 ,n1529 ,n2894);
    nand g2738(n1229 ,n25[14] ,n1032);
    dff g2739(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2321), .Q(n30[18]));
    nand g2740(n1674 ,n8[10] ,n532);
    not g2741(n2742 ,n2706);
    not g2742(n2597 ,n2598);
    nand g2743(n728 ,n31[2] ,n565);
    not g2744(n2693 ,n2694);
    nand g2745(n519 ,n455 ,n518);
    nand g2746(n1703 ,n6[17] ,n536);
    nand g2747(n1666 ,n8[16] ,n533);
    or g2748(n2221 ,n1561 ,n2065);
    nand g2749(n2805 ,n10[0] ,n525);
    dff g2750(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3189), .Q(n11[21]));
    nand g2751(n2339 ,n2048 ,n1713);
    nand g2752(n3347 ,n3221 ,n22[31]);
    nand g2753(n2736 ,n11[4] ,n2641);
    nand g2754(n2704 ,n7[0] ,n2642);
    dff g2755(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2162), .Q(n25[3]));
    nand g2756(n1565 ,n1213 ,n1224);
    nand g2757(n1281 ,n6[27] ,n533);
    dff g2758(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2024), .Q(n27[6]));
    nand g2759(n1154 ,n31[4] ,n1031);
    dff g2760(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2360), .Q(n26[11]));
    nand g2761(n1292 ,n6[21] ,n532);
    nand g2762(n1720 ,n6[19] ,n537);
    nand g2763(n2453 ,n2169 ,n1934);
    nand g2764(n2280 ,n21[2] ,n1951);
    nand g2765(n3037 ,n2730 ,n2914);
    nand g2766(n240 ,n22[4] ,n239);
    dff g2767(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1982), .Q(n27[21]));
    nand g2768(n1073 ,n938 ,n1033);
    nand g2769(n3042 ,n2855 ,n2854);
    dff g2770(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2445), .Q(n32[22]));
    nand g2771(n1303 ,n6[26] ,n532);
    nand g2772(n1693 ,n1311 ,n1255);
    not g2773(n191 ,n190);
    nand g2774(n1794 ,n3458 ,n534);
    nand g2775(n1504 ,n1183 ,n1193);
    xnor g2776(n3518 ,n204 ,n24[16]);
    nor g2777(n2962 ,n555 ,n2850);
    nand g2778(n1604 ,n3484 ,n531);
    nor g2779(n635 ,n549 ,n30[17]);
    nand g2780(n2552 ,n1778 ,n2254);
    nand g2781(n3411 ,n3330 ,n3268);
    nand g2782(n244 ,n22[6] ,n243);
    nand g2783(n1880 ,n23[31] ,n1465);
    not g2784(n557 ,n6[26]);
    dff g2785(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2515), .Q(n24[14]));
    nand g2786(n1340 ,n31[2] ,n522);
    nand g2787(n86 ,n6[29] ,n84);
    not g2788(n255 ,n254);
    xnor g2789(n3352 ,n6[7] ,n42);
    dff g2790(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2527), .Q(n24[2]));
    nand g2791(n284 ,n22[27] ,n283);
    nand g2792(n2726 ,n11[14] ,n2641);
    nand g2793(n1783 ,n3449 ,n535);
    nand g2794(n2983 ,n6[6] ,n2849);
    nand g2795(n1834 ,n22[10] ,n1464);
    nand g2796(n2314 ,n24[0] ,n1950);
    nand g2797(n759 ,n32[0] ,n540);
    nand g2798(n1835 ,n22[9] ,n1464);
    nor g2799(n2656 ,n2606 ,n2627);
    xnor g2800(n3354 ,n6[9] ,n53);
    nand g2801(n1753 ,n907 ,n1306);
    or g2802(n479 ,n456 ,n478);
    nand g2803(n3394 ,n3294 ,n3231);
    nand g2804(n762 ,n26[20] ,n538);
    nor g2805(n1243 ,n910 ,n1099);
    nand g2806(n2717 ,n11[23] ,n2641);
    dff g2807(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2542), .Q(n21[17]));
    not g2808(n165 ,n164);
    xnor g2809(n3375 ,n6[30] ,n86);
    nand g2810(n3248 ,n23[13] ,n3222);
    dff g2811(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2353), .Q(n26[18]));
    nor g2812(n1306 ,n1041 ,n1091);
    nand g2813(n330 ,n21[21] ,n329);
    nand g2814(n1839 ,n22[6] ,n1464);
    dff g2815(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2534), .Q(n21[9]));
    xnor g2816(n3543 ,n156 ,n23[22]);
    nand g2817(n1309 ,n27[30] ,n1146);
    nand g2818(n2450 ,n2174 ,n1725);
    nor g2819(n662 ,n542 ,n29[13]);
    nand g2820(n2346 ,n2069 ,n1763);
    nand g2821(n306 ,n21[8] ,n305);
    or g2822(n2237 ,n1750 ,n1244);
    not g2823(n345 ,n344);
    nand g2824(n1587 ,n30[1] ,n1150);
    nand g2825(n920 ,n648 ,n803);
    nand g2826(n1623 ,n8[28] ,n533);
    nand g2827(n74 ,n6[20] ,n73);
    nand g2828(n1512 ,n1215 ,n1238);
    nand g2829(n1093 ,n1013 ,n1030);
    nand g2830(n2815 ,n27[27] ,n2694);
    nand g2831(n1866 ,n3521 ,n536);
    not g2832(n292 ,n291);
    not g2833(n539 ,n1);
    nand g2834(n2326 ,n1994 ,n1720);
    nand g2835(n496 ,n434 ,n495);
    nor g2836(n641 ,n555 ,n31[21]);
    nand g2837(n2534 ,n1833 ,n2273);
    nor g2838(n2940 ,n1511 ,n2883);
    dff g2839(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2390), .Q(n22[10]));
    not g2840(n350 ,n3406);
    nand g2841(n1173 ,n25[9] ,n529);
    nand g2842(n2075 ,n1400 ,n1461);
    nor g2843(n2834 ,n581 ,n2693);
    nand g2844(n998 ,n809 ,n721);
    dff g2845(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1975), .Q(n27[23]));
    nand g2846(n3117 ,n2804 ,n2956);
    nand g2847(n3318 ,n3220 ,n22[6]);
    nand g2848(n2975 ,n6[14] ,n2849);
    not g2849(n388 ,n3380);
    nand g2850(n2255 ,n21[27] ,n1951);
    nand g2851(n1429 ,n25[27] ,n521);
    nand g2852(n1094 ,n1055 ,n1048);
    nand g2853(n393 ,n3422 ,n370);
    dff g2854(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2072), .Q(n27[18]));
    nand g2855(n1167 ,n29[6] ,n1032);
    dff g2856(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2015), .Q(n29[21]));
    nand g2857(n909 ,n658 ,n746);
    nor g2858(n2843 ,n582 ,n2695);
    nand g2859(n3409 ,n3324 ,n3261);
    dff g2860(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3142), .Q(n9[3]));
    nand g2861(n3198 ,n2816 ,n3048);
    nand g2862(n1359 ,n27[4] ,n1146);
    xnor g2863(n3499 ,n238 ,n22[4]);
    nand g2864(n1214 ,n25[28] ,n529);
    nand g2865(n2832 ,n27[21] ,n2694);
    nand g2866(n3116 ,n2803 ,n2955);
    dff g2867(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1970), .Q(n31[10]));
    nand g2868(n2487 ,n1649 ,n1900);
    nand g2869(n2038 ,n1373 ,n1541);
    nand g2870(n1920 ,n4 ,n1467);
    nor g2871(n2927 ,n1520 ,n2870);
    dff g2872(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3088), .Q(n10[30]));
    xnor g2873(n3456 ,n320 ,n21[16]);
    nand g2874(n739 ,n29[21] ,n555);
    nand g2875(n2981 ,n6[8] ,n2849);
    nand g2876(n844 ,n35[0] ,n1);
    nor g2877(n3152 ,n2221 ,n3125);
    nand g2878(n784 ,n28[3] ,n6[5]);
    dff g2879(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2470), .Q(n28[26]));
    nand g2880(n2291 ,n24[23] ,n1950);
    dff g2881(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3117), .Q(n10[1]));
    nand g2882(n808 ,n29[3] ,n560);
    nand g2883(n2857 ,n25[4] ,n2696);
    nand g2884(n2549 ,n1782 ,n2258);
    dff g2885(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2123), .Q(n25[20]));
    nand g2886(n791 ,n29[11] ,n554);
    nand g2887(n3099 ,n2786 ,n2938);
    nand g2888(n3306 ,n3221 ,n22[11]);
    nand g2889(n3382 ,n3332 ,n3255);
    nor g2890(n2766 ,n932 ,n2691);
    nand g2891(n2131 ,n1444 ,n1671);
    nand g2892(n2621 ,n830 ,n2609);
    nand g2893(n2780 ,n10[25] ,n525);
    nand g2894(n1840 ,n22[5] ,n1464);
    nand g2895(n1211 ,n1008 ,n1033);
    nand g2896(n1398 ,n32[10] ,n1149);
    nand g2897(n1831 ,n3462 ,n534);
    nand g2898(n2087 ,n1358 ,n1527);
    nand g2899(n1904 ,n23[7] ,n1465);
    nand g2900(n824 ,n91 ,n1);
    nor g2901(n3066 ,n2825 ,n3024);
    nand g2902(n3207 ,n3001 ,n3158);
    nand g2903(n1944 ,n8[1] ,n535);
    dff g2904(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2492), .Q(n23[16]));
    nand g2905(n1437 ,n25[18] ,n521);
    nand g2906(n2281 ,n21[1] ,n1951);
    dff g2907(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1956), .Q(n31[20]));
    or g2908(n3167 ,n2980 ,n3135);
    nand g2909(n3341 ,n3220 ,n22[18]);
    dff g2910(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3176), .Q(n11[5]));
    nand g2911(n3022 ,n2820 ,n2819);
    nand g2912(n2092 ,n26[16] ,n520);
    nand g2913(n729 ,n31[20] ,n557);
    nand g2914(n1262 ,n6[21] ,n530);
    nand g2915(n1212 ,n27[30] ,n527);
    nand g2916(n2529 ,n1803 ,n2278);
    dff g2917(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2035), .Q(n27[2]));
    nand g2918(n1305 ,n6[18] ,n533);
    nand g2919(n2719 ,n11[0] ,n2641);
    nand g2920(n2093 ,n26[15] ,n1463);
    nand g2921(n1833 ,n3463 ,n534);
    xnor g2922(n3469 ,n294 ,n21[3]);
    nand g2923(n2978 ,n6[11] ,n2849);
    nand g2924(n2028 ,n1420 ,n1297);
    nand g2925(n1444 ,n25[13] ,n1147);
    nand g2926(n484 ,n415 ,n481);
    nor g2927(n613 ,n538 ,n28[27]);
    xnor g2928(n3366 ,n6[21] ,n74);
    nand g2929(n2283 ,n24[31] ,n1950);
    nand g2930(n778 ,n26[23] ,n538);
    nand g2931(n2526 ,n1877 ,n2311);
    nand g2932(n2330 ,n2163 ,n1724);
    nand g2933(n1296 ,n6[17] ,n532);
    nor g2934(n3164 ,n2232 ,n3138);
    nor g2935(n485 ,n464 ,n480);
    nand g2936(n2150 ,n28[22] ,n523);
    nand g2937(n1439 ,n27[9] ,n522);
    dff g2938(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2485), .Q(n23[9]));
    nand g2939(n733 ,n31[6] ,n562);
    nand g2940(n296 ,n21[3] ,n295);
    nand g2941(n2903 ,n6[2] ,n2697);
    dff g2942(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2111), .Q(n25[31]));
    nand g2943(n3421 ,n3309 ,n3243);
    nand g2944(n2724 ,n11[16] ,n2641);
    nand g2945(n2064 ,n1391 ,n1558);
    not g2946(n2748 ,n2722);
    or g2947(n2224 ,n1569 ,n2074);
    nand g2948(n3002 ,n9[13] ,n2848);
    nand g2949(n495 ,n431 ,n494);
    nand g2950(n3145 ,n2758 ,n3062);
    nor g2951(n1247 ,n977 ,n1064);
    nand g2952(n2053 ,n1547 ,n1375);
    nand g2953(n460 ,n398 ,n394);
    nand g2954(n1185 ,n25[21] ,n1032);
    nand g2955(n1042 ,n902 ,n903);
    nor g2956(n614 ,n538 ,n28[25]);
    nand g2957(n1761 ,n8[26] ,n537);
    nand g2958(n1563 ,n1155 ,n1233);
    nand g2959(n2830 ,n1003 ,n2692);
    nand g2960(n1176 ,n996 ,n1033);
    nand g2961(n3209 ,n2998 ,n3155);
    nand g2962(n1818 ,n22[22] ,n1464);
    nand g2963(n2732 ,n11[8] ,n2641);
    nand g2964(n2683 ,n7[12] ,n2642);
    not g2965(n570 ,n25[7]);
    nand g2966(n1067 ,n944 ,n1033);
    dff g2967(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1966), .Q(n27[26]));
    nand g2968(n2915 ,n1008 ,n2692);
    nand g2969(n3278 ,n23[25] ,n3222);
    nand g2970(n2600 ,n937 ,n2596);
    xor g2971(n3533 ,n24[1] ,n24[0]);
    nand g2972(n2325 ,n2160 ,n1723);
    not g2973(n569 ,n25[31]);
    nand g2974(n3283 ,n23[6] ,n3222);
    nand g2975(n2869 ,n1134 ,n2699);
    not g2976(n366 ,n3403);
    nand g2977(n2680 ,n7[14] ,n2642);
    nand g2978(n2032 ,n1361 ,n1283);
    nand g2979(n1318 ,n27[27] ,n522);
    nand g2980(n2892 ,n1173 ,n2686);
    dff g2981(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2331), .Q(n30[6]));
    dff g2982(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3114), .Q(n10[4]));
    nand g2983(n2155 ,n1419 ,n1496);
    xnor g2984(n3520 ,n200 ,n24[14]);
    dff g2985(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2355), .Q(n26[16]));
    nor g2986(n2696 ,n2589 ,n2641);
    xor g2987(n3454 ,n21[18] ,n322);
    nand g2988(n2384 ,n2107 ,n1827);
    nand g2989(n3261 ,n23[0] ,n3219);
    xor g2990(n862 ,n6[18] ,n30[12]);
    nand g2991(n1961 ,n1321 ,n1261);
    nand g2992(n3187 ,n2826 ,n3066);
    nand g2993(n1461 ,n3360 ,n1148);
    nand g2994(n2533 ,n1800 ,n2274);
    nand g2995(n160 ,n23[23] ,n159);
    nand g2996(n2207 ,n26[19] ,n520);
    nand g2997(n1770 ,n8[17] ,n536);
    nand g2998(n1985 ,n30[25] ,n1463);
    not g2999(n542 ,n6[19]);
    nor g3000(n3069 ,n2834 ,n3027);
    xor g3001(n3516 ,n24[18] ,n206);
    dff g3002(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2043), .Q(n27[1]));
    nand g3003(n3144 ,n2761 ,n3064);
    nand g3004(n2779 ,n10[26] ,n2690);
    nand g3005(n3113 ,n2800 ,n2952);
    nor g3006(n2568 ,n1497 ,n2243);
    xnor g3007(n3576 ,n35[3] ,n109);
    nand g3008(n2429 ,n2195 ,n1942);
    nand g3009(n1393 ,n32[14] ,n1149);
    nand g3010(n798 ,n12 ,n1);
    nand g3011(n2974 ,n6[15] ,n2849);
    xnor g3012(n3358 ,n6[13] ,n62);
    nor g3013(n2939 ,n1501 ,n2882);
    nand g3014(n1201 ,n27[25] ,n527);
    nand g3015(n1734 ,n6[22] ,n534);
    nor g3016(n2926 ,n1495 ,n2869);
    nand g3017(n867 ,n1 ,n720);
    nand g3018(n1618 ,n8[31] ,n533);
    nand g3019(n2307 ,n24[7] ,n1950);
    nand g3020(n3426 ,n3331 ,n3270);
    nand g3021(n2703 ,n7[1] ,n2642);
    nand g3022(n2139 ,n28[29] ,n523);
    nand g3023(n2518 ,n1867 ,n2302);
    not g3024(n2647 ,n2636);
    nand g3025(n1945 ,n8[0] ,n535);
    nand g3026(n3058 ,n3010 ,n2925);
    dff g3027(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3187), .Q(n11[23]));
    xnor g3028(n3490 ,n256 ,n22[13]);
    dff g3029(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2456), .Q(n28[14]));
    nand g3030(n1003 ,n786 ,n772);
    nand g3031(n2421 ,n2203 ,n1745);
    nand g3032(n3277 ,n24[9] ,n3222);
    dff g3033(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2031), .Q(n29[10]));
    or g3034(n628 ,n558 ,n30[8]);
    nor g3035(n518 ,n487 ,n517);
    xnor g3036(n3484 ,n266 ,n22[19]);
    nand g3037(n1123 ,n29[24] ,n529);
    nand g3038(n2991 ,n9[24] ,n2848);
    dff g3039(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2347), .Q(n26[23]));
    xnor g3040(n3559 ,n126 ,n23[6]);
    nand g3041(n3139 ,n2904 ,n3015);
    nand g3042(n1446 ,n27[19] ,n1146);
    nand g3043(n3332 ,n3220 ,n21[5]);
    nand g3044(n1584 ,n30[2] ,n1150);
    not g3045(n217 ,n216);
    nand g3046(n735 ,n31[17] ,n549);
    nand g3047(n1609 ,n3491 ,n530);
    nand g3048(n1938 ,n8[7] ,n535);
    nand g3049(n2250 ,n1582 ,n2216);
    nand g3050(n2921 ,n27[12] ,n2694);
    nand g3051(n1934 ,n8[11] ,n534);
    not g3052(n281 ,n280);
    nand g3053(n1635 ,n3542 ,n532);
    nand g3054(n1538 ,n1105 ,n1131);
    nand g3055(n180 ,n24[3] ,n179);
    nand g3056(n723 ,n29[22] ,n550);
    dff g3057(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2384), .Q(n26[3]));
    xnor g3058(n3446 ,n338 ,n21[26]);
    nand g3059(n3218 ,n3007 ,n3162);
    nand g3060(n3030 ,n2723 ,n2842);
    nor g3061(n1054 ,n864 ,n954);
    nand g3062(n1415 ,n27[12] ,n1146);
    nand g3063(n1564 ,n30[12] ,n1150);
    nor g3064(n1039 ,n870 ,n955);
    dff g3065(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2522), .Q(n24[7]));
    nand g3066(n1979 ,n1337 ,n1272);
    nand g3067(n1390 ,n3366 ,n1148);
    dff g3068(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2494), .Q(n23[18]));
    or g3069(n2569 ,n1548 ,n2244);
    nand g3070(n1143 ,n31[15] ,n527);
    nand g3071(n1657 ,n8[20] ,n533);
    dff g3072(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2437), .Q(n32[16]));
    nand g3073(n2670 ,n7[24] ,n2642);
    xnor g3074(n3371 ,n6[26] ,n82);
    not g3075(n219 ,n218);
    nand g3076(n3108 ,n2794 ,n2946);
    nand g3077(n3114 ,n2801 ,n2953);
    nand g3078(n2611 ,n35[0] ,n2597);
    not g3079(n559 ,n6[20]);
    nand g3080(n224 ,n24[26] ,n223);
    nand g3081(n1932 ,n8[13] ,n534);
    xnor g3082(n3491 ,n254 ,n22[12]);
    nand g3083(n3319 ,n3221 ,n22[23]);
    dff g3084(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2446), .Q(n28[7]));
    nand g3085(n2556 ,n1775 ,n2251);
    or g3086(n2575 ,n1549 ,n2245);
    nand g3087(n776 ,n29[15] ,n541);
    nand g3088(n2260 ,n21[22] ,n1951);
    nand g3089(n254 ,n22[11] ,n253);
    nand g3090(n3046 ,n2865 ,n2772);
    nor g3091(n2929 ,n1499 ,n2872);
    nand g3092(n1179 ,n25[26] ,n1032);
    or g3093(n648 ,n555 ,n30[21]);
    nand g3094(n37[0] ,n445 ,n519);
    dff g3095(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2560), .Q(n24[0]));
    nand g3096(n1230 ,n27[12] ,n1031);
    dff g3097(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2381), .Q(n22[17]));
    nand g3098(n1481 ,n27[31] ,n522);
    nand g3099(n2999 ,n9[16] ,n2848);
    nand g3100(n235 ,n22[17] ,n22[16]);
    nand g3101(n2034 ,n1364 ,n1284);
    nor g3102(n611 ,n538 ,n28[31]);
    nand g3103(n1984 ,n1253 ,n1493);
    nand g3104(n2050 ,n1349 ,n1542);
    dff g3105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2323), .Q(n30[1]));
    nand g3106(n1591 ,n3480 ,n530);
    nor g3107(n607 ,n26[25] ,n6[5]);
    nor g3108(n2694 ,n2593 ,n2641);
    dff g3109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2516), .Q(n24[11]));
    nor g3110(n476 ,n412 ,n470);
    not g3111(n568 ,n25[19]);
    nand g3112(n3431 ,n3311 ,n3241);
    nand g3113(n3342 ,n3220 ,n21[1]);
    nand g3114(n1410 ,n32[4] ,n1149);
    nand g3115(n1822 ,n8[4] ,n537);
    nand g3116(n3044 ,n2737 ,n2859);
    nand g3117(n2012 ,n1351 ,n1280);
    nand g3118(n2063 ,n26[25] ,n520);
    not g3119(n520 ,n537);
    nand g3120(n1643 ,n3548 ,n533);
    not g3121(n563 ,n6[7]);
    nand g3122(n2564 ,n1037 ,n2239);
    nand g3123(n1170 ,n27[24] ,n1031);
    nand g3124(n2186 ,n28[5] ,n523);
    not g3125(n96 ,n95);
    nor g3126(n2934 ,n1504 ,n2877);
    nor g3127(n935 ,n608 ,n602);
    nor g3128(n3059 ,n2806 ,n3016);
    nand g3129(n2702 ,n7[2] ,n2642);
    or g3130(n1250 ,n23[0] ,n521);
    nor g3131(n2952 ,n1531 ,n2895);
    not g3132(n521 ,n533);
    nand g3133(n1981 ,n1340 ,n1274);
    not g3134(n2749 ,n2724);
    nand g3135(n2094 ,n30[9] ,n520);
    dff g3136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1967), .Q(n31[12]));
    nand g3137(n2439 ,n2185 ,n1733);
    nand g3138(n1827 ,n8[3] ,n536);
    xnor g3139(n3460 ,n312 ,n21[12]);
    dff g3140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2495), .Q(n23[19]));
    nand g3141(n2171 ,n823 ,n523);
    nand g3142(n1160 ,n1007 ,n1033);
    xnor g3143(n3522 ,n196 ,n24[12]);
    not g3144(n380 ,n3381);
    not g3145(n267 ,n266);
    nand g3146(n1492 ,n8[21] ,n530);
    nand g3147(n1128 ,n27[20] ,n1031);
    nand g3148(n821 ,n28[5] ,n6[5]);
    nand g3149(n3344 ,n3220 ,n22[25]);
    nand g3150(n3401 ,n3308 ,n3244);
    not g3151(n522 ,n531);
    nand g3152(n3000 ,n9[15] ,n2848);
    nand g3153(n1719 ,n6[29] ,n536);
    nand g3154(n1585 ,n8[17] ,n531);
    not g3155(n327 ,n326);
    nand g3156(n228 ,n24[28] ,n227);
    nand g3157(n1124 ,n25[2] ,n529);
    nand g3158(n1750 ,n1243 ,n1092);
    nand g3159(n2973 ,n6[16] ,n2849);
    nand g3160(n3395 ,n3296 ,n3232);
    nand g3161(n3348 ,n3221 ,n21[11]);
    nand g3162(n2333 ,n2005 ,n1711);
    nand g3163(n1354 ,n29[19] ,n1147);
    nand g3164(n1539 ,n30[25] ,n1150);
    nand g3165(n1678 ,n8[8] ,n533);
    nor g3166(n51 ,n40 ,n45);
    nand g3167(n1559 ,n1143 ,n1111);
    nand g3168(n1181 ,n29[0] ,n1032);
    nand g3169(n2778 ,n10[27] ,n525);
    nand g3170(n2417 ,n2079 ,n1749);
    nand g3171(n2410 ,n1634 ,n1887);
    nand g3172(n1789 ,n3454 ,n534);
    dff g3173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3100), .Q(n10[18]));
    dff g3174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2656), .Q(n34[2]));
    nand g3175(n3414 ,n3345 ,n3279);
    not g3176(n285 ,n284);
    nand g3177(n2687 ,n7[8] ,n2642);
    nand g3178(n2122 ,n1422 ,n1654);
    nand g3179(n1688 ,n1231 ,n1179);
    nand g3180(n2837 ,n1000 ,n2692);
    nand g3181(n1687 ,n30[13] ,n1150);
    nand g3182(n2567 ,n884 ,n2235);
    nand g3183(n2787 ,n10[18] ,n2690);
    not g3184(n1036 ,n1035);
    nand g3185(n2812 ,n25[29] ,n2696);
    nand g3186(n922 ,n702 ,n764);
    nand g3187(n822 ,n28[22] ,n6[5]);
    nand g3188(n3112 ,n2799 ,n2951);
    nand g3189(n1991 ,n30[17] ,n1463);
    nor g3190(n2613 ,n3575 ,n2598);
    nand g3191(n1153 ,n994 ,n1033);
    nand g3192(n2116 ,n1476 ,n1626);
    dff g3193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2387), .Q(n22[13]));
    xnor g3194(n887 ,n6[16] ,n32[10]);
    xnor g3195(n3577 ,n35[2] ,n107);
    nand g3196(n763 ,n29[13] ,n542);
    nand g3197(n1594 ,n3473 ,n531);
    nand g3198(n210 ,n24[19] ,n209);
    nand g3199(n1310 ,n31[24] ,n1146);
    nand g3200(n1425 ,n25[31] ,n521);
    nor g3201(n1754 ,n1246 ,n1096);
    nand g3202(n1644 ,n3549 ,n532);
    nand g3203(n1414 ,n32[1] ,n1149);
    dff g3204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2017), .Q(n29[20]));
    not g3205(n589 ,n34[5]);
    dff g3206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3215), .Q(n9[15]));
    nor g3207(n1044 ,n882 ,n979);
    nand g3208(n2277 ,n21[5] ,n1951);
    dff g3209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2351), .Q(n30[5]));
    nor g3210(n85 ,n6[29] ,n84);
    nand g3211(n1597 ,n3476 ,n531);
    dff g3212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3171), .Q(n11[24]));
    not g3213(n163 ,n162);
    dff g3214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3209), .Q(n9[17]));
    nand g3215(n2722 ,n11[18] ,n2641);
    nand g3216(n2247 ,n1553 ,n2213);
    nand g3217(n3177 ,n2858 ,n3082);
    nand g3218(n1634 ,n3541 ,n532);
    dff g3219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2457), .Q(n28[15]));
    nand g3220(n1562 ,n1128 ,n1192);
    nand g3221(n2141 ,n1456 ,n1679);
    nand g3222(n1892 ,n23[19] ,n1465);
    not g3223(n303 ,n302);
    nand g3224(n1423 ,n25[22] ,n1147);
    nand g3225(n1908 ,n23[3] ,n1465);
    dff g3226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2549), .Q(n21[24]));
    nand g3227(n1098 ,n1058 ,n1047);
    nand g3228(n1249 ,n872 ,n1065);
    nand g3229(n3400 ,n3307 ,n3242);
    dff g3230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3095), .Q(n10[21]));
    nand g3231(n2128 ,n30[23] ,n520);
    not g3232(n849 ,n848);
    nand g3233(n725 ,n30[5] ,n544);
    not g3234(n105 ,n35[4]);
    nand g3235(n2844 ,n999 ,n2692);
    dff g3236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2414), .Q(n23[20]));
    nand g3237(n2982 ,n6[7] ,n2849);
    nand g3238(n2102 ,n26[8] ,n1463);
    nand g3239(n1282 ,n6[22] ,n532);
    nand g3240(n1008 ,n817 ,n805);
    nand g3241(n2836 ,n27[19] ,n2694);
    nand g3242(n3301 ,n3221 ,n22[10]);
    nand g3243(n2786 ,n10[19] ,n525);
    nand g3244(n2578 ,n2557 ,n2562);
    not g3245(n377 ,n3429);
    nor g3246(n517 ,n469 ,n516);
    buf g3247(n18[3], 1'b0);
    xor g3248(n3485 ,n22[18] ,n264);
    xnor g3249(n3473 ,n288 ,n22[30]);
    dff g3250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2466), .Q(n28[23]));
    not g3251(n2646 ,n2635);
    nand g3252(n2156 ,n28[19] ,n523);
    nand g3253(n439 ,n3418 ,n363);
    nand g3254(n1859 ,n3514 ,n536);
    nor g3255(n600 ,n26[17] ,n6[5]);
    nand g3256(n2166 ,n28[13] ,n1462);
    nand g3257(n3028 ,n2721 ,n2836);
    or g3258(n2223 ,n1567 ,n2070);
    nand g3259(n2077 ,n1402 ,n1572);
    nand g3260(n1104 ,n25[5] ,n529);
    dff g3261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2467), .Q(n28[24]));
    nand g3262(n3410 ,n3335 ,n3265);
    dff g3263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2427), .Q(n28[2]));
    nand g3264(n781 ,n29[25] ,n548);
    nand g3265(n1787 ,n3452 ,n534);
    nand g3266(n174 ,n23[30] ,n173);
    not g3267(n167 ,n166);
    nand g3268(n1386 ,n27[14] ,n1146);
    nand g3269(n1108 ,n25[17] ,n1032);
    dff g3270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2621), .Q(n16));
    nand g3271(n3334 ,n3220 ,n21[6]);
    nand g3272(n1405 ,n29[16] ,n521);
    nand g3273(n3233 ,n23[9] ,n3222);
    dff g3274(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2551), .Q(n21[26]));
    nand g3275(n1127 ,n25[4] ,n1032);
    dff g3276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2023), .Q(n29[15]));
    nand g3277(n1924 ,n8[21] ,n535);
    nand g3278(n3280 ,n24[0] ,n3222);
    dff g3279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2531), .Q(n21[6]));
    nand g3280(n2106 ,n26[4] ,n1463);
    xnor g3281(n905 ,n6[7] ,n29[1]);
    nand g3282(n2083 ,n1410 ,n1408);
    nand g3283(n2899 ,n1114 ,n2703);
    nand g3284(n2524 ,n1875 ,n2309);
    nand g3285(n777 ,n31[7] ,n561);
    not g3286(n43 ,n42);
    dff g3287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2373), .Q(n22[24]));
    nand g3288(n3333 ,n3220 ,n22[28]);
    nand g3289(n2609 ,n1 ,n2599);
    dff g3290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2404), .Q(n23[30]));
    nand g3291(n2517 ,n1866 ,n2301);
    dff g3292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3111), .Q(n10[7]));
    not g3293(n574 ,n33[2]);
    nand g3294(n988 ,n654 ,n731);
    nand g3295(n1364 ,n29[8] ,n521);
    nand g3296(n2412 ,n1636 ,n1889);
    nand g3297(n2667 ,n7[27] ,n2642);
    nand g3298(n3424 ,n3321 ,n3257);
    nand g3299(n813 ,n28[18] ,n6[5]);
    nand g3300(n398 ,n3407 ,n369);
    not g3301(n78 ,n77);
    or g3302(n1081 ,n932 ,n1034);
    nor g3303(n872 ,n638 ,n642);
    nand g3304(n1852 ,n3507 ,n537);
    nor g3305(n937 ,n33[1] ,n761);
    nand g3306(n1349 ,n32[23] ,n1149);
    nand g3307(n3244 ,n24[24] ,n3222);
    nor g3308(n3073 ,n2749 ,n3031);
    not g3309(n153 ,n152);
    dff g3310(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2429), .Q(n28[3]));
    nand g3311(n1895 ,n23[16] ,n1465);
    nand g3312(n3440 ,n3347 ,n3249);
    nand g3313(n2699 ,n7[31] ,n2642);
    nand g3314(n2561 ,n1695 ,n2282);
    xnor g3315(n3365 ,n6[20] ,n72);
    nand g3316(n3310 ,n3220 ,n21[25]);
    nand g3317(n3297 ,n3220 ,n22[9]);
    dff g3318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2444), .Q(n32[21]));
    not g3319(n2741 ,n2705);
    xnor g3320(n3445 ,n340 ,n21[27]);
    nor g3321(n1950 ,n539 ,n537);
    nand g3322(n423 ,n3437 ,n352);
    nand g3323(n2047 ,n1371 ,n1279);
    nand g3324(n3241 ,n23[22] ,n3222);
    buf g3325(n19[1], 1'b0);
    nand g3326(n2781 ,n10[24] ,n2690);
    nand g3327(n3435 ,n3298 ,n3223);
    nor g3328(n933 ,n618 ,n594);
    nand g3329(n2007 ,n1360 ,n1507);
    nand g3330(n3128 ,n1398 ,n2973);
    nand g3331(n175 ,n24[1] ,n24[0]);
    nor g3332(n2652 ,n2607 ,n2622);
    nand g3333(n3088 ,n2775 ,n2927);
    dff g3334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1971), .Q(n31[9]));
    nand g3335(n3406 ,n3350 ,n3266);
    not g3336(n309 ,n308);
    nand g3337(n2788 ,n10[17] ,n525);
    nand g3338(n1453 ,n32[12] ,n1149);
    nand g3339(n2328 ,n2094 ,n1715);
    nand g3340(n3340 ,n3220 ,n21[9]);
    not g3341(n273 ,n272);
    nand g3342(n2462 ,n2156 ,n1926);
    or g3343(n2593 ,n1307 ,n2592);
    nand g3344(n2111 ,n1425 ,n1618);
    dff g3345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2548), .Q(n21[23]));
    nor g3346(n941 ,n612 ,n599);
    not g3347(n546 ,n6[22]);
    nand g3348(n53 ,n6[8] ,n50);
    nand g3349(n1518 ,n8[7] ,n530);
    dff g3350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1957), .Q(n27[28]));
    nand g3351(n1304 ,n6[9] ,n533);
    nand g3352(n1567 ,n1157 ,n1200);
    nand g3353(n1964 ,n1324 ,n1291);
    or g3354(n894 ,n699 ,n685);
    nand g3355(n2909 ,n25[8] ,n2696);
    nand g3356(n2403 ,n1691 ,n1880);
    nand g3357(n2827 ,n27[22] ,n2694);
    or g3358(n2220 ,n1559 ,n2064);
    nand g3359(n1554 ,n1140 ,n1203);
    nand g3360(n984 ,n686 ,n763);
    nand g3361(n2801 ,n10[4] ,n2690);
    nand g3362(n2443 ,n2181 ,n1730);
    nand g3363(n2243 ,n1346 ,n2209);
    nand g3364(n2701 ,n7[3] ,n2642);
    or g3365(n889 ,n640 ,n682);
    nand g3366(n2509 ,n1859 ,n2294);
    or g3367(n2232 ,n1590 ,n2091);
    nand g3368(n977 ,n647 ,n727);
    nand g3369(n1285 ,n6[16] ,n533);
    not g3370(n75 ,n74);
    nand g3371(n2542 ,n1790 ,n2265);
    nand g3372(n2298 ,n24[16] ,n1950);
    nand g3373(n3350 ,n3221 ,n21[29]);
    nand g3374(n1136 ,n31[21] ,n1031);
    dff g3375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2000), .Q(n27[14]));
    nand g3376(n1916 ,n8[27] ,n535);
    dff g3377(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n837), .Q(n20[11]));
    nand g3378(n1765 ,n8[22] ,n536);
    not g3379(n371 ,n3404);
    nand g3380(n2176 ,n28[8] ,n523);
    nor g3381(n2690 ,n925 ,n2642);
    dff g3382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2513), .Q(n24[16]));
    nand g3383(n1156 ,n27[21] ,n527);
    nand g3384(n2249 ,n1543 ,n2215);
    nand g3385(n1286 ,n6[11] ,n532);
    dff g3386(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2120), .Q(n25[23]));
    nand g3387(n2154 ,n28[20] ,n523);
    nand g3388(n1649 ,n3554 ,n532);
    dff g3389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2502), .Q(n24[28]));
    not g3390(n843 ,n842);
    not g3391(n183 ,n182);
    dff g3392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2343), .Q(n26[26]));
    nand g3393(n2866 ,n27[0] ,n2694);
    nand g3394(n2406 ,n1630 ,n1883);
    or g3395(n878 ,n655 ,n646);
    or g3396(n1014 ,n6[5] ,n952);
    nand g3397(n2822 ,n1007 ,n2692);
    nand g3398(n1870 ,n3524 ,n537);
    nand g3399(n1034 ,n566 ,n925);
    nand g3400(n1263 ,n6[19] ,n531);
    nand g3401(n1142 ,n29[16] ,n529);
    nor g3402(n3077 ,n2750 ,n3036);
    not g3403(n560 ,n6[9]);
    nand g3404(n1379 ,n29[14] ,n521);
    nand g3405(n2800 ,n10[5] ,n525);
    not g3406(n205 ,n204);
    nand g3407(n1860 ,n3515 ,n537);
    nand g3408(n2069 ,n26[24] ,n520);
    nor g3409(n1012 ,n914 ,n974);
    nand g3410(n2274 ,n21[8] ,n1951);
    dff g3411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2394), .Q(n22[7]));
    nand g3412(n3323 ,n3221 ,n21[0]);
    dff g3413(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2652), .Q(n34[7]));
    nor g3414(n3079 ,n2751 ,n3039);
    nand g3415(n1941 ,n8[4] ,n534);
    nand g3416(n1099 ,n808 ,n1026);
    nand g3417(n1690 ,n3498 ,n531);
    not g3418(n525 ,n524);
    or g3419(n2231 ,n1588 ,n2090);
    nand g3420(n97 ,n34[2] ,n96);
    nand g3421(n2127 ,n1438 ,n1665);
    nand g3422(n2538 ,n1795 ,n2269);
    nand g3423(n962 ,n90 ,n722);
    dff g3424(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2432), .Q(n32[12]));
    nand g3425(n1751 ,n891 ,n1241);
    nand g3426(n3269 ,n24[4] ,n3222);
    nor g3427(n2946 ,n1519 ,n2889);
    nand g3428(n3136 ,n1411 ,n2981);
    not g3429(n2644 ,n2633);
    or g3430(n875 ,n670 ,n701);
    nand g3431(n2502 ,n1851 ,n2286);
    nand g3432(n304 ,n21[7] ,n303);
    nand g3433(n1220 ,n27[27] ,n1031);
    nor g3434(n206 ,n177 ,n204);
    nand g3435(n1763 ,n8[24] ,n537);
    nor g3436(n1694 ,n1249 ,n1086);
    nand g3437(n150 ,n23[18] ,n148);
    nor g3438(n694 ,n552 ,n32[4]);
    nand g3439(n2396 ,n1690 ,n1840);
    nor g3440(n943 ,n611 ,n597);
    not g3441(n315 ,n314);
    nand g3442(n1515 ,n8[8] ,n530);
    nor g3443(n2616 ,n3578 ,n2598);
    nand g3444(n1890 ,n23[21] ,n1465);
    not g3445(n580 ,n27[3]);
    nand g3446(n2768 ,n930 ,n2692);
    or g3447(n698 ,n552 ,n29[4]);
    nand g3448(n1691 ,n3534 ,n533);
    nor g3449(n3084 ,n2860 ,n3044);
    nand g3450(n156 ,n23[21] ,n155);
    nand g3451(n1960 ,n1320 ,n1260);
    nor g3452(n644 ,n557 ,n31[20]);
    nand g3453(n1448 ,n32[19] ,n1149);
    not g3454(n295 ,n294);
    nand g3455(n742 ,n30[25] ,n548);
    nand g3456(n72 ,n6[19] ,n68);
    nand g3457(n2459 ,n2161 ,n1929);
    nand g3458(n1125 ,n27[3] ,n1031);
    xnor g3459(n3545 ,n152 ,n23[20]);
    nand g3460(n2969 ,n6[20] ,n2849);
    nand g3461(n2099 ,n26[12] ,n1463);
    nor g3462(n701 ,n557 ,n30[20]);
    nand g3463(n1667 ,n8[19] ,n530);
    xnor g3464(n3496 ,n244 ,n22[7]);
    nand g3465(n188 ,n24[7] ,n187);
    nor g3466(n443 ,n363 ,n3418);
    nand g3467(n1041 ,n897 ,n905);
    dff g3468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2040), .Q(n12));
    nand g3469(n2173 ,n28[9] ,n1462);
    nand g3470(n1218 ,n31[19] ,n1031);
    xnor g3471(n3506 ,n226 ,n24[28]);
    nand g3472(n2289 ,n24[25] ,n1950);
    nand g3473(n1628 ,n3535 ,n532);
    nand g3474(n3094 ,n2781 ,n2933);
    nand g3475(n1208 ,n29[19] ,n1032);
    nand g3476(n1401 ,n3359 ,n1148);
    nand g3477(n1638 ,n3545 ,n532);
    nand g3478(n3200 ,n2912 ,n3050);
    nand g3479(n1315 ,n31[20] ,n1146);
    nand g3480(n1376 ,n32[21] ,n1149);
    nand g3481(n3387 ,n3343 ,n3230);
    dff g3482(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2464), .Q(n28[21]));
    nand g3483(n1841 ,n8[1] ,n537);
    nand g3484(n2135 ,n28[31] ,n1462);
    nand g3485(n2359 ,n2099 ,n1774);
    nand g3486(n218 ,n24[23] ,n217);
    not g3487(n2596 ,n2595);
    xnor g3488(n3531 ,n178 ,n24[3]);
    dff g3489(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1962), .Q(n31[15]));
    nand g3490(n1132 ,n31[25] ,n527);
    nand g3491(n2373 ,n1600 ,n1816);
    not g3492(n375 ,n3395);
    dff g3493(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2030), .Q(n29[11]));
    nand g3494(n985 ,n651 ,n723);
    not g3495(n213 ,n212);
    nand g3496(n465 ,n410 ,n407);
    nand g3497(n2147 ,n1458 ,n1680);
    xnor g3498(n3537 ,n168 ,n23[28]);
    nand g3499(n2279 ,n21[3] ,n1951);
    nand g3500(n1470 ,n25[1] ,n1147);
    nand g3501(n2700 ,n7[4] ,n2642);
    nand g3502(n1348 ,n29[10] ,n521);
    not g3503(n275 ,n274);
    nand g3504(n3183 ,n2990 ,n3055);
    dff g3505(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2357), .Q(n26[15]));
    nand g3506(n2765 ,n933 ,n2692);
    dff g3507(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2741), .Q(n35[0]));
    nand g3508(n1488 ,n8[25] ,n531);
    nand g3509(n2120 ,n1431 ,n1642);
    nand g3510(n1996 ,n1347 ,n1669);
    nor g3511(n682 ,n551 ,n31[24]);
    nand g3512(n789 ,n29[4] ,n552);
    nand g3513(n252 ,n22[10] ,n251);
    not g3514(n63 ,n62);
    nand g3515(n830 ,n16 ,n1);
    nand g3516(n55 ,n6[23] ,n51);
    nor g3517(n452 ,n441 ,n392);
    nand g3518(n2163 ,n30[7] ,n1463);
    not g3519(n123 ,n122);
    dff g3520(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2440), .Q(n28[6]));
    nand g3521(n2878 ,n1175 ,n2672);
    nand g3522(n1838 ,n22[7] ,n1464);
    nand g3523(n1825 ,n22[16] ,n1464);
    nand g3524(n996 ,n819 ,n769);
    xnor g3525(n3459 ,n314 ,n21[13]);
    nand g3526(n1137 ,n31[20] ,n527);
    dff g3527(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2122), .Q(n25[21]));
    dff g3528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3181), .Q(n9[27]));
    dff g3529(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2349), .Q(n26[21]));
    nor g3530(n1951 ,n539 ,n535);
    nand g3531(n2358 ,n2096 ,n1773);
    nand g3532(n2413 ,n1637 ,n1890);
    nand g3533(n2777 ,n10[28] ,n2690);
    nand g3534(n1661 ,n3563 ,n533);
    dff g3535(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2500), .Q(n24[27]));
    nand g3536(n2760 ,n939 ,n2692);
    nand g3537(n3010 ,n9[5] ,n2848);
    nand g3538(n1394 ,n3364 ,n1148);
    nor g3539(n80 ,n47 ,n78);
    nand g3540(n3412 ,n3336 ,n3272);
    nand g3541(n2467 ,n2145 ,n1919);
    nand g3542(n344 ,n21[28] ,n343);
    nand g3543(n1257 ,n6[27] ,n530);
    nand g3544(n2813 ,n27[28] ,n2694);
    nand g3545(n2295 ,n24[19] ,n1950);
    nand g3546(n2718 ,n11[22] ,n2641);
    nand g3547(n709 ,n31[18] ,n545);
    nor g3548(n703 ,n26[4] ,n6[5]);
    nand g3549(n2126 ,n1440 ,n1666);
    nor g3550(n1032 ,n834 ,n924);
    dff g3551(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1978), .Q(n27[22]));
    nand g3552(n3390 ,n3287 ,n3254);
    nand g3553(n2313 ,n24[1] ,n1950);
    or g3554(n627 ,n565 ,n32[2]);
    dff g3555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3098), .Q(n10[20]));
    nand g3556(n428 ,n3427 ,n375);
    nand g3557(n2497 ,n1807 ,n2281);
    nand g3558(n2772 ,n927 ,n2692);
    dff g3559(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2126), .Q(n25[16]));
    nand g3560(n2165 ,n28[14] ,n1462);
    nand g3561(n470 ,n403 ,n465);
    dff g3562(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3140), .Q(n9[0]));
    nand g3563(n1482 ,n32[3] ,n1149);
    xnor g3564(n3441 ,n348 ,n21[31]);
    nand g3565(n3253 ,n23[23] ,n3222);
    nor g3566(n700 ,n552 ,n31[4]);
    nor g3567(n100 ,n93 ,n99);
    nand g3568(n2172 ,n825 ,n520);
    nor g3569(n907 ,n645 ,n671);
    nand g3570(n1909 ,n23[2] ,n1465);
    not g3571(n223 ,n222);
    nand g3572(n2482 ,n1656 ,n1905);
    nand g3573(n3031 ,n2845 ,n2844);
    not g3574(n195 ,n194);
    nand g3575(n1836 ,n8[2] ,n536);
    dff g3576(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2504), .Q(n24[25]));
    dff g3577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3166), .Q(n9[13]));
    nand g3578(n722 ,n30[8] ,n558);
    nor g3579(n389 ,n359 ,n3420);
    dff g3580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2014), .Q(n29[22]));
    dff g3581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2521), .Q(n24[8]));
    nand g3582(n3095 ,n2784 ,n2936);
    not g3583(n558 ,n6[14]);
    nand g3584(n1200 ,n29[11] ,n1032);
    nand g3585(n168 ,n23[27] ,n167);
    nor g3586(n2828 ,n578 ,n2695);
    nand g3587(n1547 ,n30[21] ,n1150);
    nand g3588(n1911 ,n23[0] ,n1465);
    nand g3589(n1489 ,n8[24] ,n530);
    nand g3590(n3005 ,n9[10] ,n2848);
    nand g3591(n2338 ,n1988 ,n1700);
    nand g3592(n3299 ,n3220 ,n21[19]);
    nand g3593(n3211 ,n2994 ,n3153);
    dff g3594(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3201), .Q(n11[6]));
    nand g3595(n1792 ,n3456 ,n534);
    dff g3596(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1480), .Q(n89));
    nand g3597(n2466 ,n2148 ,n1921);
    dff g3598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2578), .Q(n36[0]));
    nand g3599(n60 ,n6[11] ,n57);
    dff g3600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2397), .Q(n22[4]));
    nor g3601(n2619 ,n3573 ,n2598);
    dff g3602(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2141), .Q(n25[7]));
    nand g3603(n1758 ,n8[29] ,n537);
    nand g3604(n1267 ,n6[15] ,n531);
    not g3605(n718 ,n717);
    nand g3606(n2451 ,n2173 ,n1936);
    nor g3607(n715 ,n26[2] ,n6[5]);
    dff g3608(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2561), .Q(n21[0]));
    nand g3609(n3127 ,n1566 ,n2972);
    nand g3610(n1558 ,n30[15] ,n1150);
    nand g3611(n2912 ,n27[10] ,n2694);
    not g3612(n373 ,n3432);
    dff g3613(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2157), .Q(n25[4]));
    nand g3614(n1101 ,n31[14] ,n527);
    nor g3615(n2630 ,n838 ,n2608);
    nand g3616(n720 ,n33[1] ,n574);
    xnor g3617(n3525 ,n190 ,n24[9]);
    nand g3618(n504 ,n450 ,n503);
    nand g3619(n2795 ,n10[10] ,n2690);
    nand g3620(n3014 ,n9[2] ,n2848);
    nand g3621(n918 ,n650 ,n725);
    not g3622(n261 ,n260);
    nand g3623(n1186 ,n25[3] ,n1032);
    nand g3624(n1677 ,n8[9] ,n531);
    nand g3625(n1663 ,n3494 ,n531);
    not g3626(n2649 ,n2640);
    nand g3627(n1400 ,n32[9] ,n1149);
    dff g3628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3202), .Q(n9[11]));
    xnor g3629(n3450 ,n330 ,n21[22]);
    nand g3630(n1595 ,n3474 ,n531);
    nand g3631(n3224 ,n24[14] ,n3219);
    nand g3632(n1653 ,n3557 ,n533);
    dff g3633(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2412), .Q(n23[22]));
    nand g3634(n1426 ,n25[30] ,n1147);
    nand g3635(n1110 ,n31[23] ,n527);
    nor g3636(n506 ,n391 ,n505);
    nand g3637(n2203 ,n32[5] ,n523);
    nor g3638(n667 ,n564 ,n30[9]);
    nor g3639(n617 ,n538 ,n28[14]);
    xor g3640(n865 ,n6[17] ,n31[11]);
    nand g3641(n2862 ,n25[2] ,n2696);
    nand g3642(n1570 ,n30[9] ,n1150);
    nand g3643(n2688 ,n7[7] ,n2642);
    dff g3644(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3058), .Q(n9[5]));
    nand g3645(n3325 ,n3221 ,n22[16]);
    nand g3646(n2264 ,n21[18] ,n1951);
    nor g3647(n2663 ,n2615 ,n2647);
    nand g3648(n1842 ,n22[4] ,n1464);
    nand g3649(n3125 ,n1560 ,n2969);
    not g3650(n2753 ,n2736);
    nand g3651(n1494 ,n8[1] ,n530);
    nand g3652(n2030 ,n1381 ,n1296);
    nand g3653(n805 ,n26[11] ,n538);
    nor g3654(n3083 ,n2867 ,n3017);
    nand g3655(n1982 ,n1341 ,n1492);
    nand g3656(n1294 ,n6[30] ,n531);
    nor g3657(n695 ,n540 ,n31[0]);
    xnor g3658(n3544 ,n154 ,n23[21]);
    buf g3659(n18[4], 1'b0);
    nor g3660(n2617 ,n3572 ,n2598);
    dff g3661(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2354), .Q(n26[17]));
    nand g3662(n2757 ,n942 ,n2692);
    not g3663(n2743 ,n2710);
    or g3664(n658 ,n560 ,n31[3]);
    nand g3665(n1888 ,n23[23] ,n1465);
    xnor g3666(n3498 ,n240 ,n22[5]);
    nand g3667(n2729 ,n11[11] ,n2641);
    nand g3668(n2713 ,n11[27] ,n2641);
    nand g3669(n2816 ,n25[27] ,n2696);
    nand g3670(n2357 ,n2093 ,n1772);
    not g3671(n372 ,n3385);
    dff g3672(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2129), .Q(n25[15]));
    not g3673(n311 ,n310);
    not g3674(n3222 ,n6[5]);
    nand g3675(n1533 ,n1129 ,n1127);
    or g3676(n668 ,n546 ,n29[16]);
    nand g3677(n2353 ,n2085 ,n1769);
    nand g3678(n2907 ,n27[7] ,n2694);
    xnor g3679(n3452 ,n326 ,n21[20]);
    nand g3680(n761 ,n33[0] ,n574);
    dff g3681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1952), .Q(n27[30]));
    nand g3682(n2344 ,n2046 ,n1712);
    dff g3683(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3116), .Q(n10[2]));
    dff g3684(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2518), .Q(n24[12]));
    nand g3685(n3143 ,n2903 ,n3014);
    nand g3686(n976 ,n681 ,n752);
    buf g3687(n18[7], 1'b0);
    not g3688(n241 ,n240);
    nand g3689(n3226 ,n23[20] ,n3219);
    nand g3690(n1772 ,n8[15] ,n536);
    nand g3691(n1344 ,n29[5] ,n1147);
    nand g3692(n3184 ,n2991 ,n3056);
    nand g3693(n960 ,n737 ,n789);
    nand g3694(n752 ,n31[4] ,n552);
    nor g3695(n3074 ,n2847 ,n3032);
    nand g3696(n2062 ,n1389 ,n1557);
    dff g3697(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2241), .Q(n23[0]));
    nand g3698(n1580 ,n8[31] ,n530);
    nand g3699(n1874 ,n3528 ,n537);
    dff g3700(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3108), .Q(n10[11]));
    nand g3701(n2167 ,n1469 ,n1684);
    dff g3702(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2396), .Q(n22[5]));
    nor g3703(n1151 ,n37[0] ,n1062);
    nand g3704(n994 ,n821 ,n771);
    not g3705(n87 ,n86);
    nand g3706(n1921 ,n8[23] ,n535);
    nand g3707(n2968 ,n6[21] ,n2849);
    nand g3708(n2177 ,n32[23] ,n1462);
    nand g3709(n1353 ,n32[24] ,n1149);
    nand g3710(n95 ,n34[1] ,n34[0]);
    nand g3711(n2893 ,n1232 ,n2688);
    nand g3712(n1117 ,n995 ,n1033);
    nand g3713(n194 ,n24[10] ,n193);
    nand g3714(n2967 ,n6[22] ,n2849);
    nand g3715(n1486 ,n8[27] ,n531);
    dff g3716(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n836), .Q(n20[10]));
    nand g3717(n3131 ,n2571 ,n3002);
    nand g3718(n787 ,n30[17] ,n549);
    nand g3719(n427 ,n3382 ,n349);
    not g3720(n231 ,n230);
    nand g3721(n2174 ,n32[25] ,n523);
    nand g3722(n1778 ,n3444 ,n535);
    nand g3723(n1219 ,n25[15] ,n529);
    nand g3724(n3171 ,n2823 ,n3065);
    nand g3725(n2058 ,n1382 ,n1449);
    nand g3726(n1202 ,n27[19] ,n1031);
    nand g3727(n1701 ,n6[22] ,n536);
    nand g3728(n1319 ,n31[18] ,n522);
    not g3729(n851 ,n850);
    nand g3730(n1672 ,n8[12] ,n532);
    not g3731(n40 ,n6[24]);
    nand g3732(n3289 ,n3220 ,n21[14]);
    nand g3733(n3179 ,n2863 ,n3085);
    dff g3734(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2007), .Q(n27[11]));
    nand g3735(n1169 ,n31[5] ,n1031);
    nand g3736(n3026 ,n2740 ,n2830);
    nand g3737(n2065 ,n1393 ,n1392);
    nand g3738(n1745 ,n6[11] ,n535);
    nand g3739(n1273 ,n6[9] ,n531);
    nor g3740(n1049 ,n873 ,n947);
    dff g3741(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2426), .Q(n32[8]));
    not g3742(n2208 ,n2045);
    nor g3743(n2964 ,n556 ,n2850);
    nand g3744(n3142 ,n2902 ,n3013);
    nand g3745(n3423 ,n3317 ,n3251);
    nor g3746(n2933 ,n1503 ,n2876);
    nand g3747(n1265 ,n6[17] ,n531);
    dff g3748(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2151), .Q(n25[5]));
    not g3749(n367 ,n3377);
    nor g3750(n2944 ,n1516 ,n2887);
    nand g3751(n190 ,n24[8] ,n189);
    nand g3752(n1592 ,n3490 ,n531);
    nor g3753(n2957 ,n1538 ,n2900);
    not g3754(n39 ,n6[16]);
    nor g3755(n841 ,n588 ,n539);
    nor g3756(n413 ,n381 ,n3393);
    nand g3757(n2478 ,n1661 ,n1909);
    nand g3758(n2297 ,n24[17] ,n1950);
    nand g3759(n1165 ,n31[7] ,n1031);
    or g3760(n409 ,n375 ,n3427);
    dff g3761(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1947), .Q(n27[31]));
    nand g3762(n2499 ,n1849 ,n2284);
    not g3763(n378 ,n3419);
    nand g3764(n2415 ,n1084 ,n1920);
    dff g3765(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2402), .Q(n26[0]));
    dff g3766(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2359), .Q(n26[12]));
    nand g3767(n1196 ,n29[7] ,n529);
    or g3768(n625 ,n544 ,n30[5]);
    not g3769(n2642 ,n2643);
    nand g3770(n2199 ,n32[7] ,n523);
    or g3771(n2580 ,n895 ,n2564);
    dff g3772(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2448), .Q(n28[8]));
    not g3773(n209 ,n208);
    nand g3774(n1952 ,n1309 ,n1483);
    nand g3775(n1873 ,n3527 ,n536);
    or g3776(n931 ,n620 ,n592);
    nand g3777(n88 ,n6[30] ,n87);
    dff g3778(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2382), .Q(n26[4]));
    xnor g3779(n3500 ,n236 ,n22[3]);
    not g3780(n145 ,n144);
    xnor g3781(n3511 ,n216 ,n24[23]);
    nand g3782(n1572 ,n30[8] ,n1150);
    nand g3783(n3303 ,n3221 ,n22[21]);
    nand g3784(n516 ,n453 ,n515);
    dff g3785(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2463), .Q(n28[20]));
    nor g3786(n670 ,n540 ,n30[0]);
    or g3787(n1307 ,n1063 ,n1094);
    dff g3788(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2147), .Q(n25[6]));
    nand g3789(n1805 ,n3470 ,n534);
    nand g3790(n2206 ,n32[2] ,n523);
    not g3791(n73 ,n72);
    dff g3792(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2034), .Q(n29[8]));
    dff g3793(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2451), .Q(n28[9]));
    nand g3794(n2441 ,n2184 ,n1732);
    nand g3795(n1469 ,n25[2] ,n1147);
    nand g3796(n1237 ,n25[13] ,n529);
    nor g3797(n3161 ,n2229 ,n3134);
    dff g3798(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2324), .Q(n30[15]));
    nand g3799(n2997 ,n9[18] ,n2848);
    nand g3800(n2706 ,n2618 ,n2629);
    nand g3801(n449 ,n3435 ,n366);
    nand g3802(n1116 ,n1002 ,n1033);
    nand g3803(n3260 ,n23[24] ,n3219);
    nor g3804(n2938 ,n1510 ,n2881);
    nand g3805(n3035 ,n2728 ,n2921);
    dff g3806(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2506), .Q(n24[23]));
    nor g3807(n2955 ,n1535 ,n2898);
    nand g3808(n1459 ,n25[5] ,n521);
    nand g3809(n1113 ,n25[29] ,n529);
    nand g3810(n1496 ,n8[10] ,n530);
    nor g3811(n1053 ,n885 ,n969);
    nand g3812(n1252 ,n1044 ,n1083);
    nand g3813(n1650 ,n8[22] ,n533);
    xnor g3814(n3467 ,n298 ,n21[5]);
    nand g3815(n2723 ,n11[17] ,n2641);
    nand g3816(n2385 ,n1593 ,n1826);
    nand g3817(n2185 ,n32[17] ,n523);
    nand g3818(n1291 ,n6[20] ,n531);
    nand g3819(n2248 ,n1687 ,n2214);
    not g3820(n579 ,n25[15]);
    nor g3821(n892 ,n700 ,n684);
    nand g3822(n1790 ,n3455 ,n534);
    nand g3823(n1746 ,n6[10] ,n535);
    nand g3824(n2256 ,n21[26] ,n1951);
    nand g3825(n1607 ,n3487 ,n531);
    xnor g3826(n3527 ,n186 ,n24[7]);
    xnor g3827(n3535 ,n172 ,n23[30]);
    nand g3828(n109 ,n35[2] ,n108);
    nand g3829(n2545 ,n1787 ,n2262);
    nand g3830(n2251 ,n21[31] ,n1951);
    dff g3831(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2431), .Q(n32[11]));
    nand g3832(n2548 ,n1783 ,n2259);
    nand g3833(n1686 ,n8[0] ,n533);
    nor g3834(n2847 ,n579 ,n2695);
    nand g3835(n1557 ,n30[16] ,n1150);
    nor g3836(n604 ,n26[12] ,n6[5]);
    nand g3837(n2682 ,n7[30] ,n2642);
    nand g3838(n3379 ,n3326 ,n3264);
    xnor g3839(n884 ,n6[31] ,n32[25]);
    nand g3840(n79 ,n6[21] ,n75);
    nand g3841(n3415 ,n3318 ,n3283);
    nand g3842(n3212 ,n2993 ,n3151);
    nand g3843(n2205 ,n32[3] ,n523);
    nand g3844(n743 ,n29[19] ,n556);
    or g3845(n1091 ,n960 ,n1014);
    dff g3846(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2376), .Q(n26[5]));
    nor g3847(n501 ,n443 ,n500);
    nand g3848(n3170 ,n2818 ,n3063);
    not g3849(n566 ,n37[0]);
    nor g3850(n52 ,n39 ,n48);
    nand g3851(n2402 ,n2110 ,n1848);
    xor g3852(n3547 ,n23[18] ,n148);
    xnor g3853(n3457 ,n318 ,n21[15]);
    nand g3854(n1882 ,n23[29] ,n1465);
    nand g3855(n3304 ,n3221 ,n21[21]);
    nand g3856(n3380 ,n3328 ,n3267);
    nor g3857(n880 ,n663 ,n643);
    nand g3858(n3214 ,n2984 ,n3148);
    nand g3859(n1441 ,n25[15] ,n521);
    nand g3860(n3109 ,n2795 ,n2949);
    nand g3861(n2418 ,n2206 ,n1748);
    nand g3862(n2880 ,n1116 ,n2674);
    nand g3863(n2669 ,n7[25] ,n2642);
    nor g3864(n2615 ,n3577 ,n2598);
    nand g3865(n1060 ,n91 ,n950);
    dff g3866(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2480), .Q(n23[4]));
    nand g3867(n1381 ,n29[11] ,n1147);
    nand g3868(n2856 ,n27[5] ,n2694);
    nand g3869(n1671 ,n8[13] ,n533);
    nand g3870(n1087 ,n1024 ,n1019);
    nand g3871(n164 ,n23[25] ,n163);
    nand g3872(n1331 ,n27[24] ,n522);
    dff g3873(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2004), .Q(n27[13]));
    nand g3874(n1669 ,n8[15] ,n530);
    nand g3875(n2789 ,n10[16] ,n2690);
    nand g3876(n1129 ,n27[4] ,n527);
    dff g3877(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2018), .Q(n27[7]));
    not g3878(n299 ,n298);
    not g3879(n335 ,n334);
    dff g3880(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2501), .Q(n24[29]));
    dff g3881(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2019), .Q(n29[19]));
    nand g3882(n1965 ,n1325 ,n1263);
    nand g3883(n3324 ,n3221 ,n22[0]);
    nor g3884(n1047 ,n878 ,n957);
    dff g3885(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2318), .Q(n30[24]));
    nand g3886(n1430 ,n25[25] ,n1147);
    nand g3887(n2710 ,n11[30] ,n2641);
    nand g3888(n1568 ,n30[10] ,n1150);
    nand g3889(n1742 ,n6[14] ,n535);
    nand g3890(n286 ,n22[28] ,n285);
    xnor g3891(n3528 ,n184 ,n24[6]);
    xnor g3892(n3503 ,n232 ,n24[31]);
    dff g3893(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2379), .Q(n22[19]));
    nor g3894(n432 ,n380 ,n3413);
    nand g3895(n3208 ,n2999 ,n3156);
    nand g3896(n2820 ,n27[25] ,n2694);
    nor g3897(n601 ,n2 ,n3);
    nor g3898(n399 ,n374 ,n3392);
    nand g3899(n1800 ,n3464 ,n534);
    dff g3900(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2653), .Q(n34[5]));
    xnor g3901(n3367 ,n6[22] ,n79);
    xnor g3902(n3489 ,n258 ,n22[14]);
    nand g3903(n1511 ,n1195 ,n1069);
    nand g3904(n1552 ,n1218 ,n1208);
    nand g3905(n969 ,n750 ,n709);
    nor g3906(n2932 ,n1502 ,n2875);
    nand g3907(n2716 ,n11[24] ,n2641);
    or g3908(n882 ,n677 ,n660);
    dff g3909(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2659), .Q(n35[6]));
    nand g3910(n1972 ,n1331 ,n1489);
    nand g3911(n737 ,n29[7] ,n561);
    xnor g3912(n3369 ,n6[24] ,n81);
    nand g3913(n2303 ,n24[11] ,n1950);
    nand g3914(n979 ,n676 ,n733);
    nand g3915(n1600 ,n3479 ,n531);
    nand g3916(n2194 ,n32[11] ,n523);
    nand g3917(n3234 ,n23[29] ,n3222);
    or g3918(n636 ,n558 ,n29[8]);
    nand g3919(n2715 ,n11[25] ,n2641);
    nand g3920(n1440 ,n25[16] ,n521);
    nand g3921(n2853 ,n27[6] ,n2694);
    nand g3922(n1631 ,n3538 ,n532);
    nand g3923(n3255 ,n24[5] ,n3222);
    dff g3924(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3210), .Q(n9[20]));
    nor g3925(n3081 ,n2752 ,n3042);
    nand g3926(n158 ,n23[22] ,n157);
    nand g3927(n828 ,n33[0] ,n1);
    nand g3928(n1962 ,n1322 ,n1262);
    nand g3929(n1327 ,n31[12] ,n1146);
    nand g3930(n2071 ,n26[23] ,n1463);
    dff g3931(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2320), .Q(n30[19]));
    nand g3932(n1343 ,n32[6] ,n1149);
    dff g3933(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1479), .Q(n91));
    nand g3934(n2363 ,n2104 ,n1809);
    nand g3935(n1174 ,n31[3] ,n527);
    nand g3936(n1491 ,n8[22] ,n530);
    nand g3937(n1320 ,n31[17] ,n522);
    nand g3938(n1845 ,n22[1] ,n1464);
    dff g3939(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3212), .Q(n9[22]));
    nand g3940(n951 ,n5 ,n829);
    nor g3941(n2584 ,n2583 ,n2234);
    nor g3942(n660 ,n553 ,n31[23]);
    nand g3943(n1378 ,n32[20] ,n1149);
    nor g3944(n3056 ,n2573 ,n2965);
    nand g3945(n2060 ,n1385 ,n1384);
    nand g3946(n3314 ,n3220 ,n22[27]);
    nand g3947(n2471 ,n2142 ,n1916);
    nand g3948(n3438 ,n3302 ,n3234);
    nor g3949(n2604 ,n3568 ,n2600);
    nand g3950(n2244 ,n1376 ,n2210);
    not g3951(n179 ,n178);
    or g3952(n693 ,n558 ,n32[8]);
    nand g3953(n1893 ,n23[18] ,n1465);
    nand g3954(n1726 ,n6[30] ,n534);
    nand g3955(n2164 ,n28[15] ,n523);
    nand g3956(n1931 ,n8[14] ,n535);
    nand g3957(n1698 ,n6[6] ,n534);
    nand g3958(n2468 ,n1992 ,n1701);
    nand g3959(n770 ,n32[20] ,n557);
    nand g3960(n1928 ,n8[17] ,n535);
    nor g3961(n2627 ,n836 ,n2608);
    nand g3962(n1997 ,n1415 ,n1505);
    nand g3963(n2684 ,n7[11] ,n2642);
    nand g3964(n1853 ,n3508 ,n537);
    nand g3965(n2266 ,n21[16] ,n1951);
    dff g3966(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2399), .Q(n26[1]));
    nand g3967(n2445 ,n2178 ,n1728);
    nand g3968(n291 ,n21[1] ,n21[0]);
    nor g3969(n2838 ,n568 ,n2695);
    nand g3970(n1274 ,n6[8] ,n530);
    not g3971(n369 ,n3439);
    nand g3972(n990 ,n675 ,n788);
    nand g3973(n1477 ,n27[7] ,n1146);
    nor g3974(n113 ,n35[5] ,n112);
    xnor g3975(n900 ,n6[25] ,n30[19]);
    nor g3976(n928 ,n623 ,n715);
    nor g3977(n2954 ,n1534 ,n2897);
    nand g3978(n1780 ,n3446 ,n535);
    nand g3979(n1499 ,n1121 ,n1214);
    buf g3980(n18[2], 1'b0);
    nand g3981(n3408 ,n3322 ,n3259);
    nand g3982(n1550 ,n30[19] ,n1150);
    nand g3983(n2498 ,n1847 ,n2283);
    nor g3984(n1010 ,n988 ,n958);
    nand g3985(n3335 ,n3221 ,n22[1]);
    nor g3986(n1148 ,n716 ,n1036);
    nor g3987(n3155 ,n2223 ,n3127);
    nor g3988(n2976 ,n561 ,n2850);
    nand g3989(n1843 ,n22[3] ,n1464);
    dff g3990(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2471), .Q(n28[27]));
    nand g3991(n731 ,n29[20] ,n557);
    not g3992(n530 ,n522);
    nand g3993(n3215 ,n2974 ,n3157);
    nand g3994(n2988 ,n9[27] ,n2848);
    nor g3995(n2606 ,n3570 ,n2600);
    nand g3996(n2104 ,n26[6] ,n520);
    not g3997(n159 ,n158);
    nand g3998(n3271 ,n24[6] ,n3222);
    nand g3999(n1714 ,n6[11] ,n536);
    nor g4000(n1026 ,n869 ,n983);
    dff g4001(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2529), .Q(n21[4]));
    nand g4002(n138 ,n23[11] ,n137);
    nand g4003(n914 ,n627 ,n804);
    not g4004(n534 ,n523);
    dff g4005(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2361), .Q(n26[10]));
    nand g4006(n3428 ,n3288 ,n3285);
    nor g4007(n926 ,n33[1] ,n719);
    not g4008(n2599 ,n2600);
    nand g4009(n859 ,n35[5] ,n1);
    nor g4010(n3065 ,n2747 ,n3023);
    nand g4011(n1233 ,n29[13] ,n529);
    nor g4012(n620 ,n538 ,n28[10]);
    nand g4013(n1876 ,n3530 ,n536);
    nand g4014(n2115 ,n1429 ,n1625);
    nand g4015(n804 ,n32[23] ,n553);
    nand g4016(n3201 ,n2853 ,n3051);
    nand g4017(n2731 ,n11[9] ,n2641);
    xnor g4018(n3495 ,n246 ,n22[8]);
    nand g4019(n772 ,n26[21] ,n538);
    dff g4020(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2514), .Q(n24[15]));
    nand g4021(n2924 ,n27[15] ,n2694);
    dff g4022(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3178), .Q(n11[2]));
    nor g4023(n639 ,n547 ,n31[10]);
    nor g4024(n2806 ,n569 ,n2695);
    nand g4025(n1369 ,n3375 ,n1148);
    nand g4026(n1316 ,n27[28] ,n1146);
    nand g4027(n2002 ,n30[6] ,n520);
    nand g4028(n2270 ,n21[12] ,n1951);
    nand g4029(n2299 ,n24[15] ,n1950);
    nand g4030(n3337 ,n3221 ,n21[7]);
    not g4031(n847 ,n846);
    nand g4032(n1990 ,n30[18] ,n1463);
    nand g4033(n3393 ,n3292 ,n3229);
    xnor g4034(n3560 ,n124 ,n23[5]);
    nand g4035(n3377 ,n3323 ,n3280);
    dff g4036(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2127), .Q(n25[17]));
    not g4037(n363 ,n3386);
    nand g4038(n1856 ,n3511 ,n537);
    nand g4039(n2414 ,n1638 ,n1891);
    nor g4040(n472 ,n396 ,n467);
    nand g4041(n1458 ,n25[6] ,n1147);
    nand g4042(n1449 ,n3369 ,n1148);
    xnor g4043(n3569 ,n34[3] ,n97);
    nand g4044(n1846 ,n22[0] ,n1464);
    dff g4045(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2032), .Q(n29[9]));
    nand g4046(n3384 ,n3337 ,n3274);
    not g4047(n98 ,n97);
    nor g4048(n2930 ,n1500 ,n2873);
    nand g4049(n2294 ,n24[20] ,n1950);
    nand g4050(n130 ,n23[7] ,n129);
    nand g4051(n1374 ,n32[22] ,n1149);
    dff g4052(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2428), .Q(n32[9]));
    nand g4053(n842 ,n34[0] ,n1);
    nand g4054(n3282 ,n24[11] ,n3219);
    nand g4055(n2031 ,n1348 ,n1285);
    not g4056(n127 ,n126);
    nand g4057(n2852 ,n25[6] ,n2696);
endmodule
