module top (n0, n1, n2, n3, n4, n5, n6);
    input n0, n1;
    input [13:0] n2;
    input [12:0] n3;
    output [12:0] n4, n5, n6;
    wire n0, n1;
    wire [13:0] n2;
    wire [12:0] n3;
    wire [12:0] n4, n5, n6;
    wire [12:0] n7;
    wire [12:0] n8;
    wire [12:0] n9;
    wire [12:0] n10;
    wire [12:0] n11;
    wire [12:0] n12;
    wire [2:0] n13;
    wire [3:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695;
    xnor g0(n141 ,n2[2] ,n3[2]);
    xnor g1(n37 ,n659 ,n12[7]);
    xnor g2(n130 ,n2[11] ,n3[11]);
    dff g3(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n436), .Q(n13[2]));
    nand g4(n321 ,n267 ,n300);
    nand g5(n51 ,n19 ,n50);
    nor g6(n117 ,n2[8] ,n3[8]);
    nand g7(n306 ,n11[2] ,n285);
    xnor g8(n92 ,n636 ,n12[11]);
    xnor g9(n5[11] ,n570 ,n7[11]);
    not g10(n673 ,n672);
    not g11(n668 ,n3[8]);
    xnor g12(n644 ,n30 ,n53);
    xor g13(n577 ,n563 ,n10[5]);
    nand g14(n473 ,n439 ,n407);
    nand g15(n464 ,n7[7] ,n329);
    nor g16(n296 ,n1 ,n283);
    nor g17(n343 ,n262 ,n313);
    nand g18(n540 ,n513 ,n536);
    xnor g19(n5[0] ,n565 ,n7[0]);
    not g20(n252 ,n639);
    nor g21(n380 ,n233 ,n295);
    dff g22(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n505), .Q(n9[4]));
    not g23(n287 ,n286);
    xor g24(n607 ,n608 ,n10[9]);
    nand g25(n440 ,n8[0] ,n334);
    nor g26(n362 ,n241 ,n295);
    nand g27(n480 ,n452 ,n416);
    nor g28(n325 ,n231 ,n295);
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n545), .Q(n11[5]));
    xnor g30(n4[11] ,n570 ,n8[11]);
    xnor g31(n5[5] ,n577 ,n7[5]);
    xor g32(n657 ,n2[5] ,n10[5]);
    not g33(n233 ,n626);
    nor g34(n326 ,n252 ,n295);
    nand g35(n20 ,n662 ,n12[10]);
    xor g36(n593 ,n594 ,n10[2]);
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n541), .Q(n11[10]));
    xnor g38(n612 ,n130 ,n165);
    xnor g39(n604 ,n139 ,n157);
    not g40(n246 ,n620);
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n467), .Q(n7[5]));
    nor g42(n297 ,n1 ,n293);
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n479), .Q(n9[10]));
    nor g44(n164 ,n134 ,n163);
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n499), .Q(n9[2]));
    nand g46(n60 ,n28 ,n59);
    nand g47(n496 ,n465 ,n430);
    nand g48(n490 ,n460 ,n424);
    nand g49(n431 ,n7[5] ,n336);
    nand g50(n554 ,n11[6] ,n12[6]);
    nor g51(n102 ,n68 ,n101);
    xor g52(n568 ,n557 ,n10[7]);
    xnor g53(n5[12] ,n566 ,n7[12]);
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n485), .Q(n9[6]));
    nor g55(n384 ,n232 ,n295);
    nand g56(n485 ,n451 ,n417);
    xnor g57(n179 ,n613 ,n12[11]);
    nor g58(n374 ,n229 ,n295);
    not g59(n140 ,n139);
    xor g60(n613 ,n614 ,n10[12]);
    nand g61(n491 ,n461 ,n425);
    nand g62(n541 ,n509 ,n525);
    nand g63(n318 ,n270 ,n306);
    not g64(n229 ,n585);
    nand g65(n494 ,n463 ,n408);
    nand g66(n74 ,n635 ,n12[10]);
    nand g67(n457 ,n9[0] ,n334);
    nand g68(n171 ,n599 ,n12[4]);
    xor g69(n634 ,n3[8] ,n10[8]);
    nand g70(n506 ,n464 ,n428);
    nand g71(n691 ,n2[13] ,n2[12]);
    xnor g72(n625 ,n95 ,n114);
    nor g73(n371 ,n224 ,n295);
    xor g74(n596 ,n143 ,n148);
    not g75(n80 ,n79);
    nand g76(n77 ,n631 ,n12[6]);
    nor g77(n151 ,n124 ,n150);
    xnor g78(n10[7] ,n3[7] ,n679);
    nand g79(n558 ,n11[2] ,n12[2]);
    xnor g80(n6[10] ,n571 ,n9[10]);
    nor g81(n521 ,n14[0] ,n466);
    nand g82(n66 ,n42 ,n65);
    nand g83(n686 ,n3[10] ,n685);
    nor g84(n404 ,n356 ,n339);
    nor g85(n353 ,n250 ,n295);
    not g86(n87 ,n86);
    nand g87(n486 ,n442 ,n409);
    xnor g88(n131 ,n2[4] ,n3[4]);
    xnor g89(n10[8] ,n3[8] ,n681);
    nand g90(n406 ,n365 ,n351);
    xnor g91(n43 ,n655 ,n12[3]);
    nor g92(n119 ,n2[9] ,n3[9]);
    nand g93(n320 ,n265 ,n306);
    nand g94(n322 ,n615 ,n296);
    xor g95(n581 ,n196 ,n200);
    xnor g96(n6[7] ,n568 ,n9[7]);
    not g97(n181 ,n180);
    nand g98(n471 ,n435 ,n403);
    xnor g99(n589 ,n180 ,n216);
    not g100(n259 ,n11[10]);
    nand g101(n443 ,n9[12] ,n338);
    xnor g102(n587 ,n182 ,n212);
    nand g103(n498 ,n322 ,n393);
    nor g104(n299 ,n1 ,n292);
    nor g105(n17 ,n657 ,n12[5]);
    not g106(n225 ,n646);
    xnor g107(n143 ,n2[3] ,n3[3]);
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n500), .Q(n8[1]));
    xor g109(n654 ,n2[2] ,n10[2]);
    nor g110(n386 ,n236 ,n295);
    xor g111(n567 ,n556 ,n10[1]);
    nand g112(n463 ,n7[8] ,n349);
    nand g113(n205 ,n185 ,n204);
    not g114(n295 ,n296);
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n489), .Q(n7[12]));
    xor g116(n605 ,n606 ,n10[8]);
    xor g117(n597 ,n598 ,n10[4]);
    xnor g118(n95 ,n637 ,n10[11]);
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n473), .Q(n8[10]));
    nand g120(n688 ,n3[11] ,n687);
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n538), .Q(n14[0]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n471), .Q(n8[12]));
    xnor g123(n133 ,n2[5] ,n3[5]);
    xnor g124(n10[6] ,n3[6] ,n677);
    not g125(n234 ,n619);
    nand g126(n489 ,n459 ,n423);
    nand g127(n301 ,n284 ,n289);
    xnor g128(n82 ,n631 ,n12[6]);
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n501), .Q(n9[1]));
    xor g130(n662 ,n2[10] ,n10[10]);
    nor g131(n419 ,n354 ,n335);
    xor g132(n626 ,n638 ,n116);
    nor g133(n382 ,n245 ,n295);
    nor g134(n420 ,n373 ,n335);
    not g135(n221 ,n582);
    xor g136(n601 ,n602 ,n10[6]);
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n474), .Q(n8[9]));
    not g138(n251 ,n618);
    not g139(n237 ,n650);
    nor g140(n123 ,n2[10] ,n3[10]);
    not g141(n91 ,n90);
    nor g142(n387 ,n246 ,n295);
    not g143(n231 ,n617);
    or g144(n201 ,n196 ,n200);
    xor g145(n591 ,n592 ,n10[1]);
    nor g146(n421 ,n375 ,n330);
    nor g147(n413 ,n368 ,n343);
    nor g148(n162 ,n132 ,n161);
    xnor g149(n4[6] ,n575 ,n8[6]);
    nand g150(n47 ,n16 ,n46);
    nand g151(n694 ,n1 ,n693);
    nand g152(n211 ,n198 ,n210);
    not g153(n236 ,n621);
    xnor g154(n6[3] ,n572 ,n9[3]);
    nand g155(n305 ,n10[12] ,n285);
    nand g156(n345 ,n284 ,n314);
    xnor g157(n5[8] ,n573 ,n7[8]);
    nand g158(n58 ,n38 ,n57);
    nand g159(n98 ,n69 ,n97);
    xor g160(n653 ,n2[1] ,n10[1]);
    nand g161(n338 ,n284 ,n305);
    nand g162(n492 ,n440 ,n402);
    nand g163(n499 ,n378 ,n394);
    not g164(n240 ,n645);
    nor g165(n358 ,n248 ,n295);
    xnor g166(n586 ,n197 ,n210);
    nand g167(n207 ,n191 ,n206);
    xor g168(n632 ,n3[6] ,n10[6]);
    nand g169(n355 ,n13[1] ,n299);
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n486), .Q(n8[8]));
    nor g171(n120 ,n2[11] ,n3[11]);
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n470), .Q(n7[0]));
    xnor g173(n6[1] ,n567 ,n9[1]);
    nand g174(n444 ,n8[7] ,n329);
    nand g175(n309 ,n10[7] ,n285);
    nand g176(n562 ,n11[4] ,n12[4]);
    nand g177(n488 ,n458 ,n422);
    xor g178(n635 ,n3[9] ,n10[9]);
    xnor g179(n6[5] ,n577 ,n9[5]);
    nand g180(n447 ,n8[6] ,n342);
    nand g181(n484 ,n450 ,n415);
    not g182(n232 ,n623);
    xnor g183(n192 ,n603 ,n12[6]);
    nand g184(n495 ,n456 ,n420);
    nand g185(n310 ,n10[4] ,n285);
    nand g186(n302 ,n284 ,n290);
    xor g187(n636 ,n3[10] ,n10[10]);
    nor g188(n381 ,n243 ,n295);
    xnor g189(n196 ,n595 ,n12[2]);
    nor g190(n407 ,n358 ,n340);
    xnor g191(n10[3] ,n3[3] ,n672);
    or g192(n12[10] ,n10[11] ,n10[9]);
    nand g193(n204 ,n170 ,n203);
    nand g194(n156 ,n138 ,n155);
    xnor g195(n606 ,n159 ,n144);
    xnor g196(n4[8] ,n573 ,n8[8]);
    nand g197(n551 ,n517 ,n534);
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n477), .Q(n9[12]));
    xor g199(n609 ,n610 ,n10[10]);
    nor g200(n294 ,n11[12] ,n291);
    nor g201(n166 ,n130 ,n165);
    xnor g202(n5[7] ,n568 ,n7[7]);
    xnor g203(n197 ,n605 ,n12[7]);
    nand g204(n561 ,n11[8] ,n12[8]);
    nor g205(n348 ,n255 ,n308);
    xor g206(n655 ,n2[3] ,n10[3]);
    xnor g207(n619 ,n82 ,n102);
    nand g208(n524 ,n11[7] ,n520);
    nand g209(n546 ,n515 ,n532);
    nor g210(n369 ,n235 ,n295);
    not g211(n183 ,n182);
    nand g212(n114 ,n71 ,n113);
    nand g213(n316 ,n269 ,n306);
    nand g214(n557 ,n11[7] ,n12[7]);
    nor g215(n409 ,n363 ,n348);
    nand g216(n545 ,n514 ,n531);
    nand g217(n217 ,n181 ,n216);
    nand g218(n493 ,n462 ,n426);
    xnor g219(n4[1] ,n567 ,n8[1]);
    xnor g220(n134 ,n2[10] ,n3[10]);
    nor g221(n153 ,n126 ,n152);
    nand g222(n433 ,n7[3] ,n332);
    not g223(n235 ,n584);
    xnor g224(n137 ,n2[6] ,n3[6]);
    nand g225(n67 ,n25 ,n66);
    nand g226(n300 ,n11[1] ,n285);
    nor g227(n408 ,n385 ,n348);
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n548), .Q(n11[3]));
    nor g229(n690 ,n2[13] ,n2[12]);
    xor g230(n633 ,n3[7] ,n10[7]);
    nand g231(n446 ,n9[10] ,n341);
    xor g232(n616 ,n88 ,n78);
    nand g233(n313 ,n10[6] ,n285);
    or g234(n12[8] ,n10[9] ,n10[7]);
    xnor g235(n33 ,n653 ,n12[1]);
    xor g236(n631 ,n3[5] ,n10[5]);
    nor g237(n410 ,n364 ,n350);
    nand g238(n206 ,n171 ,n205);
    not g239(n142 ,n141);
    nand g240(n475 ,n453 ,n418);
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n495), .Q(n8[4]));
    nand g242(n314 ,n10[9] ,n285);
    not g243(n222 ,n583);
    not g244(n38 ,n37);
    nand g245(n170 ,n597 ,n12[3]);
    nor g246(n430 ,n387 ,n343);
    not g247(n263 ,n11[7]);
    xnor g248(n4[0] ,n565 ,n8[0]);
    nand g249(n461 ,n7[10] ,n341);
    or g250(n12[6] ,n10[7] ,n10[5]);
    nand g251(n107 ,n91 ,n106);
    xnor g252(n585 ,n192 ,n208);
    nor g253(n400 ,n325 ,n330);
    nor g254(n676 ,n3[5] ,n675);
    nand g255(n435 ,n8[12] ,n338);
    xor g256(n573 ,n561 ,n10[8]);
    or g257(n12[5] ,n10[6] ,n10[4]);
    or g258(n12[7] ,n10[8] ,n10[6]);
    nand g259(n478 ,n445 ,n405);
    or g260(n121 ,n2[2] ,n3[2]);
    not g261(n228 ,n643);
    nor g262(n522 ,n287 ,n521);
    not g263(n40 ,n39);
    nor g264(n126 ,n2[4] ,n3[4]);
    not g265(n250 ,n587);
    nand g266(n513 ,n10[6] ,n487);
    xor g267(n576 ,n564 ,n10[9]);
    nand g268(n360 ,n665 ,n297);
    not g269(n138 ,n137);
    nand g270(n213 ,n183 ,n212);
    nor g271(n152 ,n131 ,n151);
    or g272(n391 ,n13[1] ,n351);
    xnor g273(n10[2] ,n3[2] ,n670);
    nand g274(n458 ,n8[3] ,n332);
    nand g275(n157 ,n125 ,n156);
    nand g276(n383 ,n641 ,n296);
    xor g277(n579 ,n10[1] ,n591);
    xnor g278(n643 ,n29 ,n51);
    nand g279(n23 ,n660 ,n12[8]);
    xor g280(n652 ,n2[0] ,n3[0]);
    nor g281(n402 ,n326 ,n333);
    xor g282(n666 ,n13[1] ,n13[0]);
    xnor g283(n5[4] ,n574 ,n7[4]);
    nand g284(n560 ,n11[3] ,n12[3]);
    xor g285(n651 ,n664 ,n67);
    nand g286(n109 ,n80 ,n108);
    not g287(n279 ,n278);
    nand g288(n503 ,n383 ,n396);
    xnor g289(n6[0] ,n565 ,n9[0]);
    xor g290(n639 ,n10[1] ,n652);
    nor g291(n689 ,n2[11] ,n2[10]);
    nand g292(n49 ,n18 ,n48);
    nor g293(n163 ,n119 ,n162);
    nor g294(n167 ,n120 ,n166);
    nor g295(n423 ,n380 ,n337);
    nand g296(n331 ,n284 ,n310);
    xor g297(n659 ,n2[7] ,n10[7]);
    nand g298(n177 ,n601 ,n12[5]);
    nand g299(n510 ,n10[9] ,n487);
    or g300(n390 ,n288 ,n317);
    nand g301(n200 ,n168 ,n199);
    dff g302(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n551), .Q(n11[2]));
    not g303(n695 ,n694);
    xnor g304(n621 ,n90 ,n106);
    nand g305(n208 ,n177 ,n207);
    xor g306(n594 ,n141 ,n146);
    xor g307(n642 ,n43 ,n49);
    nand g308(n534 ,n11[2] ,n520);
    or g309(n12[4] ,n10[5] ,n10[3]);
    nand g310(n556 ,n11[1] ,n12[1]);
    not g311(n149 ,n148);
    xnor g312(n4[2] ,n569 ,n8[2]);
    xor g313(n599 ,n600 ,n10[5]);
    nor g314(n379 ,n223 ,n295);
    nand g315(n452 ,n8[5] ,n336);
    xnor g316(n35 ,n661 ,n12[9]);
    xor g317(n627 ,n3[1] ,n10[1]);
    xor g318(n595 ,n596 ,n10[3]);
    dff g319(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n490), .Q(n7[11]));
    nor g320(n273 ,n11[10] ,n11[11]);
    xnor g321(n186 ,n597 ,n12[3]);
    nand g322(n97 ,n78 ,n89);
    nor g323(n340 ,n259 ,n304);
    xnor g324(n588 ,n188 ,n214);
    not g325(n256 ,n11[4]);
    nand g326(n514 ,n10[5] ,n487);
    or g327(n122 ,n2[1] ,n3[1]);
    nor g328(n415 ,n374 ,n350);
    xor g329(n572 ,n560 ,n10[3]);
    not g330(n224 ,n644);
    xor g331(n656 ,n2[4] ,n10[4]);
    xor g332(n615 ,n12[2] ,n627);
    nand g333(n175 ,n595 ,n12[2]);
    xnor g334(n5[2] ,n569 ,n7[2]);
    xnor g335(n180 ,n611 ,n12[10]);
    xor g336(n566 ,n552 ,n10[12]);
    not g337(n226 ,n586);
    xnor g338(n88 ,n628 ,n12[3]);
    nor g339(n424 ,n381 ,n339);
    nand g340(n59 ,n24 ,n58);
    nand g341(n547 ,n512 ,n524);
    nand g342(n544 ,n508 ,n528);
    not g343(n265 ,n8[2]);
    nand g344(n470 ,n434 ,n401);
    nor g345(n403 ,n362 ,n337);
    xor g346(n617 ,n94 ,n98);
    not g347(n45 ,n44);
    nand g348(n670 ,n3[1] ,n695);
    nor g349(n368 ,n240 ,n295);
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n498), .Q(n7[1]));
    xnor g351(n4[7] ,n568 ,n8[7]);
    not g352(n253 ,n11[12]);
    not g353(n32 ,n31);
    nand g354(n327 ,n616 ,n296);
    or g355(n12[3] ,n10[4] ,n10[2]);
    xnor g356(n10[12] ,n3[12] ,n688);
    or g357(n12[9] ,n10[10] ,n10[8]);
    nand g358(n105 ,n85 ,n104);
    nand g359(n500 ,n352 ,n397);
    nand g360(n61 ,n23 ,n60);
    nand g361(n438 ,n8[11] ,n347);
    not g362(n671 ,n670);
    xor g363(n571 ,n559 ,n10[10]);
    or g364(n69 ,n628 ,n12[3]);
    nor g365(n323 ,n234 ,n295);
    nand g366(n512 ,n10[7] ,n487);
    nand g367(n278 ,n14[1] ,n220);
    xnor g368(n282 ,n3[0] ,n578);
    nand g369(n218 ,n173 ,n217);
    nor g370(n356 ,n237 ,n295);
    nor g371(n418 ,n372 ,n346);
    dff g372(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n537), .Q(n14[1]));
    dff g373(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n481), .Q(n9[9]));
    nor g374(n344 ,n257 ,n314);
    dff g375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n468), .Q(n7[4]));
    not g376(n136 ,n135);
    xnor g377(n86 ,n635 ,n12[10]);
    nand g378(n518 ,n10[1] ,n487);
    nand g379(n392 ,n301 ,n316);
    nor g380(n361 ,n247 ,n295);
    nand g381(n56 ,n32 ,n55);
    xor g382(n663 ,n2[11] ,n10[11]);
    nand g383(n455 ,n9[3] ,n332);
    xnor g384(n41 ,n663 ,n12[11]);
    dff g385(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n469), .Q(n7[3]));
    xnor g386(n623 ,n86 ,n110);
    nand g387(n147 ,n142 ,n146);
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n546), .Q(n11[4]));
    xor g389(n660 ,n2[8] ,n10[8]);
    nand g390(n526 ,n11[9] ,n520);
    dff g391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n494), .Q(n7[8]));
    nand g392(n467 ,n431 ,n398);
    nor g393(n10[5] ,n676 ,n678);
    nand g394(n76 ,n632 ,n12[7]);
    nor g395(n150 ,n143 ,n149);
    not g396(n189 ,n188);
    nor g397(n160 ,n144 ,n159);
    xnor g398(n29 ,n656 ,n12[4]);
    nand g399(n530 ,n11[0] ,n520);
    xnor g400(n84 ,n632 ,n12[7]);
    nor g401(n285 ,n280 ,n278);
    xor g402(n592 ,n135 ,n128);
    dff g403(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n475), .Q(n9[5]));
    dff g404(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n497), .Q(n7[2]));
    nand g405(n456 ,n8[4] ,n331);
    xnor g406(n624 ,n92 ,n112);
    not g407(n248 ,n649);
    nand g408(n550 ,n519 ,n530);
    nand g409(n100 ,n70 ,n99);
    xnor g410(n144 ,n2[8] ,n3[8]);
    not g411(n254 ,n11[3]);
    nor g412(n68 ,n630 ,n12[5]);
    xnor g413(n129 ,n2[12] ,n3[12]);
    nand g414(n523 ,n11[12] ,n520);
    nand g415(n552 ,n10[11] ,n11[12]);
    not g416(n281 ,n280);
    not g417(n243 ,n625);
    nand g418(n215 ,n189 ,n214);
    not g419(n270 ,n9[2]);
    xnor g420(n6[11] ,n570 ,n9[11]);
    nand g421(n334 ,n284 ,n303);
    nand g422(n25 ,n663 ,n12[11]);
    or g423(n12[2] ,n10[3] ,n10[1]);
    not g424(n262 ,n11[6]);
    nand g425(n553 ,n10[1] ,n11[0]);
    not g426(n187 ,n186);
    not g427(n36 ,n35);
    nor g428(n429 ,n353 ,n344);
    not g429(n245 ,n624);
    nand g430(n48 ,n40 ,n47);
    nand g431(n681 ,n3[7] ,n680);
    not g432(n267 ,n8[1]);
    nand g433(n303 ,n3[0] ,n285);
    not g434(n227 ,n588);
    nand g435(n450 ,n9[7] ,n329);
    nand g436(n474 ,n441 ,n427);
    not g437(n298 ,n297);
    or g438(n16 ,n653 ,n12[1]);
    xnor g439(n614 ,n129 ,n167);
    nand g440(n288 ,n277 ,n274);
    dff g441(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n476), .Q(n8[7]));
    nor g442(n466 ,n271 ,n390);
    nor g443(n372 ,n222 ,n295);
    xnor g444(n6[8] ,n573 ,n9[8]);
    dff g445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n406), .Q(n13[0]));
    nor g446(n425 ,n382 ,n340);
    nor g447(n370 ,n226 ,n295);
    dff g448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n503), .Q(n8[2]));
    nand g449(n395 ,n302 ,n319);
    nor g450(n276 ,n11[8] ,n11[9]);
    or g451(n12[11] ,n10[12] ,n10[10]);
    nand g452(n539 ,n507 ,n523);
    nor g453(n154 ,n133 ,n153);
    nand g454(n342 ,n284 ,n313);
    nand g455(n71 ,n636 ,n12[11]);
    dff g456(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n491), .Q(n7[10]));
    nor g457(n161 ,n117 ,n160);
    nor g458(n124 ,n2[3] ,n3[3]);
    nand g459(n317 ,n273 ,n294);
    nor g460(n373 ,n228 ,n295);
    xnor g461(n190 ,n601 ,n12[5]);
    nand g462(n209 ,n193 ,n208);
    or g463(n284 ,n1 ,n281);
    xnor g464(n39 ,n654 ,n12[2]);
    xor g465(n611 ,n612 ,n10[11]);
    nand g466(n148 ,n121 ,n147);
    xnor g467(n4[3] ,n572 ,n8[3]);
    xor g468(n569 ,n558 ,n10[2]);
    nor g469(n401 ,n388 ,n333);
    nor g470(n675 ,n667 ,n674);
    xnor g471(n5[10] ,n571 ,n7[10]);
    nor g472(n53 ,n15 ,n52);
    not g473(n195 ,n194);
    nand g474(n509 ,n10[10] ,n487);
    xnor g475(n6[4] ,n574 ,n9[4]);
    nor g476(n398 ,n323 ,n346);
    or g477(n50 ,n43 ,n49);
    nand g478(n529 ,n286 ,n521);
    not g479(n680 ,n679);
    nand g480(n112 ,n74 ,n111);
    xor g481(n603 ,n604 ,n10[7]);
    not g482(n255 ,n11[8]);
    nor g483(n364 ,n225 ,n295);
    nand g484(n453 ,n9[5] ,n336);
    nand g485(n104 ,n77 ,n103);
    nand g486(n145 ,n128 ,n136);
    xnor g487(n194 ,n593 ,n12[1]);
    nand g488(n24 ,n659 ,n12[7]);
    nor g489(n339 ,n261 ,n307);
    nor g490(n118 ,n2[5] ,n3[5]);
    nor g491(n15 ,n656 ,n12[4]);
    nand g492(n319 ,n268 ,n300);
    not g493(n242 ,n589);
    nor g494(n337 ,n253 ,n305);
    xnor g495(n6[2] ,n569 ,n9[2]);
    nand g496(n22 ,n658 ,n12[6]);
    nand g497(n481 ,n448 ,n429);
    nor g498(n417 ,n369 ,n343);
    nand g499(n393 ,n302 ,n315);
    xnor g500(n4[10] ,n571 ,n8[10]);
    nand g501(n172 ,n607 ,n12[8]);
    nand g502(n528 ,n11[11] ,n520);
    not g503(n185 ,n184);
    nor g504(n367 ,n242 ,n295);
    xnor g505(n4[4] ,n574 ,n8[4]);
    dff g506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n483), .Q(n9[8]));
    nand g507(n210 ,n174 ,n209);
    dff g508(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n543), .Q(n11[8]));
    nor g509(n375 ,n230 ,n295);
    not g510(n83 ,n82);
    or g511(n168 ,n593 ,n12[1]);
    nand g512(n462 ,n7[9] ,n345);
    xor g513(n580 ,n194 ,n178);
    dff g514(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n488), .Q(n8[3]));
    xnor g515(n618 ,n81 ,n100);
    nand g516(n216 ,n176 ,n215);
    nand g517(n19 ,n655 ,n12[3]);
    nand g518(n106 ,n76 ,n105);
    xor g519(n578 ,n2[0] ,n3[0]);
    nand g520(n111 ,n87 ,n110);
    nor g521(n272 ,n11[6] ,n11[7]);
    nor g522(n366 ,n244 ,n295);
    xnor g523(n5[6] ,n575 ,n7[6]);
    nand g524(n199 ,n178 ,n195);
    not g525(n238 ,n12[1]);
    xnor g526(n5[9] ,n576 ,n7[9]);
    nor g527(n101 ,n81 ,n100);
    nand g528(n507 ,n10[12] ,n487);
    xnor g529(n582 ,n186 ,n202);
    dff g530(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n540), .Q(n11[6]));
    or g531(n12[1] ,n3[0] ,n10[2]);
    nand g532(n439 ,n8[10] ,n341);
    not g533(n230 ,n581);
    nand g534(n312 ,n10[3] ,n285);
    not g535(n28 ,n27);
    nand g536(n394 ,n301 ,n318);
    nand g537(n432 ,n7[4] ,n331);
    nand g538(n531 ,n11[5] ,n520);
    nand g539(n315 ,n266 ,n300);
    nor g540(n165 ,n123 ,n164);
    nand g541(n62 ,n36 ,n61);
    nor g542(n412 ,n376 ,n340);
    nor g543(n274 ,n11[4] ,n11[5]);
    nor g544(n487 ,n13[2] ,n391);
    nand g545(n108 ,n75 ,n107);
    nand g546(n437 ,n355 ,n357);
    nand g547(n538 ,n298 ,n529);
    xnor g548(n6[12] ,n566 ,n9[12]);
    nand g549(n549 ,n518 ,n535);
    or g550(n99 ,n94 ,n98);
    nand g551(n57 ,n22 ,n56);
    nor g552(n427 ,n361 ,n344);
    xor g553(n664 ,n10[12] ,n2[12]);
    xnor g554(n94 ,n629 ,n12[4]);
    xnor g555(n650 ,n41 ,n65);
    xnor g556(n182 ,n607 ,n12[8]);
    xnor g557(n5[3] ,n572 ,n7[3]);
    xnor g558(n6[9] ,n576 ,n9[9]);
    nand g559(n159 ,n127 ,n158);
    nand g560(n110 ,n72 ,n109);
    nor g561(n405 ,n367 ,n339);
    nor g562(n324 ,n251 ,n295);
    nand g563(n70 ,n629 ,n12[4]);
    nand g564(n674 ,n3[3] ,n673);
    nor g565(n693 ,n690 ,n692);
    nand g566(n460 ,n7[11] ,n347);
    or g567(n283 ,n14[1] ,n280);
    nand g568(n212 ,n169 ,n211);
    not g569(n85 ,n84);
    nand g570(n515 ,n10[4] ,n487);
    nor g571(n692 ,n691 ,n689);
    nand g572(n219 ,n13[1] ,n13[0]);
    nand g573(n502 ,n457 ,n389);
    nand g574(n564 ,n11[9] ,n12[9]);
    not g575(n239 ,n647);
    nand g576(n113 ,n93 ,n112);
    nand g577(n75 ,n633 ,n12[8]);
    nor g578(n277 ,n11[2] ,n11[3]);
    not g579(n193 ,n192);
    nand g580(n341 ,n284 ,n304);
    dff g581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n547), .Q(n11[7]));
    not g582(n244 ,n590);
    not g583(n268 ,n9[1]);
    not g584(n258 ,n11[0]);
    nand g585(n169 ,n605 ,n12[7]);
    or g586(n18 ,n654 ,n12[2]);
    nand g587(n459 ,n7[12] ,n338);
    nand g588(n517 ,n10[2] ,n487);
    nor g589(n376 ,n227 ,n295);
    nand g590(n542 ,n510 ,n526);
    xor g591(n658 ,n2[6] ,n10[6]);
    nand g592(n308 ,n10[8] ,n285);
    nor g593(n416 ,n371 ,n346);
    nand g594(n548 ,n516 ,n533);
    nand g595(n505 ,n454 ,n419);
    nand g596(n291 ,n272 ,n276);
    nand g597(n527 ,n11[8] ,n520);
    xnor g598(n4[9] ,n576 ,n8[9]);
    nand g599(n72 ,n634 ,n12[9]);
    nor g600(n350 ,n263 ,n309);
    xnor g601(n79 ,n634 ,n12[9]);
    xor g602(n630 ,n3[4] ,n10[4]);
    xnor g603(n27 ,n660 ,n12[8]);
    dff g604(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n504), .Q(n9[3]));
    nand g605(n26 ,n652 ,n10[1]);
    nor g606(n55 ,n17 ,n54);
    nor g607(n354 ,n221 ,n295);
    nand g608(n434 ,n7[0] ,n334);
    not g609(n266 ,n7[1]);
    xnor g610(n600 ,n133 ,n153);
    xor g611(n574 ,n562 ,n10[4]);
    xnor g612(n135 ,n2[1] ,n3[1]);
    dff g613(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n482), .Q(n8[6]));
    nor g614(n363 ,n239 ,n295);
    xor g615(n570 ,n555 ,n10[11]);
    nor g616(n292 ,n14[1] ,n275);
    nor g617(n414 ,n370 ,n348);
    xnor g618(n647 ,n27 ,n59);
    xnor g619(n44 ,n662 ,n12[10]);
    xnor g620(n10[11] ,n3[11] ,n686);
    nor g621(n669 ,n3[1] ,n695);
    xnor g622(n583 ,n184 ,n204);
    nand g623(n214 ,n172 ,n213);
    xnor g624(n188 ,n609 ,n12[9]);
    nand g625(n468 ,n432 ,n399);
    nor g626(n328 ,n282 ,n295);
    nand g627(n65 ,n20 ,n64);
    nand g628(n64 ,n45 ,n63);
    nand g629(n173 ,n611 ,n12[10]);
    not g630(n96 ,n95);
    nor g631(n426 ,n384 ,n344);
    xnor g632(n590 ,n179 ,n218);
    nor g633(n10[1] ,n671 ,n669);
    nor g634(n683 ,n3[9] ,n682);
    not g635(n261 ,n11[11]);
    xnor g636(n608 ,n132 ,n161);
    not g637(n685 ,n684);
    not g638(n198 ,n197);
    not g639(n241 ,n651);
    nand g640(n202 ,n175 ,n201);
    nand g641(n311 ,n10[5] ,n285);
    nor g642(n399 ,n324 ,n335);
    xor g643(n575 ,n554 ,n10[6]);
    dff g644(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n478), .Q(n9[11]));
    dff g645(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n522), .Q(n14[2]));
    xnor g646(n81 ,n630 ,n12[5]);
    xnor g647(n10[10] ,n3[10] ,n684);
    dff g648(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n506), .Q(n7[7]));
    not g649(n220 ,n1);
    nor g650(n388 ,n238 ,n295);
    nand g651(n559 ,n11[10] ,n12[10]);
    nand g652(n357 ,n666 ,n297);
    nor g653(n335 ,n256 ,n310);
    not g654(n89 ,n88);
    nand g655(n127 ,n2[7] ,n3[7]);
    nand g656(n146 ,n122 ,n145);
    nand g657(n116 ,n73 ,n115);
    dff g658(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n472), .Q(n8[11]));
    dff g659(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n492), .Q(n8[0]));
    nor g660(n520 ,n1 ,n487);
    nand g661(n304 ,n10[10] ,n285);
    dff g662(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n496), .Q(n7[6]));
    xor g663(n661 ,n2[9] ,n10[9]);
    nand g664(n684 ,n3[9] ,n682);
    nor g665(n428 ,n386 ,n350);
    nand g666(n332 ,n284 ,n312);
    not g667(n264 ,n14[2]);
    nand g668(n497 ,n327 ,n392);
    nand g669(n482 ,n447 ,n413);
    nand g670(n336 ,n284 ,n311);
    not g671(n257 ,n11[9]);
    nor g672(n346 ,n260 ,n311);
    xor g673(n638 ,n10[12] ,n3[12]);
    nand g674(n472 ,n438 ,n404);
    xor g675(n637 ,n3[11] ,n10[11]);
    nand g676(n128 ,n2[0] ,n3[0]);
    nand g677(n347 ,n284 ,n307);
    not g678(n191 ,n190);
    xnor g679(n30 ,n657 ,n12[5]);
    or g680(n351 ,n13[0] ,n298);
    nand g681(n448 ,n9[9] ,n345);
    nand g682(n516 ,n10[3] ,n487);
    not g683(n34 ,n33);
    xnor g684(n4[5] ,n577 ,n8[5]);
    or g685(n275 ,n14[0] ,n14[2]);
    xnor g686(n4[12] ,n566 ,n8[12]);
    nand g687(n537 ,n295 ,n529);
    nor g688(n155 ,n118 ,n154);
    xor g689(n629 ,n3[3] ,n10[3]);
    nand g690(n290 ,n10[1] ,n279);
    nand g691(n504 ,n455 ,n421);
    nand g692(n535 ,n11[1] ,n520);
    xor g693(n640 ,n33 ,n26);
    xnor g694(n139 ,n2[7] ,n3[7]);
    nor g695(n333 ,n258 ,n303);
    nand g696(n396 ,n301 ,n320);
    nand g697(n377 ,n579 ,n296);
    nand g698(n469 ,n433 ,n400);
    xnor g699(n5[1] ,n567 ,n7[1]);
    not g700(n678 ,n677);
    nand g701(n476 ,n444 ,n410);
    nand g702(n63 ,n21 ,n62);
    nand g703(n115 ,n96 ,n114);
    nand g704(n477 ,n443 ,n411);
    nand g705(n442 ,n8[8] ,n349);
    not g706(n667 ,n3[4]);
    xnor g707(n90 ,n633 ,n12[8]);
    nand g708(n441 ,n8[9] ,n345);
    nand g709(n533 ,n11[3] ,n520);
    nand g710(n174 ,n603 ,n12[6]);
    nand g711(n125 ,n2[6] ,n3[6]);
    nand g712(n511 ,n10[8] ,n487);
    not g713(n247 ,n648);
    not g714(n260 ,n11[5]);
    nand g715(n307 ,n10[11] ,n285);
    not g716(n249 ,n622);
    nand g717(n203 ,n187 ,n202);
    nand g718(n436 ,n359 ,n360);
    nand g719(n158 ,n140 ,n157);
    nand g720(n349 ,n284 ,n308);
    xnor g721(n598 ,n131 ,n151);
    nand g722(n378 ,n580 ,n296);
    dff g723(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n549), .Q(n11[1]));
    not g724(n223 ,n642);
    not g725(n93 ,n92);
    nand g726(n103 ,n83 ,n102);
    nand g727(n280 ,n14[0] ,n264);
    xnor g728(n665 ,n13[2] ,n219);
    nand g729(n454 ,n9[4] ,n331);
    xnor g730(n622 ,n79 ,n108);
    xnor g731(n184 ,n599 ,n12[4]);
    nand g732(n483 ,n449 ,n414);
    xor g733(n628 ,n3[2] ,n10[2]);
    nand g734(n445 ,n9[11] ,n347);
    nand g735(n525 ,n11[10] ,n520);
    dff g736(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n550), .Q(n11[0]));
    nor g737(n411 ,n366 ,n337);
    xnor g738(n6[6] ,n575 ,n9[6]);
    xnor g739(n620 ,n104 ,n84);
    nand g740(n677 ,n3[5] ,n675);
    nand g741(n365 ,n13[0] ,n299);
    nor g742(n682 ,n668 ,n681);
    nand g743(n679 ,n3[6] ,n678);
    xnor g744(n10[4] ,n3[4] ,n674);
    nand g745(n176 ,n609 ,n12[9]);
    nor g746(n385 ,n249 ,n295);
    xnor g747(n648 ,n35 ,n61);
    nand g748(n465 ,n7[6] ,n342);
    dff g749(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n542), .Q(n11[9]));
    nand g750(n508 ,n10[11] ,n487);
    nor g751(n330 ,n254 ,n312);
    nand g752(n555 ,n11[11] ,n12[11]);
    nand g753(n501 ,n377 ,n395);
    not g754(n269 ,n7[2]);
    xnor g755(n132 ,n2[9] ,n3[9]);
    dff g756(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n544), .Q(n11[11]));
    nand g757(n359 ,n13[2] ,n299);
    xnor g758(n31 ,n658 ,n12[6]);
    nand g759(n449 ,n9[8] ,n349);
    nand g760(n178 ,n591 ,n10[1]);
    nand g761(n519 ,n3[0] ,n487);
    not g762(n293 ,n292);
    nand g763(n479 ,n446 ,n412);
    not g764(n42 ,n41);
    xnor g765(n649 ,n44 ,n63);
    nor g766(n422 ,n379 ,n330);
    nand g767(n397 ,n302 ,n321);
    nand g768(n21 ,n661 ,n12[9]);
    nand g769(n532 ,n11[4] ,n520);
    nor g770(n389 ,n333 ,n328);
    xor g771(n641 ,n39 ,n47);
    nor g772(n54 ,n30 ,n53);
    nand g773(n352 ,n640 ,n296);
    or g774(n271 ,n11[0] ,n11[1]);
    dff g775(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n484), .Q(n9[7]));
    xnor g776(n646 ,n37 ,n57);
    nand g777(n672 ,n3[2] ,n671);
    dff g778(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n480), .Q(n8[5]));
    xor g779(n565 ,n3[0] ,n553);
    xnor g780(n610 ,n134 ,n163);
    xnor g781(n645 ,n55 ,n31);
    nor g782(n10[9] ,n683 ,n685);
    nand g783(n543 ,n511 ,n527);
    dff g784(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n539), .Q(n11[12]));
    nand g785(n289 ,n10[2] ,n279);
    nand g786(n73 ,n637 ,n10[11]);
    not g787(n687 ,n686);
    dff g788(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n437), .Q(n13[1]));
    nand g789(n536 ,n11[6] ,n520);
    nor g790(n286 ,n14[2] ,n278);
    nand g791(n78 ,n627 ,n12[2]);
    nand g792(n329 ,n284 ,n309);
    dff g793(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n502), .Q(n9[0]));
    dff g794(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n493), .Q(n7[9]));
    xnor g795(n602 ,n137 ,n155);
    nand g796(n46 ,n26 ,n34);
    nand g797(n451 ,n9[6] ,n342);
    nor g798(n52 ,n29 ,n51);
    xnor g799(n584 ,n190 ,n206);
    nand g800(n563 ,n11[5] ,n12[5]);
endmodule
