module top (n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [3:0] n6;
    wire [2:0] n7;
    wire [3:0] n8;
    wire [31:0] n9;
    wire [31:0] n10;
    wire [31:0] n11;
    wire n12, n13, n14, n15, n16, n17, n18, n19;
    wire n20, n21, n22, n23, n24, n25, n26, n27;
    wire n28, n29, n30, n31, n32, n33, n34, n35;
    wire n36, n37, n38, n39, n40, n41, n42, n43;
    wire n44, n45, n46, n47, n48, n49, n50, n51;
    wire n52, n53, n54, n55, n56, n57, n58, n59;
    wire n60, n61, n62, n63, n64, n65, n66, n67;
    wire n68, n69, n70, n71, n72, n73, n74, n75;
    wire n76, n77, n78, n79, n80, n81, n82, n83;
    wire n84, n85, n86, n87, n88, n89, n90, n91;
    wire n92, n93, n94, n95, n96, n97, n98, n99;
    wire n100, n101, n102, n103, n104, n105, n106, n107;
    wire n108, n109, n110, n111, n112, n113, n114, n115;
    wire n116, n117, n118, n119, n120, n121, n122, n123;
    wire n124, n125, n126, n127, n128, n129, n130, n131;
    wire n132, n133, n134, n135, n136, n137, n138, n139;
    wire n140, n141, n142, n143, n144, n145, n146, n147;
    wire n148, n149, n150, n151, n152, n153, n154, n155;
    wire n156, n157, n158, n159, n160, n161, n162, n163;
    wire n164, n165, n166, n167, n168, n169, n170, n171;
    wire n172, n173, n174, n175, n176, n177, n178, n179;
    wire n180, n181, n182, n183, n184, n185, n186, n187;
    wire n188, n189, n190, n191, n192, n193, n194, n195;
    wire n196, n197, n198, n199, n200, n201, n202, n203;
    wire n204, n205, n206, n207, n208, n209, n210, n211;
    wire n212, n213, n214, n215, n216, n217, n218, n219;
    wire n220, n221, n222, n223, n224, n225, n226, n227;
    wire n228, n229, n230, n231, n232, n233, n234, n235;
    wire n236, n237, n238, n239, n240, n241, n242, n243;
    wire n244, n245, n246, n247, n248, n249, n250, n251;
    wire n252, n253, n254, n255, n256, n257, n258, n259;
    wire n260, n261, n262, n263, n264, n265, n266, n267;
    wire n268, n269, n270, n271, n272, n273, n274, n275;
    wire n276, n277, n278, n279, n280, n281, n282, n283;
    wire n284, n285, n286, n287, n288, n289, n290, n291;
    wire n292, n293, n294, n295, n296, n297, n298, n299;
    wire n300, n301, n302, n303, n304, n305, n306, n307;
    wire n308, n309, n310, n311, n312, n313, n314, n315;
    wire n316, n317, n318, n319, n320, n321, n322, n323;
    wire n324, n325, n326, n327, n328, n329, n330, n331;
    wire n332, n333, n334, n335, n336, n337, n338, n339;
    wire n340, n341, n342, n343, n344, n345, n346, n347;
    wire n348, n349, n350, n351, n352, n353, n354, n355;
    wire n356, n357, n358, n359, n360, n361, n362, n363;
    wire n364, n365, n366, n367, n368, n369, n370, n371;
    wire n372, n373, n374, n375, n376, n377, n378, n379;
    wire n380, n381, n382, n383, n384, n385, n386, n387;
    wire n388, n389, n390, n391, n392, n393, n394, n395;
    wire n396, n397, n398, n399, n400, n401, n402, n403;
    wire n404, n405, n406, n407, n408, n409, n410, n411;
    wire n412, n413, n414, n415, n416, n417, n418, n419;
    wire n420, n421, n422, n423, n424, n425, n426, n427;
    wire n428, n429, n430, n431, n432, n433, n434, n435;
    wire n436, n437, n438, n439, n440, n441, n442, n443;
    wire n444, n445, n446, n447, n448, n449, n450, n451;
    wire n452, n453, n454, n455, n456, n457, n458, n459;
    wire n460, n461, n462, n463, n464, n465, n466, n467;
    wire n468, n469, n470, n471, n472, n473, n474, n475;
    wire n476, n477, n478, n479, n480, n481, n482, n483;
    wire n484, n485, n486, n487, n488, n489, n490, n491;
    wire n492, n493, n494, n495, n496, n497, n498, n499;
    wire n500, n501, n502, n503, n504, n505, n506, n507;
    wire n508, n509, n510, n511, n512, n513, n514, n515;
    wire n516, n517, n518, n519, n520, n521, n522, n523;
    wire n524, n525, n526, n527, n528, n529, n530, n531;
    wire n532, n533, n534, n535, n536, n537, n538, n539;
    wire n540, n541, n542, n543, n544, n545, n546, n547;
    wire n548, n549, n550, n551, n552, n553, n554, n555;
    wire n556, n557, n558, n559, n560, n561, n562, n563;
    wire n564, n565, n566, n567, n568, n569, n570, n571;
    wire n572, n573, n574, n575, n576, n577, n578, n579;
    wire n580, n581, n582, n583, n584, n585, n586, n587;
    wire n588, n589, n590, n591, n592, n593, n594, n595;
    wire n596, n597, n598, n599, n600, n601, n602, n603;
    wire n604, n605, n606, n607, n608, n609, n610, n611;
    wire n612, n613, n614, n615, n616, n617, n618, n619;
    wire n620, n621, n622, n623, n624, n625, n626, n627;
    wire n628, n629, n630, n631, n632, n633, n634, n635;
    wire n636, n637, n638, n639, n640, n641, n642, n643;
    wire n644, n645, n646, n647, n648, n649, n650, n651;
    wire n652, n653, n654, n655, n656, n657, n658, n659;
    wire n660, n661, n662, n663, n664, n665, n666, n667;
    wire n668, n669, n670, n671, n672, n673, n674, n675;
    wire n676, n677, n678, n679, n680, n681, n682, n683;
    wire n684, n685, n686, n687, n688, n689, n690, n691;
    wire n692, n693, n694, n695, n696, n697, n698, n699;
    wire n700, n701, n702, n703, n704, n705, n706, n707;
    wire n708, n709, n710, n711, n712, n713, n714, n715;
    wire n716, n717, n718, n719, n720, n721, n722, n723;
    wire n724, n725, n726, n727, n728, n729, n730, n731;
    wire n732, n733, n734, n735, n736, n737, n738, n739;
    wire n740, n741, n742, n743, n744, n745, n746, n747;
    wire n748, n749, n750, n751, n752, n753, n754, n755;
    wire n756, n757, n758, n759, n760, n761, n762, n763;
    wire n764, n765, n766, n767, n768, n769, n770, n771;
    wire n772, n773, n774, n775, n776, n777, n778, n779;
    wire n780, n781, n782, n783, n784, n785, n786, n787;
    wire n788, n789, n790, n791, n792, n793, n794, n795;
    wire n796, n797, n798, n799, n800, n801, n802, n803;
    wire n804, n805, n806, n807, n808, n809, n810, n811;
    wire n812, n813, n814, n815, n816, n817, n818, n819;
    wire n820, n821, n822, n823, n824, n825, n826, n827;
    wire n828, n829, n830, n831, n832, n833, n834, n835;
    wire n836, n837, n838, n839, n840, n841, n842, n843;
    wire n844, n845, n846, n847, n848, n849, n850, n851;
    wire n852, n853, n854, n855, n856, n857, n858, n859;
    wire n860, n861, n862, n863, n864, n865, n866, n867;
    wire n868, n869, n870, n871, n872, n873, n874, n875;
    wire n876, n877, n878, n879, n880, n881, n882, n883;
    wire n884, n885, n886, n887, n888, n889, n890, n891;
    wire n892, n893, n894, n895, n896, n897, n898, n899;
    wire n900, n901, n902, n903, n904, n905, n906, n907;
    wire n908, n909, n910, n911, n912, n913, n914, n915;
    wire n916, n917, n918, n919, n920, n921, n922, n923;
    wire n924, n925, n926, n927, n928, n929, n930, n931;
    wire n932, n933, n934, n935, n936, n937, n938, n939;
    wire n940, n941, n942, n943, n944, n945, n946, n947;
    wire n948, n949, n950, n951, n952, n953, n954, n955;
    wire n956, n957, n958, n959, n960, n961, n962, n963;
    wire n964, n965, n966, n967, n968, n969, n970, n971;
    wire n972, n973, n974, n975, n976, n977, n978, n979;
    wire n980, n981, n982, n983, n984, n985, n986, n987;
    wire n988, n989, n990, n991, n992, n993, n994, n995;
    wire n996, n997, n998, n999, n1000, n1001, n1002, n1003;
    wire n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011;
    wire n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
    wire n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
    wire n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
    wire n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
    wire n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051;
    wire n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059;
    wire n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067;
    wire n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075;
    wire n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083;
    wire n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091;
    wire n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099;
    wire n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107;
    wire n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115;
    wire n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123;
    wire n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131;
    wire n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139;
    wire n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147;
    wire n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155;
    wire n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163;
    wire n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171;
    wire n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179;
    wire n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187;
    wire n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195;
    wire n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203;
    wire n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
    wire n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219;
    wire n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227;
    wire n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235;
    wire n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243;
    wire n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251;
    wire n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259;
    wire n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267;
    wire n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275;
    wire n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;
    wire n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291;
    wire n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;
    wire n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307;
    wire n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315;
    wire n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323;
    wire n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331;
    wire n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;
    wire n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;
    wire n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;
    wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
    wire n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;
    wire n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;
    wire n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387;
    wire n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395;
    wire n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403;
    wire n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411;
    wire n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419;
    wire n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427;
    wire n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435;
    wire n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443;
    wire n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451;
    wire n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459;
    wire n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467;
    wire n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475;
    wire n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483;
    wire n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491;
    wire n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499;
    wire n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507;
    wire n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515;
    wire n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523;
    wire n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531;
    wire n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539;
    wire n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547;
    wire n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555;
    wire n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563;
    wire n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571;
    wire n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579;
    wire n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587;
    wire n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595;
    wire n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603;
    wire n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611;
    wire n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619;
    wire n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627;
    wire n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635;
    wire n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643;
    wire n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651;
    wire n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659;
    wire n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667;
    wire n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675;
    wire n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683;
    wire n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691;
    wire n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699;
    wire n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707;
    wire n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715;
    wire n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723;
    wire n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731;
    wire n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739;
    wire n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747;
    wire n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755;
    wire n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763;
    wire n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771;
    wire n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779;
    wire n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787;
    wire n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795;
    wire n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803;
    wire n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811;
    wire n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819;
    wire n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827;
    wire n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835;
    wire n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843;
    wire n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851;
    wire n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859;
    wire n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867;
    wire n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875;
    wire n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883;
    wire n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891;
    wire n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899;
    wire n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907;
    wire n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915;
    wire n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923;
    wire n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931;
    wire n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939;
    wire n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947;
    wire n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955;
    wire n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963;
    wire n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971;
    wire n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979;
    wire n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987;
    wire n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995;
    wire n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003;
    wire n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011;
    wire n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019;
    wire n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027;
    wire n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035;
    wire n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043;
    wire n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051;
    wire n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059;
    wire n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067;
    wire n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075;
    wire n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083;
    wire n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091;
    wire n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099;
    wire n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107;
    wire n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115;
    wire n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123;
    wire n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131;
    wire n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139;
    wire n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147;
    wire n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155;
    wire n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163;
    wire n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171;
    wire n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179;
    wire n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187;
    wire n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195;
    wire n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203;
    wire n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211;
    wire n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219;
    wire n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227;
    wire n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235;
    wire n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243;
    wire n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251;
    wire n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259;
    wire n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267;
    wire n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275;
    wire n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283;
    wire n2284;
    not g0(n1244 ,n1115);
    nand g1(n1774 ,n2005 ,n1666);
    nand g2(n396 ,n8[2] ,n395);
    nor g3(n572 ,n460 ,n1);
    nand g4(n721 ,n2[96] ,n629);
    not g5(n369 ,n368);
    nand g6(n2171 ,n4[46] ,n2168);
    dff g7(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n522), .Q(n9[3]));
    nand g8(n1166 ,n752 ,n775);
    xor g9(n2065 ,n2[0] ,n2[64]);
    nand g10(n1071 ,n1904 ,n729);
    nand g11(n1142 ,n722 ,n788);
    nor g12(n490 ,n3[1] ,n6[1]);
    not g13(n1656 ,n1651);
    or g14(n1646 ,n1616 ,n1451);
    nand g15(n895 ,n1858 ,n409);
    nand g16(n610 ,n411 ,n607);
    dff g17(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1342), .Q(n4[24]));
    nand g18(n891 ,n1845 ,n408);
    nand g19(n1838 ,n2143 ,n2142);
    dff g20(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1577), .Q(n3[48]));
    xnor g21(n103 ,n2[34] ,n2[98]);
    nor g22(n158 ,n30 ,n157);
    nand g23(n662 ,n3[13] ,n621);
    not g24(n413 ,n730);
    nand g25(n1782 ,n1669 ,n3[9]);
    nand g26(n1149 ,n834 ,n820);
    nand g27(n789 ,n3[53] ,n621);
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1632), .Q(n3[22]));
    not g29(n2216 ,n11[4]);
    not g30(n1027 ,n1028);
    nand g31(n1976 ,n1794 ,n1791);
    nor g32(n558 ,n419 ,n1);
    not g33(n1256 ,n1133);
    nand g34(n799 ,n2[86] ,n629);
    nand g35(n1716 ,n1669 ,n3[25]);
    xnor g36(n2042 ,n85 ,n224);
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1586), .Q(n3[42]));
    nand g38(n766 ,n2[71] ,n406);
    nand g39(n713 ,n2[74] ,n406);
    nand g40(n705 ,n2[109] ,n406);
    nand g41(n1860 ,n2187 ,n2186);
    nand g42(n2147 ,n4[34] ,n2144);
    nand g43(n392 ,n2000 ,n391);
    nand g44(n800 ,n3[45] ,n621);
    not g45(n1655 ,n1650);
    nand g46(n1187 ,n5[35] ,n400);
    not g47(n1553 ,n1512);
    xnor g48(n2026 ,n78 ,n192);
    nand g49(n384 ,n1996 ,n383);
    xnor g50(n75 ,n2[63] ,n2[127]);
    nand g51(n1429 ,n1160 ,n1007);
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n556), .Q(n9[9]));
    nand g53(n2091 ,n4[6] ,n2088);
    nand g54(n313 ,n1956 ,n311);
    not g55(n1410 ,n1383);
    nand g56(n587 ,n2[1] ,n6[1]);
    nand g57(n1177 ,n596 ,n647);
    nand g58(n1109 ,n803 ,n691);
    not g59(n1235 ,n1104);
    not g60(n626 ,n625);
    nor g61(n41 ,n2[25] ,n2[89]);
    nor g62(n224 ,n60 ,n223);
    nand g63(n1765 ,n2059 ,n1666);
    nand g64(n1096 ,n1894 ,n410);
    nor g65(n637 ,n497 ,n412);
    nor g66(n538 ,n483 ,n1);
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1423), .Q(n5[52]));
    nor g68(n188 ,n41 ,n187);
    nand g69(n2075 ,n6[2] ,n2070);
    nand g70(n627 ,n619 ,n618);
    nand g71(n1025 ,n1840 ,n408);
    nand g72(n1436 ,n1180 ,n937);
    xor g73(n1906 ,n1974 ,n341);
    nand g74(n1308 ,n890 ,n1237);
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1560), .Q(n3[6]));
    nor g76(n207 ,n90 ,n206);
    nand g77(n978 ,n1886 ,n405);
    not g78(n377 ,n376);
    not g79(n470 ,n2[70]);
    xnor g80(n1807 ,n2080 ,n2076);
    nand g81(n370 ,n1989 ,n369);
    nor g82(n537 ,n448 ,n1);
    not g83(n440 ,n2[35]);
    nor g84(n257 ,n95 ,n256);
    nand g85(n2161 ,n4[41] ,n2158);
    nand g86(n591 ,n8[2] ,n8[3]);
    nand g87(n786 ,n3[57] ,n398);
    nand g88(n1608 ,n934 ,n1303);
    nand g89(n1045 ,n1872 ,n405);
    nand g90(n989 ,n2[61] ,n403);
    or g91(n266 ,n1941 ,n1937);
    not g92(n1281 ,n1178);
    nand g93(n1708 ,n1668 ,n3[23]);
    nand g94(n839 ,n2[23] ,n403);
    not g95(n477 ,n2[68]);
    nor g96(n615 ,n604 ,n608);
    nand g97(n1082 ,n1899 ,n729);
    nand g98(n1743 ,n1668 ,n3[31]);
    nand g99(n1973 ,n1772 ,n1697);
    nand g100(n760 ,n2[75] ,n406);
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1479), .Q(n5[8]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1466), .Q(n5[13]));
    xnor g103(n1916 ,n1984 ,n360);
    nand g104(n1769 ,n6[1] ,n1668);
    nand g105(n1603 ,n1090 ,n1557);
    nand g106(n1170 ,n754 ,n771);
    nand g107(n1189 ,n5[34] ,n400);
    nand g108(n1423 ,n1146 ,n855);
    xor g109(n1920 ,n1988 ,n366);
    nand g110(n285 ,n267 ,n284);
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n563), .Q(n11[4]));
    nand g112(n1348 ,n985 ,n1274);
    nand g113(n1303 ,n3[2] ,n1030);
    nor g114(n220 ,n47 ,n219);
    nand g115(n1064 ,n1842 ,n729);
    nand g116(n1740 ,n1668 ,n3[47]);
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1581), .Q(n3[45]));
    nand g118(n309 ,n1953 ,n308);
    nor g119(n53 ,n2[58] ,n2[122]);
    nand g120(n1818 ,n2103 ,n2102);
    nand g121(n1633 ,n840 ,n1394);
    xnor g122(n77 ,n2[46] ,n2[110]);
    nor g123(n193 ,n78 ,n192);
    nand g124(n1839 ,n2145 ,n2144);
    nor g125(n147 ,n105 ,n146);
    nand g126(n2123 ,n4[22] ,n2120);
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1319), .Q(n4[45]));
    nand g128(n1682 ,n1669 ,n3[61]);
    nand g129(n1720 ,n1669 ,n3[26]);
    not g130(n1402 ,n1375);
    nor g131(n72 ,n2[59] ,n2[123]);
    nor g132(n203 ,n98 ,n202);
    nand g133(n2191 ,n4[56] ,n2188);
    nor g134(n561 ,n469 ,n1);
    nand g135(n1438 ,n1184 ,n941);
    not g136(n482 ,n2068);
    xnor g137(n2054 ,n94 ,n248);
    nor g138(n2230 ,n2218 ,n9[15]);
    nand g139(n814 ,n3[37] ,n398);
    nand g140(n857 ,n2[15] ,n403);
    nand g141(n678 ,n2[126] ,n406);
    nor g142(n501 ,n5[0] ,n6[0]);
    nand g143(n1457 ,n1210 ,n970);
    nand g144(n1174 ,n5[40] ,n732);
    xnor g145(n102 ,n2[4] ,n2[68]);
    nand g146(n1771 ,n1669 ,n3[6]);
    nor g147(n1295 ,n486 ,n1028);
    nand g148(n979 ,n1855 ,n410);
    nand g149(n663 ,n2[70] ,n406);
    nand g150(n1792 ,n2010 ,n1666);
    nor g151(n492 ,n8[0] ,n1);
    nand g152(n2247 ,n11[11] ,n11[10]);
    nand g153(n897 ,n1870 ,n409);
    nand g154(n690 ,n2[118] ,n406);
    nand g155(n685 ,n2[121] ,n406);
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n567), .Q(n11[8]));
    nand g157(n844 ,n1891 ,n410);
    nor g158(n2203 ,n4[62] ,n2201);
    nand g159(n757 ,n2[77] ,n629);
    nand g160(n1054 ,n2[40] ,n730);
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1346), .Q(n4[20]));
    nand g162(n1317 ,n960 ,n1245);
    not g163(n1411 ,n1384);
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n4[21]));
    xnor g165(n2080 ,n6[1] ,n4[1]);
    nand g166(n1324 ,n906 ,n1252);
    nand g167(n749 ,n2[84] ,n629);
    nand g168(n805 ,n3[42] ,n398);
    nand g169(n1980 ,n1698 ,n1695);
    or g170(n2192 ,n4[57] ,n2190);
    xnor g171(n135 ,n2[22] ,n2[86]);
    nand g172(n924 ,n1826 ,n729);
    nor g173(n352 ,n273 ,n350);
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1576), .Q(n3[49]));
    nand g175(n675 ,n3[5] ,n621);
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1311), .Q(n4[52]));
    nand g177(n929 ,n1910 ,n405);
    nor g178(n507 ,n3[3] ,n6[3]);
    nand g179(n2277 ,n2264 ,n2261);
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n4[17]));
    nand g181(n1344 ,n1016 ,n1270);
    nand g182(n305 ,n1951 ,n304);
    nand g183(n1224 ,n5[8] ,n732);
    not g184(n450 ,n2[76]);
    nand g185(n2193 ,n4[57] ,n2190);
    nand g186(n1196 ,n590 ,n637);
    nand g187(n1974 ,n1694 ,n1777);
    or g188(n2090 ,n4[6] ,n2088);
    nand g189(n74 ,n2[0] ,n2[64]);
    nor g190(n2200 ,n4[61] ,n2198);
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1485), .Q(n5[6]));
    nand g192(n1568 ,n1001 ,n1526);
    nand g193(n944 ,n1905 ,n731);
    not g194(n1266 ,n1151);
    xnor g195(n1932 ,n2000 ,n390);
    nand g196(n274 ,n1955 ,n1954);
    xnor g197(n1914 ,n1982 ,n356);
    nand g198(n1735 ,n2045 ,n1665);
    nand g199(n1059 ,n2[38] ,n403);
    nand g200(n312 ,n1954 ,n310);
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1629), .Q(n3[19]));
    nand g202(n1049 ,n2[42] ,n730);
    nand g203(n1997 ,n1718 ,n1706);
    or g204(n2092 ,n4[7] ,n2090);
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n562), .Q(n11[13]));
    nor g206(n574 ,n440 ,n1);
    nand g207(n651 ,n4[63] ,n402);
    nand g208(n1210 ,n5[22] ,n732);
    nand g209(n367 ,n1986 ,n365);
    nand g210(n976 ,n1888 ,n405);
    nand g211(n1788 ,n2009 ,n1666);
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1360), .Q(n4[6]));
    nand g213(n1309 ,n894 ,n1238);
    nor g214(n259 ,n114 ,n258);
    xnor g215(n1898 ,n1966 ,n331);
    xnor g216(n86 ,n2[54] ,n2[118]);
    nand g217(n756 ,n2[78] ,n406);
    nand g218(n761 ,n4[4] ,n620);
    nand g219(n585 ,n4[1] ,n6[1]);
    nand g220(n599 ,n3[0] ,n6[0]);
    nand g221(n671 ,n3[8] ,n621);
    xnor g222(n1928 ,n1996 ,n382);
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1438), .Q(n5[36]));
    xnor g224(n1901 ,n1969 ,n337);
    nand g225(n329 ,n1964 ,n328);
    nand g226(n1601 ,n1086 ,n1555);
    nor g227(n2237 ,n11[31] ,n11[30]);
    or g228(n2190 ,n4[56] ,n2188);
    nand g229(n1178 ,n760 ,n772);
    nand g230(n140 ,n16 ,n139);
    nand g231(n2097 ,n4[9] ,n2094);
    nor g232(n488 ,n3[0] ,n6[0]);
    not g233(n1276 ,n1168);
    nand g234(n388 ,n1998 ,n387);
    nand g235(n378 ,n1993 ,n377);
    nor g236(n508 ,n456 ,n1);
    xnor g237(n2035 ,n112 ,n210);
    nand g238(n1150 ,n5[49] ,n400);
    nand g239(n1421 ,n1144 ,n915);
    nand g240(n1190 ,n5[33] ,n400);
    xnor g241(n84 ,n2[31] ,n2[95]);
    not g242(n1405 ,n1378);
    nand g243(n1047 ,n1913 ,n408);
    nor g244(n240 ,n37 ,n239);
    nor g245(n13 ,n2[29] ,n2[93]);
    nor g246(n625 ,n7[0] ,n619);
    not g247(n363 ,n362);
    nand g248(n706 ,n4[41] ,n402);
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1587), .Q(n3[41]));
    not g250(n445 ,n2[54]);
    not g251(n451 ,n2[61]);
    nand g252(n1489 ,n793 ,n928);
    nor g253(n1029 ,n1 ,n734);
    nand g254(n1418 ,n1137 ,n912);
    nand g255(n1363 ,n4[3] ,n1029);
    nand g256(n2121 ,n4[21] ,n2118);
    nor g257(n577 ,n420 ,n1);
    nand g258(n1365 ,n4[1] ,n1029);
    nor g259(n17 ,n2[16] ,n2[80]);
    nand g260(n823 ,n3[30] ,n398);
    nand g261(n1702 ,n2041 ,n1665);
    not g262(n2204 ,n9[23]);
    dff g263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n576), .Q(n11[27]));
    xnor g264(n2059 ,n114 ,n258);
    nand g265(n142 ,n73 ,n141);
    nor g266(n243 ,n129 ,n242);
    nor g267(n159 ,n115 ,n158);
    nand g268(n289 ,n1942 ,n288);
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1453), .Q(n5[25]));
    nor g270(n496 ,n2[67] ,n6[3]);
    xnor g271(n1919 ,n367 ,n1987);
    nand g272(n1390 ,n584 ,n836);
    nor g273(n578 ,n451 ,n1);
    nor g274(n144 ,n68 ,n143);
    nor g275(n836 ,n500 ,n413);
    nor g276(n489 ,n2[64] ,n6[0]);
    nand g277(n380 ,n1994 ,n379);
    nand g278(n2181 ,n4[51] ,n2178);
    dff g279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1356), .Q(n4[10]));
    nand g280(n1466 ,n1219 ,n988);
    nand g281(n1226 ,n5[6] ,n732);
    xnor g282(n2024 ,n83 ,n188);
    nand g283(n832 ,n3[25] ,n398);
    or g284(n2274 ,n2258 ,n2265);
    nand g285(n1975 ,n1787 ,n1783);
    not g286(n340 ,n339);
    nand g287(n854 ,n1886 ,n410);
    or g288(n278 ,n275 ,n268);
    xnor g289(n1929 ,n1997 ,n384);
    or g290(n2168 ,n4[45] ,n2166);
    nand g291(n1948 ,n1786 ,n1785);
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1660), .Q(n1663));
    not g293(n455 ,n2[94]);
    nand g294(n903 ,n1932 ,n731);
    nand g295(n1736 ,n6[0] ,n1669);
    not g296(n1934 ,n1736);
    nand g297(n2105 ,n4[13] ,n2102);
    not g298(n385 ,n384);
    nand g299(n1117 ,n703 ,n770);
    nor g300(n232 ,n12 ,n231);
    nand g301(n1670 ,n1669 ,n3[13]);
    nand g302(n1191 ,n769 ,n761);
    nor g303(n513 ,n442 ,n1);
    nand g304(n2232 ,n9[5] ,n2209);
    nand g305(n1389 ,n587 ,n835);
    dff g306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n557), .Q(n11[7]));
    nand g307(n1729 ,n1668 ,n3[28]);
    nand g308(n1094 ,n1895 ,n729);
    not g309(n1413 ,n1386);
    xnor g310(n1890 ,n1958 ,n315);
    nand g311(n1479 ,n1224 ,n1005);
    nor g312(n251 ,n106 ,n250);
    nand g313(n699 ,n2[112] ,n406);
    dff g314(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1596), .Q(n3[33]));
    xnor g315(n6[1] ,n10[29] ,n2284);
    dff g316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1335), .Q(n4[30]));
    nand g317(n1325 ,n891 ,n1253);
    nand g318(n1506 ,n815 ,n1065);
    nand g319(n319 ,n1959 ,n318);
    nand g320(n1578 ,n1038 ,n1536);
    nor g321(n524 ,n470 ,n1);
    nand g322(n899 ,n1859 ,n410);
    nand g323(n1194 ,n589 ,n636);
    nand g324(n1967 ,n1734 ,n1732);
    nand g325(n1686 ,n2039 ,n1665);
    nand g326(n650 ,n3[23] ,n621);
    dff g327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1630), .Q(n3[20]));
    dff g328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1322), .Q(n4[42]));
    nand g329(n668 ,n3[10] ,n621);
    dff g330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1573), .Q(n3[52]));
    dff g331(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1358), .Q(n4[8]));
    xor g332(n1888 ,n1956 ,n311);
    nand g333(n1378 ,n665 ,n865);
    nand g334(n1192 ,n588 ,n635);
    not g335(n399 ,n732);
    nand g336(n1060 ,n1908 ,n408);
    nand g337(n1376 ,n661 ,n860);
    nor g338(n642 ,n623 ,n631);
    dff g339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1600), .Q(n3[29]));
    nand g340(n315 ,n1957 ,n314);
    not g341(n330 ,n329);
    dff g342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n555), .Q(n9[11]));
    xnor g343(n2043 ,n79 ,n226);
    nand g344(n1020 ,n2[51] ,n403);
    nand g345(n1977 ,n1674 ,n1671);
    not g346(n304 ,n303);
    xnor g347(n107 ,n2[48] ,n2[112]);
    nand g348(n1705 ,n1668 ,n3[43]);
    nand g349(n1715 ,n2023 ,n1665);
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1658), .Q(n5[1]));
    nand g351(n1133 ,n717 ,n812);
    not g352(n1251 ,n1124);
    nand g353(n1430 ,n1165 ,n1026);
    nand g354(n1299 ,n3[3] ,n1030);
    nor g355(n217 ,n96 ,n216);
    nand g356(n1590 ,n1058 ,n1544);
    nand g357(n937 ,n1908 ,n405);
    nand g358(n1026 ,n1914 ,n405);
    nor g359(n525 ,n435 ,n1);
    xnor g360(n129 ,n2[53] ,n2[117]);
    not g361(n322 ,n321);
    dff g362(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1604), .Q(n3[25]));
    nand g363(n1075 ,n2[32] ,n403);
    xnor g364(n2018 ,n131 ,n176);
    nor g365(n250 ,n67 ,n249);
    nand g366(n1813 ,n2093 ,n2092);
    xnor g367(n2060 ,n91 ,n260);
    nand g368(n683 ,n2[122] ,n629);
    nand g369(n945 ,n1812 ,n410);
    nand g370(n1381 ,n669 ,n871);
    or g371(n2106 ,n4[14] ,n2104);
    xnor g372(n1895 ,n1963 ,n325);
    nand g373(n694 ,n2[115] ,n406);
    nor g374(n205 ,n103 ,n204);
    nand g375(n1820 ,n2107 ,n2106);
    nor g376(n201 ,n89 ,n200);
    nand g377(n2149 ,n4[35] ,n2146);
    dff g378(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n525), .Q(n9[8]));
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n578), .Q(n11[29]));
    dff g380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n508), .Q(n9[25]));
    nand g381(n1599 ,n1077 ,n1552);
    nand g382(n1991 ,n1699 ,n1693);
    xnor g383(n2006 ,n126 ,n152);
    nor g384(n623 ,n7[0] ,n618);
    nand g385(n1783 ,n2035 ,n1666);
    not g386(n1664 ,n7[1]);
    xnor g387(n1877 ,n1945 ,n293);
    nand g388(n1155 ,n5[48] ,n732);
    dff g389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1567), .Q(n3[58]));
    xnor g390(n2029 ,n84 ,n198);
    nand g391(n2185 ,n4[53] ,n2182);
    nand g392(n1949 ,n1789 ,n1788);
    nand g393(n1834 ,n2135 ,n2134);
    dff g394(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1447), .Q(n5[29]));
    nand g395(n1010 ,n1877 ,n405);
    nand g396(n1211 ,n5[21] ,n732);
    nand g397(n2243 ,n11[27] ,n2207);
    not g398(n1541 ,n1498);
    not g399(n1252 ,n1126);
    dff g400(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1302), .Q(n4[61]));
    not g401(n1238 ,n1108);
    dff g402(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1583), .Q(n3[44]));
    xnor g403(n2044 ,n77 ,n228);
    dff g404(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1595), .Q(n3[34]));
    nor g405(n227 ,n79 ,n226);
    nand g406(n1492 ,n5[3] ,n1032);
    nand g407(n1213 ,n5[19] ,n400);
    not g408(n1243 ,n1114);
    dff g409(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1434), .Q(n5[40]));
    xnor g410(n2036 ,n117 ,n212);
    nor g411(n495 ,n4[3] ,n6[3]);
    nand g412(n1340 ,n918 ,n1266);
    nand g413(n1943 ,n1767 ,n1766);
    nand g414(n893 ,n1862 ,n410);
    nor g415(n635 ,n496 ,n412);
    nand g416(n1305 ,n950 ,n1233);
    not g417(n2069 ,n4[1]);
    dff g418(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n536), .Q(n8[3]));
    not g419(n1524 ,n1471);
    nand g420(n1040 ,n1916 ,n729);
    not g421(n1278 ,n1172);
    nand g422(n772 ,n4[11] ,n402);
    nor g423(n59 ,n2[53] ,n2[117]);
    nand g424(n796 ,n3[47] ,n621);
    xnor g425(n1872 ,n279 ,n284);
    nand g426(n804 ,n3[43] ,n621);
    nand g427(n2081 ,n2076 ,n2080);
    dff g428(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1328), .Q(n4[36]));
    xnor g429(n111 ,n2[9] ,n2[73]);
    nand g430(n619 ,n1663 ,n609);
    dff g431(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1351), .Q(n4[15]));
    not g432(n1551 ,n1510);
    dff g433(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1348), .Q(n4[18]));
    nand g434(n658 ,n4[6] ,n402);
    nand g435(n386 ,n1997 ,n385);
    nor g436(n2279 ,n2273 ,n2275);
    nand g437(n1361 ,n917 ,n1287);
    not g438(n1556 ,n1515);
    xnor g439(n1887 ,n312 ,n1955);
    nand g440(n711 ,n2[103] ,n406);
    xnor g441(n1927 ,n1995 ,n380);
    not g442(n416 ,n2[64]);
    nor g443(n1292 ,n501 ,n1031);
    nand g444(n2197 ,n4[59] ,n2194);
    not g445(n1262 ,n1143);
    nand g446(n1745 ,n2054 ,n1665);
    nand g447(n688 ,n4[40] ,n402);
    nand g448(n2125 ,n4[23] ,n2122);
    nand g449(n702 ,n4[38] ,n620);
    nand g450(n1372 ,n664 ,n850);
    nand g451(n1465 ,n1218 ,n981);
    nand g452(n774 ,n4[14] ,n620);
    nand g453(n364 ,n1985 ,n363);
    nand g454(n1942 ,n1712 ,n1761);
    nand g455(n2074 ,n6[3] ,n2072);
    nor g456(n22 ,n2[34] ,n2[98]);
    not g457(n296 ,n295);
    nor g458(n2280 ,n2277 ,n2271);
    nor g459(n161 ,n116 ,n160);
    xnor g460(n2005 ,n108 ,n150);
    not g461(n433 ,n2[91]);
    nand g462(n1704 ,n1668 ,n3[22]);
    nand g463(n1145 ,n725 ,n726);
    not g464(n389 ,n388);
    dff g465(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1593), .Q(n3[36]));
    nand g466(n1068 ,n1905 ,n408);
    not g467(n1398 ,n1371);
    not g468(n1542 ,n1500);
    nand g469(n1004 ,n1879 ,n405);
    nand g470(n810 ,n3[40] ,n621);
    nand g471(n1195 ,n5[31] ,n732);
    xnor g472(n1915 ,n1983 ,n358);
    nand g473(n1132 ,n5[58] ,n732);
    nand g474(n333 ,n1966 ,n332);
    dff g475(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1435), .Q(n5[39]));
    nand g476(n1488 ,n1033 ,n1024);
    nor g477(n252 ,n34 ,n251);
    nand g478(n1728 ,n2026 ,n1666);
    nand g479(n1114 ,n697 ,n698);
    nand g480(n2131 ,n4[26] ,n2128);
    dff g481(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n541), .Q(n9[27]));
    nand g482(n608 ,n486 ,n607);
    nand g483(n1864 ,n2195 ,n2194);
    nand g484(n1448 ,n1201 ,n1200);
    dff g485(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1575), .Q(n3[50]));
    nand g486(n2202 ,n4[61] ,n2198);
    not g487(n1528 ,n1478);
    nor g488(n529 ,n475 ,n1);
    nand g489(n654 ,n4[60] ,n402);
    nand g490(n1816 ,n2099 ,n2098);
    or g491(n646 ,n1 ,n627);
    nor g492(n249 ,n94 ,n248);
    nand g493(n1627 ,n853 ,n1400);
    dff g494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1565), .Q(n3[60]));
    nand g495(n1775 ,n1669 ,n3[7]);
    not g496(n734 ,n733);
    not g497(n469 ,n2[41]);
    nor g498(n1297 ,n487 ,n1027);
    nand g499(n1965 ,n1725 ,n1722);
    not g500(n332 ,n331);
    nand g501(n738 ,n2[89] ,n629);
    xnor g502(n137 ,n2[6] ,n2[70]);
    nand g503(n1821 ,n2109 ,n2108);
    nand g504(n1050 ,n1912 ,n729);
    nand g505(n1175 ,n759 ,n743);
    dff g506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1424), .Q(n5[50]));
    nand g507(n1186 ,n663 ,n658);
    or g508(n2188 ,n4[55] ,n2186);
    nor g509(n162 ,n32 ,n161);
    nor g510(n510 ,n454 ,n1);
    not g511(n316 ,n315);
    nand g512(n981 ,n1884 ,n405);
    nand g513(n938 ,n1816 ,n409);
    nand g514(n325 ,n1962 ,n324);
    nor g515(n39 ,n2[39] ,n2[103]);
    nand g516(n787 ,n3[56] ,n398);
    nand g517(n1147 ,n728 ,n649);
    dff g518(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n528), .Q(n9[16]));
    nand g519(n2236 ,n11[15] ,n2219);
    xnor g520(n1884 ,n1952 ,n305);
    nand g521(n1001 ,n1927 ,n408);
    nand g522(n1785 ,n2008 ,n1666);
    not g523(n447 ,n2[62]);
    xnor g524(n1896 ,n1964 ,n327);
    nand g525(n1460 ,n1213 ,n974);
    xnor g526(n2067 ,n8[2] ,n394);
    dff g527(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1340), .Q(n4[26]));
    dff g528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1623), .Q(n3[13]));
    nand g529(n1863 ,n2193 ,n2192);
    not g530(n338 ,n337);
    nand g531(n1829 ,n2125 ,n2124);
    not g532(n430 ,n2[50]);
    not g533(n318 ,n317);
    nand g534(n594 ,n2[64] ,n6[0]);
    nor g535(n143 ,n100 ,n142);
    nand g536(n1228 ,n1919 ,n408);
    nand g537(n1777 ,n2034 ,n1666);
    nand g538(n673 ,n4[8] ,n620);
    nand g539(n1369 ,n653 ,n843);
    xnor g540(n2007 ,n111 ,n154);
    nand g541(n1414 ,n832 ,n1091);
    nand g542(n1770 ,n2004 ,n1666);
    or g543(n2148 ,n4[35] ,n2146);
    nor g544(n731 ,n1 ,n624);
    not g545(n476 ,n2[48]);
    nand g546(n1355 ,n936 ,n1281);
    nor g547(n18 ,n2[48] ,n2[112]);
    nand g548(n963 ,n1806 ,n410);
    not g549(n1653 ,n1645);
    nand g550(n1956 ,n1689 ,n1688);
    nand g551(n614 ,n544 ,n611);
    nor g552(n256 ,n72 ,n255);
    dff g553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1301), .Q(n4[62]));
    xnor g554(n1882 ,n1950 ,n301);
    nand g555(n1091 ,n2[25] ,n403);
    nand g556(n880 ,n1876 ,n408);
    xnor g557(n1892 ,n1960 ,n319);
    nand g558(n916 ,n1834 ,n409);
    nor g559(n190 ,n61 ,n189);
    nand g560(n876 ,n2[7] ,n730);
    xnor g561(n1808 ,n2079 ,n2082);
    nand g562(n1208 ,n5[24] ,n400);
    nand g563(n1354 ,n927 ,n1280);
    nand g564(n919 ,n1920 ,n731);
    xor g565(n1868 ,n4[62] ,n2200);
    nand g566(n2155 ,n4[38] ,n2152);
    nand g567(n962 ,n1896 ,n405);
    nand g568(n1938 ,n1784 ,n1802);
    or g569(n2196 ,n4[59] ,n2194);
    nand g570(n1063 ,n1907 ,n408);
    nor g571(n180 ,n55 ,n179);
    xnor g572(n2034 ,n109 ,n208);
    nand g573(n977 ,n1887 ,n731);
    not g574(n1231 ,n1100);
    not g575(n1287 ,n1188);
    nand g576(n1610 ,n909 ,n1339);
    nand g577(n1952 ,n1673 ,n1672);
    nand g578(n830 ,n4[39] ,n620);
    nand g579(n1439 ,n1190 ,n947);
    dff g580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1477), .Q(n5[9]));
    nand g581(n862 ,n2[13] ,n730);
    nand g582(n1464 ,n778 ,n982);
    nor g583(n210 ,n36 ,n209);
    nand g584(n1490 ,n794 ,n1034);
    nand g585(n841 ,n2[22] ,n730);
    nand g586(n655 ,n3[20] ,n621);
    not g587(n1534 ,n1489);
    or g588(n2170 ,n4[46] ,n2168);
    nand g589(n710 ,n2[104] ,n629);
    nand g590(n1513 ,n825 ,n1081);
    nand g591(n1984 ,n1730 ,n1727);
    nand g592(n1335 ,n864 ,n1262);
    not g593(n373 ,n372);
    nor g594(n543 ,n2[2] ,n6[2]);
    nand g595(n1734 ,n1669 ,n3[29]);
    nand g596(n299 ,n1948 ,n298);
    nor g597(n150 ,n24 ,n149);
    nand g598(n1202 ,n5[28] ,n732);
    or g599(n2178 ,n4[50] ,n2176);
    nand g600(n1795 ,n1668 ,n3[51]);
    not g601(n1261 ,n1142);
    nand g602(n997 ,n1880 ,n405);
    dff g603(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n530), .Q(n9[22]));
    nand g604(n1607 ,n1106 ,n1388);
    nor g605(n567 ,n465 ,n1);
    not g606(n454 ,n2[30]);
    dff g607(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1659), .Q(n5[3]));
    nor g608(n576 ,n421 ,n1);
    not g609(n1286 ,n1186);
    dff g610(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1327), .Q(n4[37]));
    nand g611(n323 ,n1961 ,n322);
    nand g612(n687 ,n4[50] ,n402);
    nand g613(n347 ,n1974 ,n341);
    nand g614(n1583 ,n1044 ,n1539);
    nand g615(n1742 ,n2029 ,n1665);
    not g616(n1666 ,n1664);
    nand g617(n742 ,n2[87] ,n629);
    nand g618(n970 ,n1892 ,n731);
    xnor g619(n125 ,n2[17] ,n2[81]);
    nand g620(n1426 ,n1155 ,n1048);
    nor g621(n12 ,n2[47] ,n2[111]);
    nor g622(n523 ,n463 ,n1);
    not g623(n545 ,n544);
    not g624(n328 ,n327);
    nand g625(n833 ,n4[34] ,n402);
    nand g626(n2235 ,n9[16] ,n2221);
    nand g627(n1689 ,n1668 ,n3[18]);
    xor g628(n1908 ,n1976 ,n345);
    xnor g629(n2079 ,n6[2] ,n4[2]);
    nor g630(n530 ,n422 ,n1);
    not g631(n1239 ,n1109);
    nand g632(n2241 ,n9[25] ,n2214);
    nand g633(n1477 ,n1223 ,n1004);
    not g634(n2071 ,n6[0]);
    dff g635(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1446), .Q(n5[30]));
    nand g636(n1162 ,n750 ,n716);
    nand g637(n1107 ,n746 ,n718);
    not g638(n436 ,n2[75]);
    nand g639(n768 ,n4[5] ,n402);
    nor g640(n244 ,n59 ,n243);
    nand g641(n902 ,n1850 ,n410);
    nand g642(n1425 ,n1150 ,n920);
    nand g643(n1349 ,n969 ,n1275);
    nand g644(n2095 ,n4[8] ,n2092);
    or g645(n2136 ,n4[29] ,n2134);
    not g646(n412 ,n629);
    nand g647(n984 ,n1924 ,n731);
    xnor g648(n1900 ,n1968 ,n335);
    buf g649(n7[1] ,n1662);
    nand g650(n695 ,n4[51] ,n620);
    nand g651(n908 ,n1929 ,n731);
    nand g652(n1168 ,n753 ,n773);
    xnor g653(n131 ,n2[20] ,n2[84]);
    dff g654(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n518), .Q(n8[1]));
    dff g655(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1634), .Q(n3[24]));
    dff g656(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1483), .Q(n5[5]));
    nand g657(n1778 ,n2006 ,n1666);
    nand g658(n1353 ,n931 ,n1279);
    or g659(n267 ,n1940 ,n1936);
    nor g660(n229 ,n77 ,n228);
    nand g661(n2127 ,n4[24] ,n2124);
    not g662(n446 ,n2[33]);
    nor g663(n730 ,n1 ,n630);
    not g664(n1254 ,n1129);
    nand g665(n667 ,n3[11] ,n398);
    nand g666(n686 ,n2[120] ,n406);
    nand g667(n999 ,n2[57] ,n730);
    nand g668(n1083 ,n1837 ,n729);
    nand g669(n1358 ,n940 ,n1284);
    xnor g670(n2031 ,n98 ,n202);
    nor g671(n2239 ,n2205 ,n11[16]);
    nor g672(n536 ,n484 ,n1);
    nand g673(n1858 ,n2183 ,n2182);
    not g674(n1275 ,n1166);
    xnor g675(n2049 ,n118 ,n238);
    nand g676(n1037 ,n2[47] ,n730);
    xnor g677(n2046 ,n107 ,n232);
    xor g678(n1880 ,n1948 ,n298);
    nor g679(n632 ,n485 ,n618);
    nand g680(n1505 ,n814 ,n1061);
    nand g681(n1789 ,n1668 ,n3[11]);
    dff g682(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1597), .Q(n3[32]));
    nor g683(n58 ,n2[22] ,n2[86]);
    nand g684(n1594 ,n1068 ,n1548);
    nor g685(n165 ,n120 ,n164);
    nand g686(n1759 ,n1669 ,n3[3]);
    dff g687(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1458), .Q(n5[20]));
    not g688(n426 ,n2[93]);
    nand g689(n1203 ,n5[27] ,n400);
    dff g690(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1518), .Q(n5[60]));
    xnor g691(n127 ,n2[41] ,n2[105]);
    dff g692(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n4[11]));
    nand g693(n1515 ,n828 ,n1087);
    nand g694(n2117 ,n4[19] ,n2114);
    nor g695(n559 ,n414 ,n1);
    nand g696(n1483 ,n1227 ,n1019);
    nand g697(n1791 ,n2036 ,n1666);
    nand g698(n826 ,n3[54] ,n398);
    nand g699(n728 ,n2[92] ,n406);
    nor g700(n21 ,n2[40] ,n2[104]);
    nand g701(n1609 ,n1177 ,n1389);
    nand g702(n1005 ,n1878 ,n731);
    dff g703(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1661), .Q(n5[2]));
    nor g704(n160 ,n65 ,n159);
    dff g705(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n572), .Q(n11[12]));
    nand g706(n1969 ,n1743 ,n1742);
    nand g707(n1793 ,n1668 ,n3[12]);
    nand g708(n2077 ,n6[1] ,n2069);
    not g709(n1248 ,n1119);
    nand g710(n887 ,n1873 ,n410);
    nand g711(n1333 ,n1083 ,n1261);
    nor g712(n570 ,n432 ,n1);
    nand g713(n949 ,n1810 ,n409);
    nand g714(n1019 ,n1875 ,n731);
    not g715(n1241 ,n1111);
    dff g716(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1422), .Q(n5[51]));
    xnor g717(n2066 ,n8[3] ,n396);
    nor g718(n555 ,n436 ,n1);
    not g719(n411 ,n1663);
    nand g720(n1321 ,n942 ,n1249);
    xnor g721(n1886 ,n1954 ,n309);
    nand g722(n987 ,n1932 ,n409);
    nand g723(n1718 ,n1669 ,n3[59]);
    nand g724(n793 ,n3[49] ,n621);
    nor g725(n239 ,n118 ,n238);
    or g726(n2108 ,n4[15] ,n2106);
    dff g727(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1443), .Q(n5[32]));
    nand g728(n1570 ,n1008 ,n1528);
    or g729(n2150 ,n4[36] ,n2148);
    dff g730(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1463), .Q(n5[15]));
    nand g731(n831 ,n3[26] ,n621);
    nand g732(n955 ,n1808 ,n410);
    not g733(n1548 ,n1507);
    xor g734(n1806 ,n6[0] ,n4[0]);
    not g735(n1519 ,n1414);
    nor g736(n34 ,n2[57] ,n2[121]);
    dff g737(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1317), .Q(n4[47]));
    nor g738(n1296 ,n411 ,n1028);
    nor g739(n148 ,n23 ,n147);
    nor g740(n2263 ,n2249 ,n2233);
    nor g741(n167 ,n122 ,n166);
    nand g742(n2246 ,n9[22] ,n2204);
    nand g743(n1840 ,n2147 ,n2146);
    nand g744(n2248 ,n9[3] ,n9[2]);
    nand g745(n900 ,n1852 ,n409);
    nand g746(n888 ,n1815 ,n408);
    not g747(n467 ,n2[55]);
    xnor g748(n2011 ,n119 ,n162);
    not g749(n1282 ,n1179);
    nand g750(n657 ,n3[17] ,n621);
    not g751(n424 ,n2[34]);
    nand g752(n1559 ,n877 ,n1410);
    not g753(n410 ,n407);
    nand g754(n1222 ,n5[10] ,n400);
    nand g755(n1183 ,n765 ,n673);
    nor g756(n35 ,n2[13] ,n2[77]);
    nand g757(n1787 ,n1669 ,n3[37]);
    nand g758(n280 ,n276 ,n266);
    nand g759(n1330 ,n1025 ,n1258);
    or g760(n2198 ,n4[60] ,n2196);
    nand g761(n1827 ,n2121 ,n2120);
    nand g762(n1151 ,n737 ,n824);
    not g763(n1288 ,n1191);
    nand g764(n1140 ,n721 ,n784);
    nand g765(n2103 ,n4[12] ,n2100);
    nand g766(n1659 ,n1492 ,n1654);
    dff g767(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1642), .Q(n3[0]));
    nor g768(n33 ,n2[54] ,n2[118]);
    nand g769(n1176 ,n5[39] ,n400);
    nand g770(n1328 ,n1064 ,n1256);
    not g771(n1558 ,n1517);
    xnor g772(n2055 ,n106 ,n250);
    dff g773(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1571), .Q(n3[54]));
    dff g774(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1572), .Q(n3[53]));
    nand g775(n1996 ,n1687 ,n1675);
    nor g776(n528 ,n428 ,n1);
    dff g777(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1631), .Q(n3[21]));
    dff g778(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1420), .Q(n5[54]));
    nand g779(n1307 ,n943 ,n1235);
    nand g780(n1435 ,n1176 ,n953);
    nand g781(n2086 ,n2074 ,n2085);
    xnor g782(n1873 ,n280 ,n286);
    nand g783(n1982 ,n1713 ,n1710);
    nand g784(n1600 ,n1082 ,n1554);
    or g785(n2116 ,n4[19] ,n2114);
    nor g786(n551 ,n418 ,n1);
    nand g787(n894 ,n1860 ,n410);
    nand g788(n301 ,n1949 ,n300);
    xnor g789(n2032 ,n103 ,n204);
    nand g790(n1017 ,n2[52] ,n730);
    nor g791(n493 ,n4[2] ,n6[2]);
    nand g792(n1588 ,n598 ,n1291);
    nand g793(n765 ,n2[72] ,n406);
    not g794(n1532 ,n1486);
    not g795(n1546 ,n1505);
    nand g796(n1717 ,n2043 ,n1665);
    not g797(n457 ,n2[90]);
    nand g798(n1517 ,n735 ,n1095);
    nand g799(n1126 ,n710 ,n688);
    dff g800(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n550), .Q(n9[18]));
    not g801(n306 ,n305);
    not g802(n294 ,n293);
    not g803(n290 ,n289);
    nand g804(n1051 ,n1871 ,n731);
    nand g805(n1100 ,n680 ,n679);
    nor g806(n641 ,n499 ,n622);
    nor g807(n236 ,n25 ,n235);
    not g808(n1401 ,n1374);
    not g809(n1242 ,n1112);
    nand g810(n2082 ,n2077 ,n2081);
    nand g811(n1216 ,n5[16] ,n732);
    not g812(n1520 ,n1464);
    nand g813(n1727 ,n2044 ,n1665);
    nor g814(n152 ,n56 ,n151);
    nand g815(n1566 ,n996 ,n1524);
    nand g816(n901 ,n2[58] ,n730);
    nand g817(n1796 ,n2011 ,n1665);
    nor g818(n14 ,n2[55] ,n2[119]);
    or g819(n2144 ,n4[33] ,n2142);
    nand g820(n1772 ,n1669 ,n3[35]);
    not g821(n1550 ,n1509);
    nor g822(n63 ,n2[38] ,n2[102]);
    dff g823(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1640), .Q(n3[1]));
    nand g824(n1944 ,n1771 ,n1770);
    nand g825(n1347 ,n1000 ,n1273);
    nand g826(n871 ,n2[9] ,n403);
    nor g827(n522 ,n417 ,n1);
    dff g828(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1330), .Q(n4[34]));
    xnor g829(n2003 ,n105 ,n146);
    or g830(n2098 ,n4[10] ,n2096);
    nand g831(n1786 ,n1669 ,n3[10]);
    nand g832(n1006 ,n2[55] ,n730);
    nand g833(n276 ,n1941 ,n1937);
    nand g834(n1634 ,n1096 ,n1558);
    not g835(n2212 ,n9[6]);
    nand g836(n1845 ,n2157 ,n2156);
    or g837(n2112 ,n4[17] ,n2110);
    nand g838(n2183 ,n4[52] ,n2180);
    xor g839(n1871 ,n281 ,n275);
    dff g840(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1334), .Q(n4[56]));
    dff g841(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1562), .Q(n3[63]));
    nor g842(n26 ,n2[8] ,n2[72]);
    nand g843(n1757 ,n1669 ,n3[60]);
    nand g844(n1000 ,n1825 ,n729);
    nand g845(n1852 ,n2171 ,n2170);
    nand g846(n1182 ,n5[37] ,n732);
    nor g847(n503 ,n5[3] ,n6[3]);
    nand g848(n803 ,n2[117] ,n406);
    nand g849(n990 ,n1882 ,n405);
    dff g850(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n510), .Q(n10[30]));
    nand g851(n1624 ,n861 ,n1403);
    nand g852(n1197 ,n586 ,n633);
    xnor g853(n95 ,n2[60] ,n2[124]);
    nand g854(n1375 ,n660 ,n857);
    nor g855(n213 ,n117 ,n212);
    nor g856(n838 ,n506 ,n413);
    xnor g857(n2045 ,n82 ,n230);
    dff g858(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1627), .Q(n3[17]));
    nand g859(n1362 ,n949 ,n1288);
    not g860(n1538 ,n1494);
    nand g861(n1709 ,n2052 ,n1665);
    xnor g862(n96 ,n2[40] ,n2[104]);
    not g863(n1269 ,n1156);
    nand g864(n829 ,n4[62] ,n402);
    nand g865(n1120 ,n5[63] ,n400);
    nand g866(n582 ,n3[2] ,n6[2]);
    dff g867(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1325), .Q(n4[39]));
    nor g868(n174 ,n46 ,n173);
    not g869(n1246 ,n1117);
    nand g870(n1122 ,n727 ,n723);
    nand g871(n701 ,n4[47] ,n402);
    xnor g872(n1918 ,n1986 ,n364);
    nor g873(n151 ,n108 ,n150);
    not g874(n438 ,n2[42]);
    not g875(n1397 ,n1370);
    dff g876(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n549), .Q(n9[19]));
    nand g877(n684 ,n4[57] ,n620);
    dff g878(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1617), .Q(n3[4]));
    nand g879(n1086 ,n1898 ,n729);
    nor g880(n540 ,n426 ,n1);
    nor g881(n502 ,n3[2] ,n6[2]);
    nand g882(n1582 ,n601 ,n1290);
    nand g883(n764 ,n2[73] ,n406);
    nand g884(n809 ,n2[99] ,n629);
    nand g885(n1377 ,n662 ,n862);
    nand g886(n961 ,n1897 ,n731);
    nand g887(n886 ,n1904 ,n405);
    nor g888(n2229 ,n2217 ,n9[13]);
    nand g889(n1458 ,n1212 ,n973);
    dff g890(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n492), .Q(n8[0]));
    nor g891(n37 ,n2[51] ,n2[115]);
    nor g892(n68 ,n2[3] ,n2[67]);
    xnor g893(n2058 ,n95 ,n256);
    nor g894(n504 ,n5[2] ,n6[2]);
    nand g895(n693 ,n3[58] ,n621);
    nand g896(n1867 ,n2202 ,n2201);
    not g897(n1412 ,n1385);
    nand g898(n1106 ,n582 ,n645);
    nand g899(n1576 ,n1228 ,n1534);
    nand g900(n1828 ,n2123 ,n2122);
    dff g901(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n569), .Q(n11[15]));
    dff g902(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1430), .Q(n5[44]));
    nand g903(n1137 ,n5[56] ,n732);
    nand g904(n286 ,n270 ,n285);
    nor g905(n181 ,n135 ,n180);
    nand g906(n1722 ,n2025 ,n1665);
    nand g907(n1336 ,n859 ,n1263);
    nand g908(n1115 ,n699 ,n797);
    nor g909(n2240 ,n2206 ,n11[18]);
    nand g910(n2262 ,n2231 ,n2237);
    nor g911(n170 ,n17 ,n169);
    nand g912(n773 ,n4[16] ,n402);
    nand g913(n1940 ,n1753 ,n1804);
    nand g914(n1962 ,n1724 ,n1711);
    not g915(n1668 ,n1667);
    nand g916(n1710 ,n2042 ,n1666);
    nand g917(n985 ,n1824 ,n409);
    not g918(n441 ,n2[46]);
    or g919(n2130 ,n4[26] ,n2128);
    nor g920(n260 ,n38 ,n259);
    nand g921(n1741 ,n2058 ,n1665);
    dff g922(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1427), .Q(n5[47]));
    nand g923(n1319 ,n935 ,n1247);
    dff g924(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n540), .Q(n9[29]));
    xnor g925(n119 ,n2[13] ,n2[77]);
    dff g926(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1313), .Q(n4[50]));
    nand g927(n1621 ,n868 ,n1406);
    not g928(n1400 ,n1373);
    nand g929(n1573 ,n1018 ,n1531);
    not g930(n1274 ,n1164);
    nand g931(n605 ,n1663 ,n544);
    dff g932(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n509), .Q(n10[28]));
    xnor g933(n1878 ,n1946 ,n295);
    xnor g934(n2025 ,n80 ,n190);
    not g935(n1409 ,n1382);
    not g936(n442 ,n2[31]);
    nor g937(n70 ,n2[30] ,n2[94]);
    nand g938(n1784 ,n1668 ,n3[0]);
    nand g939(n649 ,n4[28] ,n620);
    nand g940(n1957 ,n1692 ,n1691);
    dff g941(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n560), .Q(n11[17]));
    nand g942(n1629 ,n849 ,n1398);
    nand g943(n1481 ,n1225 ,n1010);
    nand g944(n2169 ,n4[45] ,n2166);
    nand g945(n1595 ,n1071 ,n1549);
    dff g946(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1601), .Q(n3[28]));
    not g947(n1399 ,n1372);
    dff g948(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1336), .Q(n4[29]));
    not g949(n419 ,n2[69]);
    nor g950(n514 ,n423 ,n1);
    nand g951(n715 ,n4[37] ,n620);
    dff g952(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1592), .Q(n3[37]));
    xnor g953(n113 ,n2[10] ,n2[74]);
    nand g954(n1473 ,n693 ,n901);
    xnor g955(n2038 ,n96 ,n216);
    nand g956(n1312 ,n896 ,n1241);
    dff g957(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1598), .Q(n3[30]));
    dff g958(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1594), .Q(n3[35]));
    not g959(n458 ,n2[78]);
    nand g960(n874 ,n2[8] ,n403);
    nand g961(n1672 ,n2012 ,n1665);
    not g962(n421 ,n2[59]);
    nand g963(n943 ,n1863 ,n409);
    not g964(n324 ,n323);
    nand g965(n1227 ,n5[5] ,n400);
    nor g966(n531 ,n439 ,n1);
    nand g967(n1368 ,n652 ,n841);
    nor g968(n186 ,n40 ,n185);
    xnor g969(n80 ,n2[27] ,n2[91]);
    nand g970(n1116 ,n700 ,n701);
    nor g971(n187 ,n88 ,n186);
    nor g972(n617 ,n1662 ,n610);
    dff g973(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1454), .Q(n5[24]));
    nand g974(n983 ,n1933 ,n409);
    nand g975(n1046 ,n2[43] ,n730);
    nand g976(n2133 ,n4[27] ,n2130);
    dff g977(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n570), .Q(n11[26]));
    nand g978(n1846 ,n2159 ,n2158);
    nand g979(n718 ,n4[55] ,n402);
    nand g980(n704 ,n4[45] ,n620);
    nand g981(n1097 ,n592 ,n648);
    nor g982(n526 ,n450 ,n1);
    not g983(n1268 ,n1153);
    not g984(n1277 ,n1170);
    dff g985(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n554), .Q(n9[13]));
    nand g986(n1471 ,n783 ,n995);
    dff g987(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n516), .Q(n11[10]));
    nor g988(n245 ,n86 ,n244);
    xnor g989(n123 ,n2[58] ,n2[122]);
    nand g990(n1824 ,n2115 ,n2114);
    nand g991(n1614 ,n955 ,n1364);
    xnor g992(n2016 ,n128 ,n172);
    nand g993(n986 ,n2[62] ,n403);
    nand g994(n335 ,n1967 ,n334);
    nand g995(n1615 ,n959 ,n1365);
    nand g996(n1310 ,n899 ,n1239);
    dff g997(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1308), .Q(n4[55]));
    nand g998(n1475 ,n786 ,n999);
    not g999(n486 ,n1662);
    dff g1000(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1350), .Q(n4[16]));
    dff g1001(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1652), .Q(n4[1]));
    nand g1002(n1014 ,n1827 ,n408);
    not g1003(n1284 ,n1183);
    nand g1004(n925 ,n1902 ,n731);
    nand g1005(n1754 ,n2031 ,n1666);
    nand g1006(n1118 ,n705 ,n704);
    not g1007(n463 ,n2[71]);
    nand g1008(n1141 ,n5[54] ,n400);
    nor g1009(n581 ,n462 ,n1);
    not g1010(n302 ,n301);
    nand g1011(n1939 ,n1748 ,n1803);
    or g1012(n2154 ,n4[38] ,n2152);
    xnor g1013(n2020 ,n135 ,n180);
    nand g1014(n807 ,n4[23] ,n402);
    nor g1015(n645 ,n502 ,n622);
    xnor g1016(n2040 ,n132 ,n220);
    not g1017(n1544 ,n1503);
    xnor g1018(n1876 ,n1944 ,n291);
    nand g1019(n808 ,n3[41] ,n398);
    nand g1020(n337 ,n1968 ,n336);
    nand g1021(n845 ,n2[20] ,n730);
    nand g1022(n672 ,n3[7] ,n621);
    nand g1023(n1343 ,n1056 ,n1269);
    nand g1024(n1042 ,n1915 ,n729);
    not g1025(n359 ,n358);
    nor g1026(n176 ,n48 ,n175);
    not g1027(n402 ,n401);
    dff g1028(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1618), .Q(n3[8]));
    xor g1029(n2063 ,n97 ,n140);
    nand g1030(n1843 ,n2153 ,n2152);
    nand g1031(n1510 ,n821 ,n1075);
    xnor g1032(n6[3] ,n10[31] ,n2284);
    not g1033(n383 ,n382);
    not g1034(n1531 ,n1484);
    nand g1035(n2167 ,n4[44] ,n2164);
    nand g1036(n1493 ,n798 ,n1039);
    nand g1037(n1219 ,n5[13] ,n732);
    nand g1038(n1052 ,n2[41] ,n403);
    nand g1039(n910 ,n1841 ,n410);
    xor g1040(n1870 ,n1934 ,n1938);
    nor g1041(n633 ,n493 ,n622);
    nor g1042(n36 ,n2[36] ,n2[100]);
    nand g1043(n883 ,n2[4] ,n403);
    nor g1044(n556 ,n466 ,n1);
    nor g1045(n568 ,n480 ,n1);
    nand g1046(n1811 ,n2089 ,n2088);
    or g1047(n2223 ,n9[1] ,n9[0]);
    xnor g1048(n1902 ,n339 ,n1970);
    nor g1049(n23 ,n2[5] ,n2[69]);
    xnor g1050(n2051 ,n129 ,n242);
    nand g1051(n1995 ,n1779 ,n1768);
    nand g1052(n714 ,n2[101] ,n406);
    nand g1053(n1440 ,n1187 ,n944);
    nand g1054(n767 ,n2[69] ,n629);
    nand g1055(n1111 ,n694 ,n695);
    nand g1056(n922 ,n1917 ,n731);
    not g1057(n483 ,n2067);
    dff g1058(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1626), .Q(n3[16]));
    nand g1059(n659 ,n3[16] ,n621);
    nand g1060(n2173 ,n4[47] ,n2170);
    nand g1061(n279 ,n270 ,n267);
    nand g1062(n818 ,n3[34] ,n621);
    xnor g1063(n2009 ,n115 ,n158);
    dff g1064(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n603), .Q(n9[23]));
    dff g1065(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1312), .Q(n4[51]));
    dff g1066(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n565), .Q(n11[2]));
    nand g1067(n1172 ,n756 ,n774);
    nand g1068(n1630 ,n846 ,n1397);
    nand g1069(n596 ,n3[1] ,n6[1]);
    nand g1070(n283 ,n1972 ,n282);
    nand g1071(n1853 ,n2173 ,n2172);
    dff g1072(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1344), .Q(n4[22]));
    dff g1073(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n580), .Q(n11[22]));
    nand g1074(n583 ,n2[2] ,n6[2]);
    nand g1075(n1830 ,n2127 ,n2126);
    nand g1076(n849 ,n1889 ,n729);
    nand g1077(n995 ,n2[59] ,n730);
    nor g1078(n2231 ,n2213 ,n11[28]);
    xnor g1079(n2057 ,n101 ,n254);
    nor g1080(n242 ,n45 ,n241);
    dff g1081(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n517), .Q(n11[6]));
    nor g1082(n2281 ,n2276 ,n2274);
    not g1083(n1552 ,n1511);
    nand g1084(n781 ,n3[61] ,n621);
    nand g1085(n769 ,n2[68] ,n629);
    xnor g1086(n2010 ,n116 ,n160);
    not g1087(n1936 ,n1737);
    nand g1088(n1346 ,n924 ,n1272);
    nand g1089(n348 ,n1976 ,n345);
    nand g1090(n737 ,n2[90] ,n629);
    nor g1091(n19 ,n2[15] ,n2[79]);
    nand g1092(n1766 ,n2003 ,n1666);
    nand g1093(n1455 ,n1209 ,n968);
    nand g1094(n1334 ,n893 ,n1236);
    nand g1095(n372 ,n1990 ,n371);
    nor g1096(n509 ,n449 ,n1);
    nor g1097(n563 ,n437 ,n1);
    nand g1098(n1494 ,n800 ,n1041);
    nor g1099(n518 ,n482 ,n1);
    nand g1100(n2250 ,n9[27] ,n9[26]);
    nand g1101(n1171 ,n5[41] ,n732);
    nand g1102(n1008 ,n1925 ,n408);
    nand g1103(n939 ,n1907 ,n405);
    not g1104(n1547 ,n1506);
    nand g1105(n1586 ,n1050 ,n1541);
    dff g1106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1465), .Q(n5[14]));
    nand g1107(n843 ,n2[21] ,n403);
    or g1108(n2184 ,n4[53] ,n2182);
    nand g1109(n1958 ,n1744 ,n1696);
    nand g1110(n1110 ,n692 ,n689);
    nor g1111(n520 ,n415 ,n1);
    not g1112(n1407 ,n1380);
    nand g1113(n1950 ,n1793 ,n1792);
    nand g1114(n794 ,n3[48] ,n621);
    not g1115(n485 ,n7[0]);
    nand g1116(n1763 ,n1669 ,n3[40]);
    dff g1117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1337), .Q(n4[28]));
    nand g1118(n2177 ,n4[49] ,n2174);
    nand g1119(n1841 ,n2149 ,n2148);
    nand g1120(n1833 ,n2133 ,n2132);
    nand g1121(n941 ,n1906 ,n731);
    nand g1122(n1373 ,n657 ,n852);
    nor g1123(n494 ,n2[1] ,n6[1]);
    not g1124(n2219 ,n11[14]);
    nor g1125(n515 ,n473 ,n1);
    xnor g1126(n88 ,n2[25] ,n2[89]);
    nand g1127(n344 ,n1970 ,n340);
    dff g1128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1566), .Q(n3[59]));
    not g1129(n1240 ,n1110);
    nand g1130(n2101 ,n4[11] ,n2098);
    not g1131(n453 ,n2[74]);
    nor g1132(n55 ,n2[21] ,n2[85]);
    nand g1133(n1866 ,n2199 ,n2198);
    nand g1134(n1677 ,n1668 ,n3[15]);
    dff g1135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1441), .Q(n5[34]));
    nand g1136(n2258 ,n2240 ,n2239);
    nand g1137(n1994 ,n1755 ,n1745);
    not g1138(n2073 ,n4[4]);
    nand g1139(n820 ,n4[27] ,n402);
    nand g1140(n827 ,n3[28] ,n621);
    nor g1141(n1638 ,n1 ,n1637);
    xnor g1142(n104 ,n2[16] ,n2[80]);
    nand g1143(n682 ,n2[123] ,n406);
    nand g1144(n1589 ,n1055 ,n1543);
    dff g1145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1289), .Q(n5[61]));
    nand g1146(n696 ,n2[114] ,n629);
    nand g1147(n1713 ,n1668 ,n3[44]);
    nor g1148(n194 ,n50 ,n193);
    nand g1149(n1007 ,n1916 ,n731);
    not g1150(n1271 ,n1159);
    not g1151(n2214 ,n9[24]);
    nor g1152(n185 ,n87 ,n184);
    xnor g1153(n2037 ,n121 ,n214);
    nor g1154(n1637 ,n1295 ,n1293);
    nand g1155(n1738 ,n2028 ,n1665);
    nand g1156(n1604 ,n1094 ,n1519);
    nand g1157(n2189 ,n4[55] ,n2186);
    not g1158(n1529 ,n1480);
    nand g1159(n951 ,n1821 ,n409);
    not g1160(n1530 ,n1482);
    nor g1161(n564 ,n461 ,n1);
    nand g1162(n1437 ,n1182 ,n939);
    nand g1163(n376 ,n1992 ,n375);
    nor g1164(n2224 ,n11[1] ,n11[0]);
    nor g1165(n341 ,n283 ,n339);
    nor g1166(n579 ,n444 ,n1);
    nand g1167(n988 ,n1883 ,n731);
    nand g1168(n362 ,n1984 ,n361);
    nand g1169(n2238 ,n11[13] ,n11[12]);
    xnor g1170(n76 ,n2[29] ,n2[93]);
    nor g1171(n2076 ,n2071 ,n4[0]);
    nand g1172(n1451 ,n1205 ,n1204);
    xnor g1173(n138 ,n2[23] ,n2[87]);
    nand g1174(n1476 ,n787 ,n1002);
    xnor g1175(n2048 ,n110 ,n236);
    nand g1176(n1386 ,n676 ,n883);
    nand g1177(n1966 ,n1729 ,n1728);
    nand g1178(n791 ,n3[51] ,n621);
    xnor g1179(n1893 ,n1961 ,n321);
    nand g1180(n1135 ,n809 ,n719);
    xnor g1181(n2015 ,n125 ,n170);
    nand g1182(n927 ,n1818 ,n410);
    nand g1183(n1098 ,n677 ,n651);
    nand g1184(n2273 ,n2266 ,n2254);
    nor g1185(n28 ,n2[42] ,n2[106]);
    nand g1186(n1495 ,n802 ,n1043);
    xnor g1187(n134 ,n2[55] ,n2[119]);
    not g1188(n1257 ,n1135);
    not g1189(n1669 ,n1667);
    xnor g1190(n1911 ,n353 ,n1979);
    nand g1191(n822 ,n3[31] ,n621);
    nand g1192(n1673 ,n1668 ,n3[14]);
    dff g1193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1450), .Q(n5[27]));
    nand g1194(n1043 ,n2[44] ,n730);
    not g1195(n2213 ,n11[29]);
    nand g1196(n1760 ,n2032 ,n1665);
    nand g1197(n1143 ,n724 ,n670);
    not g1198(n1280 ,n1175);
    nand g1199(n724 ,n2[94] ,n629);
    nand g1200(n921 ,n1830 ,n409);
    nand g1201(n270 ,n1940 ,n1936);
    nand g1202(n1193 ,n5[32] ,n400);
    dff g1203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1563), .Q(n3[62]));
    nand g1204(n1650 ,n1045 ,n1582);
    xnor g1205(n132 ,n2[42] ,n2[106]);
    nand g1206(n1062 ,n1831 ,n729);
    nand g1207(n1383 ,n672 ,n876);
    dff g1208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1462), .Q(n5[16]));
    xnor g1209(n1881 ,n1949 ,n299);
    nand g1210(n1518 ,n1127 ,n964);
    nand g1211(n870 ,n1880 ,n409);
    nand g1212(n1301 ,n889 ,n1230);
    nand g1213(n588 ,n2[67] ,n6[3]);
    nand g1214(n303 ,n1950 ,n302);
    dff g1215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n523), .Q(n9[7]));
    nand g1216(n1679 ,n2038 ,n1666);
    nand g1217(n759 ,n2[76] ,n406);
    nand g1218(n327 ,n1963 ,n326);
    nand g1219(n1836 ,n2139 ,n2138);
    xnor g1220(n2008 ,n113 ,n156);
    nand g1221(n1469 ,n782 ,n992);
    dff g1222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1418), .Q(n5[56]));
    nand g1223(n676 ,n3[4] ,n398);
    nand g1224(n1979 ,n1690 ,n1686);
    nand g1225(n1113 ,n599 ,n634);
    nand g1226(n1491 ,n796 ,n1037);
    nand g1227(n356 ,n1981 ,n355);
    nand g1228(n374 ,n1991 ,n373);
    xnor g1229(n2013 ,n122 ,n166);
    not g1230(n444 ,n2[52]);
    nand g1231(n700 ,n2[111] ,n406);
    nor g1232(n230 ,n57 ,n229);
    or g1233(n2124 ,n4[23] ,n2122);
    nand g1234(n813 ,n3[38] ,n398);
    xnor g1235(n2062 ,n100 ,n142);
    nand g1236(n896 ,n1857 ,n409);
    nor g1237(n215 ,n121 ,n214);
    or g1238(n2174 ,n4[48] ,n2172);
    nand g1239(n982 ,n2[63] ,n403);
    nand g1240(n1139 ,n5[55] ,n400);
    nand g1241(n1711 ,n2022 ,n1666);
    nand g1242(n354 ,n1980 ,n352);
    nor g1243(n172 ,n42 ,n171);
    nand g1244(n722 ,n2[95] ,n629);
    xnor g1245(n2047 ,n99 ,n234);
    nor g1246(n15 ,n2[23] ,n2[87]);
    nor g1247(n393 ,n8[1] ,n8[0]);
    nand g1248(n1961 ,n1708 ,n1707);
    nand g1249(n968 ,n1893 ,n731);
    nand g1250(n1804 ,n1665 ,n1800);
    dff g1251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n4[9]));
    nand g1252(n1417 ,n1134 ,n911);
    nand g1253(n2143 ,n4[32] ,n2140);
    nand g1254(n697 ,n2[113] ,n629);
    nand g1255(n996 ,n1929 ,n410);
    nand g1256(n1592 ,n1063 ,n1546);
    nand g1257(n1971 ,n1756 ,n1754);
    nand g1258(n1758 ,n2047 ,n1666);
    nand g1259(n1612 ,n1113 ,n1390);
    nor g1260(n2278 ,n2272 ,n2270);
    nand g1261(n2093 ,n4[7] ,n2090);
    nand g1262(n1359 ,n875 ,n1285);
    nor g1263(n48 ,n2[19] ,n2[83]);
    dff g1264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n534), .Q(n11[30]));
    not g1265(n425 ,n2[38]);
    nor g1266(n60 ,n2[43] ,n2[107]);
    not g1267(n437 ,n2[36]);
    dff g1268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1619), .Q(n3[9]));
    dff g1269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n527), .Q(n9[10]));
    xor g1270(n1799 ,n2064 ,n6[1]);
    nand g1271(n1341 ,n1062 ,n1267);
    not g1272(n448 ,n2[29]);
    not g1273(n1283 ,n1181);
    nand g1274(n1032 ,n605 ,n646);
    nand g1275(n1622 ,n866 ,n1405);
    nand g1276(n1101 ,n681 ,n654);
    not g1277(n1526 ,n1475);
    xnor g1278(n81 ,n2[30] ,n2[94]);
    nand g1279(n1485 ,n1226 ,n1084);
    not g1280(n475 ,n2[79]);
    nand g1281(n1855 ,n2177 ,n2176);
    nand g1282(n1078 ,n1928 ,n731);
    not g1283(n387 ,n386);
    nand g1284(n1575 ,n1023 ,n1533);
    nand g1285(n1577 ,n1035 ,n1535);
    nand g1286(n1136 ,n801 ,n833);
    nand g1287(n935 ,n1851 ,n409);
    xnor g1288(n105 ,n2[5] ,n2[69]);
    dff g1289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1359), .Q(n4[7]));
    nand g1290(n776 ,n4[18] ,n402);
    nor g1291(n345 ,n265 ,n342);
    not g1292(n420 ,n2[63]);
    not g1293(n2206 ,n11[19]);
    xnor g1294(n2039 ,n127 ,n218);
    nand g1295(n947 ,n1903 ,n405);
    nand g1296(n307 ,n1952 ,n306);
    xnor g1297(n128 ,n2[18] ,n2[82]);
    nand g1298(n1508 ,n818 ,n1070);
    xor g1299(n1904 ,n1972 ,n343);
    xnor g1300(n82 ,n2[47] ,n2[111]);
    dff g1301(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n531), .Q(n9[20]));
    xnor g1302(n1913 ,n1981 ,n354);
    or g1303(n1640 ,n1610 ,n1609);
    not g1304(n1665 ,n1664);
    nand g1305(n782 ,n3[60] ,n621);
    nand g1306(n780 ,n4[56] ,n402);
    nand g1307(n1678 ,n2050 ,n1665);
    not g1308(n422 ,n2[86]);
    nor g1309(n226 ,n54 ,n225);
    not g1310(n334 ,n333);
    nor g1311(n155 ,n111 ,n154);
    nand g1312(n1565 ,n993 ,n1523);
    nor g1313(n557 ,n443 ,n1);
    nand g1314(n1511 ,n822 ,n1076);
    not g1315(n1267 ,n1152);
    nand g1316(n1748 ,n1668 ,n3[1]);
    nand g1317(n1694 ,n1669 ,n3[36]);
    nor g1318(n254 ,n53 ,n253);
    nand g1319(n748 ,n4[43] ,n402);
    nand g1320(n889 ,n1868 ,n410);
    nor g1321(n241 ,n124 ,n240);
    nand g1322(n1433 ,n1171 ,n933);
    dff g1323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n579), .Q(n11[20]));
    not g1324(n1258 ,n1136);
    nor g1325(n2256 ,n2234 ,n2232);
    not g1326(n1245 ,n1116);
    nand g1327(n1099 ,n678 ,n829);
    dff g1328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n535), .Q(n9[30]));
    nand g1329(n1865 ,n2197 ,n2196);
    nand g1330(n1156 ,n742 ,n807);
    not g1331(n1935 ,n1769);
    not g1332(n472 ,n2[45]);
    or g1333(n2140 ,n4[31] ,n2138);
    nand g1334(n1695 ,n2040 ,n1666);
    nand g1335(n1084 ,n1876 ,n731);
    nand g1336(n1188 ,n767 ,n768);
    not g1337(n460 ,n2[44]);
    nand g1338(n1503 ,n811 ,n1057);
    nand g1339(n1441 ,n1189 ,n886);
    nand g1340(n2157 ,n4[39] ,n2154);
    nand g1341(n964 ,n1930 ,n405);
    nor g1342(n2259 ,n2243 ,n2242);
    nand g1343(n590 ,n2[66] ,n6[2]);
    dff g1344(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1620), .Q(n3[10]));
    dff g1345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1338), .Q(n4[27]));
    nor g1346(n613 ,n7[0] ,n608);
    nand g1347(n953 ,n1909 ,n731);
    nand g1348(n763 ,n4[9] ,n620);
    nand g1349(n1701 ,n2061 ,n1665);
    dff g1350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n520), .Q(n9[2]));
    nand g1351(n1680 ,n2014 ,n1665);
    nor g1352(n31 ,n2[37] ,n2[101]);
    dff g1353(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1341), .Q(n4[25]));
    nand g1354(n1079 ,n2[30] ,n730);
    nor g1355(n65 ,n2[11] ,n2[75]);
    or g1356(n2146 ,n4[34] ,n2144);
    dff g1357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n558), .Q(n9[5]));
    nand g1358(n1826 ,n2119 ,n2118);
    nand g1359(n878 ,n1844 ,n409);
    nand g1360(n1731 ,n1669 ,n3[55]);
    nand g1361(n1831 ,n2129 ,n2128);
    dff g1362(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1326), .Q(n4[38]));
    nor g1363(n27 ,n2[45] ,n2[109]);
    not g1364(n1527 ,n1476);
    or g1365(n1643 ,n1613 ,n1442);
    nand g1366(n1797 ,n1669 ,n3[49]);
    dff g1367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1440), .Q(n5[35]));
    nand g1368(n936 ,n1817 ,n729);
    or g1369(n2284 ,n2283 ,n2282);
    nand g1370(n2234 ,n9[7] ,n2212);
    nand g1371(n670 ,n4[30] ,n620);
    nand g1372(n881 ,n2[5] ,n403);
    or g1373(n141 ,n97 ,n140);
    nand g1374(n798 ,n3[46] ,n621);
    nand g1375(n1128 ,n711 ,n830);
    not g1376(n1230 ,n1099);
    nand g1377(n1815 ,n2097 ,n2096);
    nand g1378(n1752 ,n1669 ,n3[63]);
    xnor g1379(n606 ,n486 ,n485);
    nor g1380(n534 ,n447 ,n1);
    dff g1381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1331), .Q(n4[33]));
    xnor g1382(n1925 ,n1993 ,n376);
    nand g1383(n1737 ,n6[2] ,n1669);
    nor g1384(n216 ,n39 ,n215);
    nor g1385(n171 ,n125 ,n170);
    not g1386(n484 ,n2066);
    nor g1387(n202 ,n44 ,n201);
    or g1388(n2122 ,n4[22] ,n2120);
    nand g1389(n1628 ,n851 ,n1399);
    dff g1390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1648), .Q(n7[0]));
    nand g1391(n1392 ,n1123 ,n903);
    nand g1392(n2083 ,n2079 ,n2082);
    nand g1393(n1463 ,n1217 ,n980);
    dff g1394(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n512), .Q(n11[0]));
    not g1395(n1259 ,n1138);
    not g1396(n1536 ,n1491);
    nor g1397(n634 ,n488 ,n622);
    or g1398(n1642 ,n1611 ,n1612);
    nand g1399(n848 ,n1869 ,n410);
    nand g1400(n1388 ,n583 ,n837);
    nor g1401(n282 ,n263 ,n271);
    nor g1402(n629 ,n1662 ,n614);
    nand g1403(n1832 ,n2131 ,n2130);
    nand g1404(n851 ,n1888 ,n409);
    nand g1405(n1978 ,n1763 ,n1679);
    xnor g1406(n121 ,n2[39] ,n2[103]);
    nor g1407(n32 ,n2[12] ,n2[76]);
    xnor g1408(n109 ,n2[36] ,n2[100]);
    dff g1409(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1657), .Q(n5[0]));
    dff g1410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1416), .Q(n5[58]));
    nand g1411(n892 ,n1864 ,n410);
    dff g1412(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n559), .Q(n9[1]));
    not g1413(n342 ,n341);
    nand g1414(n712 ,n4[10] ,n402);
    nor g1415(n222 ,n28 ,n221);
    not g1416(n300 ,n299);
    nand g1417(n1322 ,n907 ,n1250);
    nand g1418(n911 ,n1927 ,n731);
    or g1419(n2194 ,n4[58] ,n2192);
    dff g1420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n511), .Q(n11[1]));
    nor g1421(n51 ,n2[35] ,n2[99]);
    nand g1422(n1474 ,n1222 ,n997);
    nand g1423(n1311 ,n895 ,n1240);
    not g1424(n1525 ,n1473);
    nand g1425(n1951 ,n1670 ,n1796);
    dff g1426(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1343), .Q(n4[23]));
    nand g1427(n828 ,n3[27] ,n398);
    not g1428(n452 ,n2[32]);
    xnor g1429(n2021 ,n138 ,n182);
    dff g1430(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1428), .Q(n5[45]));
    not g1431(n2218 ,n9[14]);
    nand g1432(n1744 ,n1669 ,n3[20]);
    nand g1433(n719 ,n4[35] ,n620);
    nor g1434(n157 ,n113 ,n156);
    nand g1435(n681 ,n2[124] ,n629);
    xnor g1436(n2041 ,n136 ,n222);
    nand g1437(n816 ,n3[35] ,n621);
    nand g1438(n1093 ,n1843 ,n729);
    nand g1439(n360 ,n1983 ,n359);
    nor g1440(n573 ,n441 ,n1);
    not g1441(n1539 ,n1495);
    not g1442(n397 ,n621);
    nor g1443(n548 ,n471 ,n1);
    dff g1444(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1323), .Q(n4[41]));
    nand g1445(n1315 ,n3[0] ,n1030);
    xnor g1446(n106 ,n2[57] ,n2[121]);
    nand g1447(n1351 ,n951 ,n1277);
    dff g1448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1622), .Q(n3[12]));
    nand g1449(n1038 ,n1917 ,n729);
    not g1450(n404 ,n731);
    nand g1451(n1972 ,n1762 ,n1760);
    or g1452(n1639 ,n1606 ,n1605);
    nand g1453(n677 ,n2[127] ,n629);
    nand g1454(n284 ,n277 ,n278);
    nand g1455(n821 ,n3[32] ,n621);
    nand g1456(n1998 ,n1757 ,n1741);
    dff g1457(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1417), .Q(n5[57]));
    nand g1458(n1185 ,n766 ,n666);
    not g1459(n427 ,n2[88]);
    nand g1460(n1431 ,n1167 ,n967);
    xnor g1461(n1907 ,n347 ,n1975);
    nor g1462(n607 ,n546 ,n591);
    nand g1463(n1357 ,n888 ,n1283);
    nand g1464(n1605 ,n1097 ,n1387);
    nand g1465(n1992 ,n1714 ,n1709);
    nand g1466(n1999 ,n1682 ,n1765);
    not g1467(n462 ,n2[51]);
    nand g1468(n858 ,n1885 ,n409);
    nand g1469(n958 ,n1898 ,n731);
    nand g1470(n1088 ,n1897 ,n729);
    nand g1471(n2111 ,n4[16] ,n2108);
    dff g1472(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n4[5]));
    nor g1473(n569 ,n474 ,n1);
    nand g1474(n1851 ,n2169 ,n2168);
    not g1475(n465 ,n2[40]);
    nor g1476(n732 ,n1 ,n623);
    nor g1477(n2268 ,n2248 ,n2223);
    nand g1478(n1304 ,n946 ,n1232);
    not g1479(n1249 ,n1121);
    not g1480(n471 ,n2[85]);
    xnor g1481(n83 ,n2[26] ,n2[90]);
    dff g1482(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n537), .Q(n10[29]));
    nand g1483(n825 ,n3[29] ,n398);
    xor g1484(n1869 ,n4[63] ,n2203);
    nor g1485(n255 ,n101 ,n254);
    not g1486(n381 ,n380);
    xnor g1487(n1931 ,n1999 ,n388);
    dff g1488(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n574), .Q(n11[3]));
    not g1489(n1265 ,n1149);
    nand g1490(n1988 ,n1781 ,n1776);
    xnor g1491(n1903 ,n344 ,n1971);
    nor g1492(n62 ,n2[14] ,n2[78]);
    or g1493(n2104 ,n4[13] ,n2102);
    nand g1494(n1597 ,n1074 ,n1551);
    nor g1495(n50 ,n2[28] ,n2[92]);
    nand g1496(n1380 ,n668 ,n869);
    nor g1497(n30 ,n2[10] ,n2[74]);
    nor g1498(n61 ,n2[26] ,n2[90]);
    not g1499(n428 ,n2[80]);
    nor g1500(n209 ,n109 ,n208);
    not g1501(n407 ,n729);
    nand g1502(n2113 ,n4[17] ,n2110);
    nand g1503(n1496 ,n5[2] ,n1032);
    xnor g1504(n99 ,n2[49] ,n2[113]);
    nor g1505(n311 ,n274 ,n309);
    nand g1506(n1719 ,n2024 ,n1666);
    nand g1507(n1802 ,n1666 ,n1798);
    nand g1508(n923 ,n1933 ,n731);
    nand g1509(n1794 ,n1669 ,n3[38]);
    or g1510(n2152 ,n4[37] ,n2150);
    or g1511(n2088 ,n4[5] ,n2087);
    nand g1512(n1009 ,n1925 ,n405);
    dff g1513(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1449), .Q(n5[28]));
    nand g1514(n2283 ,n2279 ,n2280);
    dff g1515(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1474), .Q(n5[10]));
    not g1516(n414 ,n2[65]);
    nand g1517(n966 ,n1894 ,n405);
    or g1518(n2182 ,n4[52] ,n2180);
    nand g1519(n287 ,n266 ,n286);
    nand g1520(n868 ,n1881 ,n410);
    nand g1521(n1379 ,n667 ,n867);
    nand g1522(n1623 ,n863 ,n1404);
    not g1523(n1229 ,n1098);
    nor g1524(n729 ,n1 ,n626);
    nand g1525(n971 ,n1867 ,n409);
    not g1526(n336 ,n335);
    nand g1527(n628 ,n485 ,n619);
    xnor g1528(n2014 ,n104 ,n168);
    nand g1529(n1625 ,n858 ,n1402);
    nand g1530(n1779 ,n1669 ,n3[57]);
    dff g1531(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1481), .Q(n5[7]));
    nor g1532(n533 ,n427 ,n1);
    nor g1533(n168 ,n19 ,n167);
    nand g1534(n859 ,n1835 ,n408);
    nand g1535(n1453 ,n1207 ,n965);
    nand g1536(n1514 ,n827 ,n1085);
    nand g1537(n865 ,n2[12] ,n403);
    nor g1538(n1030 ,n613 ,n643);
    nand g1539(n1306 ,n892 ,n1234);
    xnor g1540(n2004 ,n137 ,n148);
    xnor g1541(n2030 ,n89 ,n200);
    nand g1542(n1580 ,n600 ,n1393);
    not g1543(n371 ,n370);
    nand g1544(n275 ,n1938 ,n1934);
    nor g1545(n2264 ,n2250 ,n2241);
    nand g1546(n618 ,n1662 ,n611);
    not g1547(n2217 ,n9[12]);
    nor g1548(n539 ,n468 ,n1);
    not g1549(n401 ,n620);
    nand g1550(n1773 ,n1669 ,n3[62]);
    nand g1551(n1160 ,n5[46] ,n400);
    xnor g1552(n2012 ,n120 ,n164);
    nor g1553(n228 ,n27 ,n227);
    nand g1554(n674 ,n3[6] ,n621);
    dff g1555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n571), .Q(n11[16]));
    nand g1556(n665 ,n3[12] ,n621);
    nand g1557(n1382 ,n671 ,n874);
    dff g1558(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1432), .Q(n5[42]));
    dff g1559(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1391), .Q(n5[63]));
    dff g1560(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1425), .Q(n5[49]));
    nand g1561(n762 ,n4[59] ,n620);
    not g1562(n395 ,n394);
    dff g1563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1625), .Q(n3[15]));
    nand g1564(n1391 ,n1120 ,n923);
    not g1565(n456 ,n2[89]);
    nand g1566(n1721 ,n1669 ,n3[45]);
    xnor g1567(n117 ,n2[38] ,n2[102]);
    nor g1568(n550 ,n479 ,n1);
    nand g1569(n2109 ,n4[15] ,n2106);
    nand g1570(n860 ,n2[14] ,n403);
    nor g1571(n1660 ,n1 ,n1647);
    not g1572(n409 ,n407);
    nand g1573(n293 ,n1944 ,n292);
    not g1574(n439 ,n2[84]);
    nand g1575(n2084 ,n2075 ,n2083);
    nand g1576(n1459 ,n1214 ,n976);
    dff g1577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n532), .Q(n9[28]));
    dff g1578(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1621), .Q(n3[11]));
    nor g1579(n639 ,n498 ,n622);
    nor g1580(n211 ,n112 ,n210);
    nand g1581(n598 ,n5[1] ,n6[1]);
    nand g1582(n866 ,n1882 ,n410);
    nand g1583(n1751 ,n1668 ,n3[48]);
    nand g1584(n1739 ,n1668 ,n3[30]);
    nand g1585(n1073 ,n1903 ,n408);
    not g1586(n379 ,n378);
    xnor g1587(n130 ,n2[19] ,n2[83]);
    dff g1588(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1455), .Q(n5[23]));
    nor g1589(n238 ,n29 ,n237);
    nand g1590(n956 ,n1912 ,n731);
    nand g1591(n691 ,n4[53] ,n402);
    not g1592(n1253 ,n1128);
    dff g1593(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1439), .Q(n5[33]));
    xnor g1594(n120 ,n2[14] ,n2[78]);
    nand g1595(n852 ,n2[17] ,n730);
    nand g1596(n811 ,n3[39] ,n621);
    nand g1597(n1205 ,n595 ,n641);
    nor g1598(n24 ,n2[6] ,n2[70]);
    nor g1599(n506 ,n2[3] ,n6[3]);
    dff g1600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1431), .Q(n5[43]));
    nand g1601(n1209 ,n5[23] ,n400);
    xnor g1602(n1922 ,n1990 ,n370);
    nor g1603(n575 ,n430 ,n1);
    nand g1604(n720 ,n2[97] ,n629);
    nand g1605(n1989 ,n1795 ,n1790);
    nand g1606(n1587 ,n1053 ,n1542);
    dff g1607(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1459), .Q(n5[18]));
    not g1608(n443 ,n2[39]);
    xnor g1609(n2052 ,n86 ,n244);
    nand g1610(n1163 ,n5[45] ,n400);
    nand g1611(n812 ,n4[36] ,n402);
    nor g1612(n505 ,n5[1] ,n6[1]);
    dff g1613(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1392), .Q(n5[62]));
    nand g1614(n1221 ,n5[11] ,n400);
    nand g1615(n1658 ,n1501 ,n1656);
    nand g1616(n754 ,n2[79] ,n406);
    nor g1617(n2261 ,n2222 ,n2235);
    nand g1618(n1131 ,n714 ,n715);
    xnor g1619(n2053 ,n134 ,n246);
    dff g1620(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1436), .Q(n5[38]));
    nand g1621(n1198 ,n5[30] ,n732);
    nor g1622(n1635 ,n1294 ,n1297);
    not g1623(n1540 ,n1497);
    dff g1624(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1561), .Q(n3[5]));
    nand g1625(n2242 ,n11[25] ,n2210);
    nand g1626(n2249 ,n11[7] ,n11[6]);
    dff g1627(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1318), .Q(n4[46]));
    not g1628(n2207 ,n11[26]);
    not g1629(n1270 ,n1157);
    nand g1630(n755 ,n4[58] ,n402);
    nor g1631(n535 ,n455 ,n1);
    nand g1632(n1862 ,n2191 ,n2190);
    nand g1633(n1456 ,n1211 ,n972);
    xor g1634(n1810 ,n2086 ,n4[4]);
    nand g1635(n2260 ,n2245 ,n2228);
    nor g1636(n184 ,n15 ,n183);
    nand g1637(n1563 ,n987 ,n1521);
    nor g1638(n197 ,n81 ,n196);
    dff g1639(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1310), .Q(n4[53]));
    nand g1640(n1823 ,n2113 ,n2112);
    xnor g1641(n1910 ,n1978 ,n350);
    nand g1642(n1585 ,n602 ,n1292);
    nand g1643(n2175 ,n4[48] ,n2172);
    nand g1644(n1987 ,n1797 ,n1758);
    nand g1645(n1199 ,n5[29] ,n732);
    not g1646(n479 ,n2[82]);
    xnor g1647(n118 ,n2[51] ,n2[115]);
    nand g1648(n1849 ,n2165 ,n2164);
    xnor g1649(n98 ,n2[33] ,n2[97]);
    nand g1650(n1434 ,n1174 ,n929);
    nand g1651(n778 ,n3[63] ,n621);
    nand g1652(n1478 ,n741 ,n1006);
    nand g1653(n1445 ,n1197 ,n1196);
    nand g1654(n741 ,n3[55] ,n398);
    nand g1655(n960 ,n1853 ,n410);
    not g1656(n403 ,n413);
    nor g1657(n262 ,n49 ,n261);
    xnor g1658(n1924 ,n1992 ,n374);
    nand g1659(n1723 ,n2053 ,n1666);
    nand g1660(n1415 ,n1130 ,n908);
    nand g1661(n1681 ,n1668 ,n3[8]);
    nand g1662(n1424 ,n1154 ,n919);
    not g1663(n1667 ,n7[2]);
    nand g1664(n1119 ,n707 ,n751);
    dff g1665(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n552), .Q(n11[28]));
    not g1666(n1557 ,n1516);
    not g1667(n292 ,n291);
    not g1668(n361 ,n360);
    or g1669(n2134 ,n4[28] ,n2132);
    nand g1670(n1015 ,n1923 ,n729);
    xor g1671(n1912 ,n1980 ,n352);
    dff g1672(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n524), .Q(n9[6]));
    nand g1673(n1452 ,n1206 ,n962);
    nand g1674(n744 ,n4[54] ,n402);
    nand g1675(n1108 ,n690 ,n744);
    not g1676(n1260 ,n1140);
    nand g1677(n630 ,n485 ,n617);
    xnor g1678(n2017 ,n130 ,n174);
    nor g1679(n565 ,n424 ,n1);
    nand g1680(n1080 ,n1900 ,n729);
    nand g1681(n1154 ,n5[50] ,n400);
    nand g1682(n747 ,n4[21] ,n402);
    nor g1683(n40 ,n2[24] ,n2[88]);
    nand g1684(n1780 ,n2007 ,n1666);
    dff g1685(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1419), .Q(n5[55]));
    nand g1686(n770 ,n4[46] ,n620);
    nand g1687(n788 ,n4[31] ,n620);
    dff g1688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1321), .Q(n4[43]));
    xnor g1689(n2050 ,n124 ,n240);
    not g1690(n2205 ,n11[17]);
    dff g1691(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1347), .Q(n4[19]));
    nand g1692(n750 ,n2[83] ,n406);
    dff g1693(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n564), .Q(n11[11]));
    nand g1694(n1569 ,n1003 ,n1527);
    nand g1695(n1572 ,n1015 ,n1530);
    nand g1696(n1847 ,n2161 ,n2160);
    nand g1697(n652 ,n3[22] ,n621);
    nand g1698(n864 ,n1836 ,n729);
    nand g1699(n698 ,n4[49] ,n402);
    nor g1700(n2266 ,n2238 ,n2236);
    nor g1701(n638 ,n491 ,n412);
    nand g1702(n942 ,n1849 ,n408);
    dff g1703(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1324), .Q(n4[40]));
    nand g1704(n2187 ,n4[54] ,n2184);
    xnor g1705(n108 ,n2[7] ,n2[71]);
    nand g1706(n1986 ,n1751 ,n1746);
    nor g1707(n46 ,n2[18] ,n2[82]);
    nand g1708(n1316 ,n898 ,n1244);
    or g1709(n2271 ,n2262 ,n2257);
    nand g1710(n1034 ,n2[48] ,n730);
    nand g1711(n1593 ,n1066 ,n1547);
    nor g1712(n182 ,n58 ,n181);
    nand g1713(n1501 ,n5[1] ,n1032);
    nand g1714(n1819 ,n2105 ,n2104);
    or g1715(n2156 ,n4[39] ,n2154);
    nand g1716(n1854 ,n2175 ,n2174);
    nand g1717(n847 ,n2[19] ,n730);
    or g1718(n1644 ,n1614 ,n1445);
    nand g1719(n1130 ,n5[59] ,n732);
    nand g1720(n998 ,n1928 ,n410);
    nand g1721(n1204 ,n594 ,n640);
    nand g1722(n2000 ,n1773 ,n1726);
    nor g1723(n253 ,n123 ,n252);
    nand g1724(n824 ,n4[26] ,n620);
    dff g1725(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1602), .Q(n3[27]));
    nand g1726(n1584 ,n1047 ,n1540);
    nand g1727(n2255 ,n2230 ,n2229);
    nand g1728(n2129 ,n4[25] ,n2126);
    nand g1729(n753 ,n2[80] ,n406);
    nor g1730(n71 ,n2[4] ,n2[68]);
    nand g1731(n2139 ,n4[30] ,n2136);
    xnor g1732(n115 ,n2[11] ,n2[75]);
    nand g1733(n1781 ,n1669 ,n3[50]);
    nand g1734(n869 ,n2[10] ,n730);
    nor g1735(n644 ,n632 ,n625);
    nand g1736(n661 ,n3[14] ,n621);
    nand g1737(n795 ,n4[22] ,n620);
    not g1738(n1250 ,n1122);
    dff g1739(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n561), .Q(n11[9]));
    nand g1740(n1206 ,n5[26] ,n732);
    not g1741(n466 ,n2[73]);
    nand g1742(n1500 ,n808 ,n1052);
    nand g1743(n904 ,n1847 ,n409);
    nand g1744(n1366 ,n4[0] ,n1029);
    nor g1745(n189 ,n83 ,n188);
    nand g1746(n2222 ,n9[18] ,n2215);
    nand g1747(n1657 ,n1069 ,n1653);
    nand g1748(n703 ,n2[110] ,n629);
    nor g1749(n553 ,n458 ,n1);
    or g1750(n2132 ,n4[27] ,n2130);
    nor g1751(n1294 ,n485 ,n1028);
    xnor g1752(n101 ,n2[59] ,n2[123]);
    nand g1753(n1468 ,n781 ,n989);
    dff g1754(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n519), .Q(n9[0]));
    not g1755(n624 ,n623);
    or g1756(n2166 ,n4[44] ,n2164);
    nor g1757(n156 ,n43 ,n155);
    not g1758(n2209 ,n9[4]);
    not g1759(n1236 ,n1105);
    not g1760(n355 ,n354);
    dff g1761(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n548), .Q(n9[21]));
    nand g1762(n1036 ,n1873 ,n405);
    nand g1763(n2282 ,n2281 ,n2278);
    not g1764(n478 ,n2[57]);
    nand g1765(n1579 ,n1040 ,n1537);
    dff g1766(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1591), .Q(n3[38]));
    dff g1767(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n538), .Q(n8[2]));
    nand g1768(n288 ,n276 ,n287);
    nand g1769(n726 ,n4[29] ,n402);
    nand g1770(n707 ,n2[108] ,n406);
    nand g1771(n1134 ,n5[57] ,n732);
    dff g1772(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1603), .Q(n3[26]));
    nand g1773(n1370 ,n655 ,n845);
    nor g1774(n268 ,n1939 ,n1935);
    nand g1775(n1861 ,n2189 ,n2188);
    nand g1776(n873 ,n1878 ,n409);
    nand g1777(n739 ,n4[25] ,n402);
    or g1778(n2110 ,n4[16] ,n2108);
    not g1779(n2221 ,n9[17]);
    dff g1780(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1641), .Q(n3[2]));
    dff g1781(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1646), .Q(n4[0]));
    nand g1782(n1480 ,n826 ,n1092);
    nand g1783(n1645 ,n1499 ,n1585);
    or g1784(n2162 ,n4[42] ,n2160);
    dff g1785(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n542), .Q(n9[26]));
    nand g1786(n1732 ,n2027 ,n1665);
    nand g1787(n1613 ,n948 ,n1363);
    nor g1788(n552 ,n464 ,n1);
    nand g1789(n771 ,n4[15] ,n402);
    not g1790(n408 ,n407);
    not g1791(n2072 ,n4[3]);
    xnor g1792(n2028 ,n81 ,n196);
    nor g1793(n146 ,n71 ,n145);
    nand g1794(n797 ,n4[48] ,n620);
    nor g1795(n247 ,n134 ,n246);
    nand g1796(n1021 ,n1921 ,n729);
    nand g1797(n331 ,n1965 ,n330);
    nand g1798(n1814 ,n2095 ,n2094);
    nand g1799(n1618 ,n873 ,n1409);
    nand g1800(n1207 ,n5[25] ,n400);
    nand g1801(n1044 ,n1914 ,n408);
    xnor g1802(n2033 ,n90 ,n206);
    nand g1803(n784 ,n4[32] ,n620);
    nand g1804(n1314 ,n979 ,n1243);
    not g1805(n2211 ,n9[9]);
    nand g1806(n928 ,n2[49] ,n730);
    nand g1807(n708 ,n2[107] ,n406);
    nor g1808(n640 ,n489 ,n412);
    nand g1809(n1067 ,n2[35] ,n403);
    nand g1810(n735 ,n3[24] ,n621);
    nand g1811(n855 ,n1922 ,n731);
    nand g1812(n1691 ,n2017 ,n1666);
    nand g1813(n1954 ,n1764 ,n1680);
    nor g1814(n145 ,n102 ,n144);
    not g1815(n1237 ,n1107);
    nor g1816(n195 ,n76 ,n194);
    nand g1817(n1692 ,n1668 ,n3[19]);
    nand g1818(n931 ,n1819 ,n408);
    nand g1819(n792 ,n4[33] ,n620);
    nand g1820(n1696 ,n2018 ,n1666);
    nand g1821(n1675 ,n2056 ,n1665);
    nand g1822(n1077 ,n1901 ,n408);
    xnor g1823(n87 ,n2[24] ,n2[88]);
    nand g1824(n790 ,n3[52] ,n621);
    nor g1825(n647 ,n490 ,n622);
    nand g1826(n975 ,n1833 ,n410);
    nor g1827(n636 ,n495 ,n622);
    nor g1828(n42 ,n2[17] ,n2[81]);
    not g1829(n1264 ,n1147);
    nor g1830(n66 ,n2[60] ,n2[124]);
    nand g1831(n689 ,n4[52] ,n620);
    nand g1832(n139 ,n74 ,n93);
    nand g1833(n863 ,n1883 ,n729);
    nand g1834(n1326 ,n878 ,n1254);
    nor g1835(n258 ,n66 ,n257);
    xnor g1836(n116 ,n2[12] ,n2[76]);
    nand g1837(n1104 ,n685 ,n684);
    dff g1838(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1578), .Q(n3[47]));
    nand g1839(n957 ,n1899 ,n731);
    nor g1840(n163 ,n119 ,n162);
    nand g1841(n1562 ,n983 ,n1520);
    nand g1842(n1700 ,n2019 ,n1665);
    not g1843(n351 ,n350);
    nand g1844(n926 ,n1915 ,n731);
    dff g1845(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1444), .Q(n5[31]));
    nand g1846(n669 ,n3[9] ,n621);
    nand g1847(n709 ,n2[105] ,n629);
    nand g1848(n1125 ,n5[61] ,n400);
    nor g1849(n511 ,n446 ,n1);
    nand g1850(n840 ,n1893 ,n408);
    nand g1851(n2145 ,n4[33] ,n2142);
    nand g1852(n1724 ,n1668 ,n3[24]);
    nand g1853(n846 ,n1890 ,n410);
    nor g1854(n500 ,n2[0] ,n6[0]);
    nand g1855(n952 ,n1901 ,n405);
    not g1856(n2201 ,n2200);
    nand g1857(n1693 ,n2051 ,n1665);
    or g1858(n16 ,n2[1] ,n2[65]);
    nand g1859(n1726 ,n2060 ,n1666);
    nand g1860(n1706 ,n2057 ,n1665);
    nand g1861(n954 ,n1900 ,n731);
    nand g1862(n980 ,n1885 ,n405);
    nand g1863(n885 ,n1921 ,n731);
    nand g1864(n1983 ,n1721 ,n1717);
    nand g1865(n1085 ,n2[28] ,n403);
    nand g1866(n1487 ,n817 ,n1022);
    xnor g1867(n6[2] ,n10[30] ,n2284);
    nand g1868(n1024 ,n1874 ,n405);
    nor g1869(n1393 ,n503 ,n1031);
    nand g1870(n819 ,n3[33] ,n621);
    nand g1871(n950 ,n1865 ,n410);
    nand g1872(n1835 ,n2137 ,n2136);
    or g1873(n2270 ,n2255 ,n2260);
    nand g1874(n1631 ,n844 ,n1396);
    nand g1875(n1598 ,n1080 ,n1553);
    or g1876(n2128 ,n4[25] ,n2126);
    not g1877(n434 ,n2[83]);
    nand g1878(n584 ,n2[0] ,n6[0]);
    nand g1879(n660 ,n3[15] ,n621);
    not g1880(n449 ,n2[28]);
    xnor g1881(n1921 ,n1989 ,n368);
    xnor g1882(n2023 ,n88 ,n186);
    nand g1883(n1753 ,n1668 ,n3[2]);
    nand g1884(n666 ,n4[7] ,n620);
    nand g1885(n1767 ,n1668 ,n3[5]);
    nor g1886(n2228 ,n9[11] ,n9[10]);
    nand g1887(n321 ,n1960 ,n320);
    nand g1888(n1124 ,n709 ,n706);
    xnor g1889(n79 ,n2[45] ,n2[109]);
    nand g1890(n394 ,n8[1] ,n8[0]);
    nand g1891(n277 ,n1939 ,n1935);
    xnor g1892(n1891 ,n1959 ,n317);
    nand g1893(n1360 ,n945 ,n1286);
    nand g1894(n1028 ,n733 ,n642);
    dff g1895(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1460), .Q(n5[19]));
    nor g1896(n219 ,n127 ,n218);
    or g1897(n2158 ,n4[40] ,n2156);
    nand g1898(n1214 ,n5[18] ,n732);
    nor g1899(n57 ,n2[46] ,n2[110]);
    nand g1900(n1011 ,n1924 ,n408);
    dff g1901(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1639), .Q(n3[3]));
    nand g1902(n2251 ,n11[21] ,n11[20]);
    nand g1903(n1048 ,n1918 ,n405);
    nand g1904(n1061 ,n2[37] ,n403);
    nand g1905(n1462 ,n1216 ,n978);
    nand g1906(n1364 ,n4[2] ,n1029);
    nand g1907(n1561 ,n882 ,n1412);
    nand g1908(n1069 ,n1870 ,n731);
    xnor g1909(n124 ,n2[52] ,n2[116]);
    nand g1910(n1102 ,n682 ,n762);
    xor g1911(n1798 ,n2065 ,n6[0]);
    not g1912(n1263 ,n1145);
    nand g1913(n1620 ,n870 ,n1407);
    nand g1914(n1651 ,n1051 ,n1588);
    nor g1915(n298 ,n264 ,n297);
    dff g1916(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n521), .Q(n11[23]));
    nand g1917(n602 ,n5[0] ,n6[0]);
    nand g1918(n1730 ,n1669 ,n3[46]);
    nand g1919(n1960 ,n1704 ,n1703);
    nand g1920(n1218 ,n5[14] ,n732);
    nand g1921(n1087 ,n2[27] ,n730);
    not g1922(n2215 ,n9[19]);
    not g1923(n1543 ,n1502);
    dff g1924(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1429), .Q(n5[46]));
    nand g1925(n1220 ,n5[12] ,n732);
    not g1926(n1394 ,n1367);
    nand g1927(n1419 ,n1139 ,n1009);
    nand g1928(n1018 ,n1922 ,n408);
    nor g1929(n512 ,n452 ,n1);
    nand g1930(n717 ,n2[100] ,n629);
    not g1931(n611 ,n610);
    nand g1932(n1057 ,n2[39] ,n403);
    nand g1933(n965 ,n1895 ,n405);
    nand g1934(n1596 ,n1073 ,n1550);
    nor g1935(n837 ,n543 ,n413);
    nor g1936(n498 ,n4[1] ,n6[1]);
    xnor g1937(n1909 ,n1977 ,n348);
    nand g1938(n600 ,n5[3] ,n6[3]);
    dff g1939(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n547), .Q(n9[4]));
    not g1940(n609 ,n608);
    nand g1941(n1712 ,n1668 ,n3[4]);
    nor g1942(n544 ,n485 ,n1);
    nand g1943(n1148 ,n5[51] ,n732);
    nand g1944(n1688 ,n2016 ,n1665);
    nor g1945(n166 ,n62 ,n165);
    nand g1946(n1055 ,n1910 ,n729);
    nand g1947(n1805 ,n1665 ,n1801);
    nand g1948(n1152 ,n738 ,n739);
    nand g1949(n346 ,n1972 ,n343);
    nor g1950(n2245 ,n2211 ,n9[8]);
    nor g1951(n173 ,n128 ,n172);
    xnor g1952(n136 ,n2[43] ,n2[107]);
    not g1953(n400 ,n399);
    nand g1954(n1443 ,n1193 ,n925);
    nand g1955(n1345 ,n1014 ,n1271);
    nand g1956(n390 ,n1999 ,n389);
    nand g1957(n2179 ,n4[50] ,n2176);
    nand g1958(n1567 ,n998 ,n1525);
    nor g1959(n2253 ,n2220 ,n9[29]);
    nand g1960(n913 ,n1856 ,n409);
    nand g1961(n972 ,n1891 ,n731);
    nand g1962(n1714 ,n1668 ,n3[54]);
    nand g1963(n746 ,n2[119] ,n629);
    nand g1964(n920 ,n1919 ,n405);
    nand g1965(n716 ,n4[19] ,n402);
    nand g1966(n597 ,n2[3] ,n6[3]);
    nand g1967(n1420 ,n1141 ,n984);
    not g1968(n1396 ,n1369);
    nand g1969(n736 ,n2[102] ,n629);
    nor g1970(n1291 ,n505 ,n1031);
    or g1971(n616 ,n485 ,n611);
    dff g1972(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1421), .Q(n5[53]));
    nand g1973(n1619 ,n872 ,n1408);
    nand g1974(n1432 ,n1169 ,n956);
    dff g1975(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1426), .Q(n5[48]));
    not g1976(n269 ,n268);
    nand g1977(n2151 ,n4[36] ,n2148);
    nand g1978(n1703 ,n2020 ,n1665);
    nor g1979(n366 ,n272 ,n364);
    nand g1980(n1947 ,n1782 ,n1780);
    nand g1981(n882 ,n1875 ,n408);
    dff g1982(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1332), .Q(n4[32]));
    nand g1983(n273 ,n1979 ,n1978);
    nand g1984(n358 ,n1982 ,n357);
    nand g1985(n1602 ,n1088 ,n1556);
    nand g1986(n867 ,n2[11] ,n730);
    nand g1987(n664 ,n3[18] ,n398);
    not g1988(n314 ,n313);
    nor g1989(n177 ,n131 ,n176);
    nor g1990(n648 ,n507 ,n622);
    xor g1991(n1801 ,n2062 ,n6[3]);
    not g1992(n264 ,n1947);
    nand g1993(n265 ,n1975 ,n1974);
    nand g1994(n1035 ,n1918 ,n408);
    nand g1995(n817 ,n3[50] ,n621);
    dff g1996(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1590), .Q(n3[39]));
    dff g1997(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1354), .Q(n4[12]));
    xnor g1998(n1917 ,n1985 ,n362);
    nand g1999(n1153 ,n740 ,n806);
    nand g2000(n1352 ,n932 ,n1278);
    not g2001(n432 ,n2[58]);
    nand g2002(n842 ,n1892 ,n409);
    nand g2003(n991 ,n1931 ,n409);
    nand g2004(n1981 ,n1705 ,n1702);
    nand g2005(n898 ,n1854 ,n409);
    nand g2006(n2165 ,n4[43] ,n2162);
    xnor g2007(n1889 ,n1957 ,n313);
    nor g2008(n541 ,n433 ,n1);
    dff g2009(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1643), .Q(n4[3]));
    nor g2010(n221 ,n132 ,n220);
    nand g2011(n993 ,n1930 ,n409);
    nand g2012(n1507 ,n816 ,n1067);
    nor g2013(n43 ,n2[9] ,n2[73]);
    not g2014(n464 ,n2[60]);
    nand g2015(n2276 ,n2269 ,n2259);
    or g2016(n2114 ,n4[18] ,n2112);
    nand g2017(n1959 ,n1733 ,n1700);
    not g2018(n93 ,n92);
    nand g2019(n992 ,n2[60] ,n730);
    dff g2020(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1638), .Q(n1662));
    dff g2021(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n533), .Q(n9[24]));
    nand g2022(n727 ,n2[106] ,n629);
    nand g2023(n1698 ,n1669 ,n3[42]);
    dff g2024(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1456), .Q(n5[21]));
    dff g2025(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n568), .Q(n11[24]));
    not g2026(n398 ,n397);
    nor g2027(n208 ,n51 ,n207);
    nor g2028(n835 ,n494 ,n413);
    nand g2029(n1606 ,n887 ,n1299);
    nand g2030(n915 ,n1923 ,n405);
    nand g2031(n917 ,n1811 ,n408);
    nand g2032(n1993 ,n1731 ,n1723);
    nand g2033(n1761 ,n2002 ,n1666);
    or g2034(n2118 ,n4[20] ,n2116);
    xnor g2035(n133 ,n2[21] ,n2[85]);
    nor g2036(n175 ,n130 ,n174);
    nand g2037(n1121 ,n708 ,n748);
    not g2038(n1537 ,n1493);
    nand g2039(n2199 ,n4[60] ,n2196);
    nand g2040(n1964 ,n1720 ,n1719);
    dff g2041(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1304), .Q(n4[60]));
    or g2042(n2142 ,n4[32] ,n2140);
    nand g2043(n875 ,n1813 ,n410);
    nand g2044(n1181 ,n764 ,n763);
    nand g2045(n906 ,n1846 ,n729);
    nor g2046(n149 ,n137 ,n148);
    dff g2047(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1306), .Q(n4[58]));
    nand g2048(n1339 ,n3[1] ,n1030);
    nand g2049(n1327 ,n1093 ,n1255);
    nor g2050(n169 ,n104 ,n168);
    or g2051(n2100 ,n4[11] ,n2098);
    nor g2052(n38 ,n2[61] ,n2[125]);
    nand g2053(n946 ,n1866 ,n410);
    nand g2054(n1095 ,n2[24] ,n403);
    or g2055(n2094 ,n4[8] ,n2092);
    dff g2056(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n566), .Q(n11[25]));
    nor g2057(n178 ,n52 ,n177);
    nand g2058(n905 ,n1931 ,n405);
    or g2059(n643 ,n1 ,n632);
    nand g2060(n1617 ,n884 ,n1413);
    not g2061(n1247 ,n1118);
    xnor g2062(n2056 ,n123 ,n252);
    nand g2063(n912 ,n1926 ,n731);
    nor g2064(n56 ,n2[7] ,n2[71]);
    dff g2065(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1300), .Q(n4[63]));
    nand g2066(n1697 ,n2033 ,n1665);
    nand g2067(n1661 ,n1496 ,n1655);
    not g2068(n435 ,n2[72]);
    nor g2069(n560 ,n481 ,n1);
    nand g2070(n877 ,n1877 ,n409);
    nand g2071(n1856 ,n2179 ,n2178);
    not g2072(n481 ,n2[49]);
    nand g2073(n2159 ,n4[40] ,n2156);
    not g2074(n417 ,n2[67]);
    nand g2075(n656 ,n3[19] ,n621);
    xnor g2076(n1933 ,n392 ,n2001);
    nand g2077(n1946 ,n1681 ,n1778);
    nand g2078(n1450 ,n1203 ,n961);
    not g2079(n326 ,n325);
    nand g2080(n589 ,n4[3] ,n6[3]);
    nor g2081(n223 ,n136 ,n222);
    nand g2082(n1857 ,n2181 ,n2180);
    nand g2083(n1058 ,n1909 ,n408);
    nand g2084(n339 ,n1969 ,n338);
    nand g2085(n1516 ,n831 ,n1089);
    nand g2086(n1338 ,n975 ,n1265);
    nand g2087(n1165 ,n5[44] ,n732);
    nand g2088(n1422 ,n1148 ,n885);
    nand g2089(n1089 ,n2[26] ,n403);
    nand g2090(n1442 ,n1194 ,n1192);
    nand g2091(n752 ,n2[81] ,n629);
    nand g2092(n1953 ,n1677 ,n1676);
    dff g2093(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n515), .Q(n11[5]));
    nor g2094(n2225 ,n11[3] ,n11[2]);
    nand g2095(n723 ,n4[42] ,n620);
    not g2096(n2070 ,n4[2]);
    not g2097(n1523 ,n1469);
    nand g2098(n1963 ,n1716 ,n1715);
    nor g2099(n2254 ,n2246 ,n2244);
    nand g2100(n1649 ,n1036 ,n1580);
    nor g2101(n521 ,n467 ,n1);
    nor g2102(n1648 ,n1 ,n1635);
    nand g2103(n1070 ,n2[34] ,n403);
    nor g2104(n1647 ,n1296 ,n1636);
    nor g2105(n549 ,n434 ,n1);
    not g2106(n1233 ,n1102);
    or g2107(n2186 ,n4[54] ,n2184);
    dff g2108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n513), .Q(n10[31]));
    nand g2109(n779 ,n3[62] ,n621);
    nor g2110(n44 ,n2[32] ,n2[96]);
    nand g2111(n2195 ,n4[58] ,n2192);
    nand g2112(n758 ,n4[13] ,n620);
    not g2113(n1408 ,n1381);
    nand g2114(n1470 ,n1220 ,n990);
    nand g2115(n785 ,n4[20] ,n620);
    not g2116(n415 ,n2[66]);
    nand g2117(n806 ,n4[24] ,n620);
    xnor g2118(n2078 ,n6[3] ,n4[3]);
    nor g2119(n246 ,n33 ,n245);
    nand g2120(n948 ,n1809 ,n410);
    nor g2121(n519 ,n416 ,n1);
    nor g2122(n54 ,n2[44] ,n2[108]);
    not g2123(n1285 ,n1185);
    nor g2124(n2068 ,n395 ,n393);
    or g2125(n2096 ,n4[9] ,n2094);
    nor g2126(n562 ,n472 ,n1);
    nand g2127(n872 ,n1879 ,n409);
    xnor g2128(n1905 ,n346 ,n1973);
    xnor g2129(n1926 ,n1994 ,n378);
    nand g2130(n890 ,n1861 ,n408);
    nor g2131(n45 ,n2[52] ,n2[116]);
    nand g2132(n1023 ,n1920 ,n729);
    nand g2133(n1685 ,n1668 ,n3[17]);
    nand g2134(n1318 ,n900 ,n1246);
    nand g2135(n487 ,n485 ,n411);
    nand g2136(n1574 ,n1021 ,n1532);
    dff g2137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1452), .Q(n5[26]));
    or g2138(n621 ,n544 ,n612);
    nand g2139(n1337 ,n916 ,n1264);
    xnor g2140(n1897 ,n1965 ,n329);
    nor g2141(n52 ,n2[20] ,n2[84]);
    nor g2142(n2227 ,n9[31] ,n9[30]);
    nand g2143(n1215 ,n5[17] ,n732);
    dff g2144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1461), .Q(n5[17]));
    nand g2145(n1776 ,n2048 ,n1666);
    nor g2146(n64 ,n2[27] ,n2[91]);
    nand g2147(n1127 ,n5[60] ,n732);
    nand g2148(n933 ,n1911 ,n405);
    or g2149(n2176 ,n4[49] ,n2174);
    nand g2150(n967 ,n1913 ,n405);
    nor g2151(n516 ,n438 ,n1);
    nand g2152(n1749 ,n2030 ,n1665);
    nand g2153(n1842 ,n2151 ,n2150);
    nand g2154(n1066 ,n1906 ,n408);
    not g2155(n1522 ,n1468);
    dff g2156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n551), .Q(n9[17]));
    or g2157(n1652 ,n1615 ,n1448);
    xnor g2158(n1930 ,n1998 ,n386);
    nand g2159(n2089 ,n4[5] ,n2087);
    nor g2160(n248 ,n14 ,n247);
    nand g2161(n1331 ,n1012 ,n1259);
    nand g2162(n1747 ,n6[3] ,n1668);
    not g2163(n349 ,n348);
    or g2164(n2120 ,n4[21] ,n2118);
    nand g2165(n1289 ,n1125 ,n905);
    dff g2166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1472), .Q(n5[11]));
    nor g2167(n69 ,n2[31] ,n2[95]);
    nand g2168(n1803 ,n1666 ,n1799);
    nand g2169(n1454 ,n1208 ,n966);
    nand g2170(n2141 ,n4[31] ,n2138);
    not g2171(n1234 ,n1103);
    or g2172(n2226 ,n11[9] ,n11[8]);
    nand g2173(n1105 ,n686 ,n780);
    nand g2174(n777 ,n2[82] ,n406);
    nand g2175(n1103 ,n683 ,n755);
    or g2176(n2172 ,n4[47] ,n2170);
    nand g2177(n1356 ,n938 ,n1282);
    nand g2178(n1756 ,n1669 ,n3[33]);
    nand g2179(n1755 ,n1669 ,n3[56]);
    dff g2180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1433), .Q(n5[41]));
    nand g2181(n733 ,n616 ,n628);
    not g2182(n459 ,n2[92]);
    nand g2183(n834 ,n2[91] ,n406);
    nand g2184(n1812 ,n2091 ,n2090);
    dff g2185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1352), .Q(n4[14]));
    nand g2186(n1941 ,n1759 ,n1805);
    xnor g2187(n90 ,n2[35] ,n2[99]);
    nand g2188(n2001 ,n1752 ,n1701);
    xnor g2189(n91 ,n2[62] ,n2[126]);
    nand g2190(n1212 ,n5[20] ,n400);
    nor g2191(n233 ,n107 ,n232);
    nand g2192(n271 ,n1971 ,n1970);
    nand g2193(n1968 ,n1739 ,n1738);
    nand g2194(n1970 ,n1750 ,n1749);
    nand g2195(n1387 ,n597 ,n838);
    nand g2196(n1323 ,n904 ,n1251);
    xor g2197(n2064 ,n92 ,n74);
    nand g2198(n1428 ,n1163 ,n926);
    nand g2199(n2265 ,n2225 ,n2224);
    nand g2200(n1449 ,n1202 ,n958);
    nand g2201(n1053 ,n1911 ,n408);
    nand g2202(n1416 ,n1132 ,n1078);
    nand g2203(n1564 ,n991 ,n1522);
    not g2204(n357 ,n356);
    nand g2205(n743 ,n4[12] ,n620);
    nand g2206(n1512 ,n823 ,n1079);
    xnor g2207(n1885 ,n1953 ,n307);
    nand g2208(n2163 ,n4[42] ,n2160);
    nand g2209(n1002 ,n2[56] ,n730);
    nand g2210(n353 ,n1978 ,n351);
    nand g2211(n1184 ,n5[36] ,n400);
    nor g2212(n204 ,n20 ,n203);
    nand g2213(n1859 ,n2185 ,n2184);
    dff g2214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n539), .Q(n9[31]));
    nor g2215(n29 ,n2[50] ,n2[114]);
    dff g2216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1309), .Q(n4[54]));
    nand g2217(n1509 ,n819 ,n1072);
    nand g2218(n350 ,n1977 ,n349);
    nand g2219(n368 ,n1988 ,n366);
    not g2220(n1404 ,n1377);
    nand g2221(n1041 ,n2[45] ,n730);
    not g2222(n375 ,n374);
    nand g2223(n1461 ,n1215 ,n977);
    dff g2224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1488), .Q(n5[4]));
    xor g2225(n1874 ,n1942 ,n288);
    nor g2226(n343 ,n271 ,n339);
    nand g2227(n1837 ,n2141 ,n2140);
    nand g2228(n1298 ,n1662 ,n1028);
    dff g2229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1314), .Q(n4[49]));
    xnor g2230(n89 ,n2[32] ,n2[96]);
    or g2231(n622 ,n545 ,n618);
    nand g2232(n1201 ,n585 ,n639);
    nand g2233(n297 ,n1946 ,n296);
    dff g2234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n575), .Q(n11[18]));
    nand g2235(n1768 ,n2055 ,n1666);
    nand g2236(n1504 ,n813 ,n1059);
    xnor g2237(n1923 ,n1991 ,n372);
    dff g2238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1628), .Q(n3[18]));
    nor g2239(n612 ,n1 ,n609);
    nand g2240(n907 ,n1848 ,n410);
    nand g2241(n969 ,n1823 ,n410);
    dff g2242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1633), .Q(n3[23]));
    nand g2243(n2119 ,n4[20] ,n2116);
    not g2244(n474 ,n2[47]);
    not g2245(n365 ,n364);
    dff g2246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1569), .Q(n3[56]));
    nand g2247(n1560 ,n880 ,n1411);
    or g2248(n1031 ,n1 ,n644);
    nand g2249(n1159 ,n745 ,n747);
    nor g2250(n67 ,n2[56] ,n2[120]);
    not g2251(n1395 ,n1368);
    nand g2252(n1848 ,n2163 ,n2162);
    nand g2253(n1081 ,n2[29] ,n730);
    dff g2254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n577), .Q(n11[31]));
    dff g2255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1320), .Q(n4[44]));
    not g2256(n431 ,n2[77]);
    nand g2257(n546 ,n8[0] ,n8[1]);
    nor g2258(n491 ,n2[65] ,n6[1]);
    nand g2259(n1013 ,n2[53] ,n403);
    nand g2260(n1342 ,n921 ,n1268);
    nand g2261(n1817 ,n2101 ,n2100);
    nand g2262(n745 ,n2[85] ,n629);
    nand g2263(n1332 ,n914 ,n1260);
    nand g2264(n884 ,n1874 ,n409);
    nand g2265(n653 ,n3[21] ,n621);
    nand g2266(n73 ,n2[2] ,n2[66]);
    nor g2267(n497 ,n2[66] ,n6[2]);
    xnor g2268(n1899 ,n1967 ,n333);
    nand g2269(n1092 ,n2[54] ,n730);
    dff g2270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n529), .Q(n9[15]));
    dff g2271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1584), .Q(n3[43]));
    nand g2272(n974 ,n1889 ,n405);
    nand g2273(n1138 ,n720 ,n792);
    xnor g2274(n2027 ,n76 ,n194);
    nor g2275(n183 ,n138 ,n182);
    nor g2276(n179 ,n133 ,n178);
    nor g2277(n1293 ,n606 ,n1027);
    nand g2278(n1033 ,n5[4] ,n732);
    nand g2279(n802 ,n3[44] ,n621);
    dff g2280(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1564), .Q(n3[61]));
    nor g2281(n153 ,n126 ,n152);
    nor g2282(n218 ,n21 ,n217);
    nand g2283(n1725 ,n1669 ,n3[27]);
    not g2284(n310 ,n309);
    nand g2285(n1707 ,n2021 ,n1665);
    nand g2286(n1329 ,n910 ,n1257);
    dff g2287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n573), .Q(n11[14]));
    nor g2288(n542 ,n457 ,n1);
    nand g2289(n940 ,n1814 ,n729);
    nand g2290(n1090 ,n1896 ,n729);
    nor g2291(n603 ,n429 ,n1);
    nand g2292(n601 ,n5[2] ,n6[2]);
    nand g2293(n1012 ,n1839 ,n408);
    xnor g2294(n1883 ,n1951 ,n303);
    nand g2295(n1144 ,n5[53] ,n732);
    xnor g2296(n94 ,n2[56] ,n2[120]);
    not g2297(n1654 ,n1649);
    not g2298(n2210 ,n11[24]);
    dff g2299(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1307), .Q(n4[57]));
    nand g2300(n2257 ,n2253 ,n2227);
    nand g2301(n1180 ,n5[38] ,n400);
    nand g2302(n1499 ,n5[0] ,n1032);
    nand g2303(n1065 ,n2[36] ,n730);
    dff g2304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1624), .Q(n3[14]));
    not g2305(n418 ,n2[81]);
    not g2306(n1232 ,n1101);
    nand g2307(n1371 ,n656 ,n847);
    dff g2308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1470), .Q(n5[12]));
    nand g2309(n281 ,n277 ,n269);
    not g2310(n1521 ,n1467);
    xnor g2311(n2019 ,n133 ,n178);
    nand g2312(n382 ,n1995 ,n381);
    dff g2313(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1333), .Q(n4[31]));
    dff g2314(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1316), .Q(n4[48]));
    nand g2315(n1179 ,n713 ,n712);
    dff g2316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1589), .Q(n3[40]));
    nand g2317(n801 ,n2[98] ,n406);
    nand g2318(n1626 ,n854 ,n1401);
    xnor g2319(n1809 ,n2078 ,n2084);
    dff g2320(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1329), .Q(n4[35]));
    or g2321(n2180 ,n4[51] ,n2178);
    nand g2322(n2153 ,n4[37] ,n2150);
    nand g2323(n815 ,n3[36] ,n621);
    not g2324(n2220 ,n9[28]);
    nand g2325(n1123 ,n5[62] ,n400);
    nor g2326(n25 ,n2[49] ,n2[113]);
    nand g2327(n1616 ,n963 ,n1366);
    not g2328(n461 ,n2[43]);
    nor g2329(n547 ,n477 ,n1);
    nand g2330(n291 ,n1943 ,n290);
    nand g2331(n1581 ,n1042 ,n1538);
    not g2332(n2208 ,n9[21]);
    not g2333(n406 ,n412);
    xnor g2334(n6[0] ,n10[28] ,n2284);
    nand g2335(n1850 ,n2167 ,n2166);
    nor g2336(n206 ,n22 ,n205);
    nand g2337(n1072 ,n2[33] ,n403);
    nand g2338(n973 ,n1890 ,n405);
    nor g2339(n164 ,n35 ,n163);
    nand g2340(n592 ,n3[3] ,n6[3]);
    nand g2341(n1384 ,n674 ,n879);
    xnor g2342(n92 ,n2[1] ,n2[65]);
    nand g2343(n725 ,n2[93] ,n406);
    nor g2344(n198 ,n70 ,n197);
    dff g2345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1579), .Q(n3[46]));
    dff g2346(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1437), .Q(n5[37]));
    not g2347(n1554 ,n1513);
    nand g2348(n1762 ,n1669 ,n3[34]);
    nand g2349(n1502 ,n810 ,n1054);
    dff g2350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n581), .Q(n11[19]));
    nand g2351(n680 ,n2[125] ,n629);
    xnor g2352(n2061 ,n75 ,n262);
    nor g2353(n261 ,n91 ,n260);
    xnor g2354(n97 ,n2[2] ,n2[66]);
    nor g2355(n20 ,n2[33] ,n2[97]);
    nand g2356(n1076 ,n2[31] ,n403);
    not g2357(n480 ,n2[56]);
    nand g2358(n932 ,n1820 ,n408);
    not g2359(n263 ,n1973);
    not g2360(n473 ,n2[37]);
    not g2361(n1255 ,n1131);
    nand g2362(n2135 ,n4[28] ,n2132);
    nand g2363(n853 ,n1887 ,n410);
    nand g2364(n751 ,n4[44] ,n402);
    xnor g2365(n112 ,n2[37] ,n2[101]);
    nand g2366(n1003 ,n1926 ,n729);
    nand g2367(n1444 ,n1195 ,n952);
    not g2368(n1272 ,n1161);
    dff g2369(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1568), .Q(n3[57]));
    xnor g2370(n1894 ,n1962 ,n323);
    nand g2371(n1374 ,n659 ,n856);
    not g2372(n1533 ,n1487);
    not g2373(n631 ,n630);
    nand g2374(n1945 ,n1775 ,n1774);
    dff g2375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1570), .Q(n3[55]));
    nand g2376(n2115 ,n4[18] ,n2112);
    dff g2377(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1305), .Q(n4[59]));
    not g2378(n405 ,n404);
    xnor g2379(n1879 ,n1947 ,n297);
    nand g2380(n1056 ,n1829 ,n729);
    nand g2381(n1985 ,n1740 ,n1735);
    nand g2382(n1955 ,n1685 ,n1683);
    nand g2383(n2252 ,n11[23] ,n11[22]);
    nor g2384(n527 ,n453 ,n1);
    or g2385(n2102 ,n4[12] ,n2100);
    nand g2386(n1112 ,n696 ,n687);
    nand g2387(n2137 ,n4[29] ,n2134);
    nand g2388(n692 ,n2[116] ,n629);
    nand g2389(n1129 ,n736 ,n702);
    nand g2390(n1217 ,n5[15] ,n732);
    nand g2391(n1671 ,n2037 ,n1666);
    dff g2392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n514), .Q(n11[21]));
    nand g2393(n1039 ,n2[46] ,n730);
    nand g2394(n1167 ,n5[43] ,n400);
    nand g2395(n856 ,n2[16] ,n403);
    nor g2396(n580 ,n445 ,n1);
    nor g2397(n225 ,n85 ,n224);
    nor g2398(n571 ,n476 ,n1);
    not g2399(n468 ,n2[95]);
    nand g2400(n1447 ,n1199 ,n957);
    nand g2401(n1225 ,n5[7] ,n400);
    xnor g2402(n100 ,n2[3] ,n2[67]);
    nor g2403(n517 ,n425 ,n1);
    nand g2404(n1350 ,n930 ,n1276);
    nand g2405(n1173 ,n757 ,n758);
    nand g2406(n2233 ,n11[5] ,n2216);
    not g2407(n1273 ,n1162);
    nor g2408(n200 ,n69 ,n199);
    not g2409(n1545 ,n1504);
    nor g2410(n2267 ,n2247 ,n2226);
    nand g2411(n775 ,n4[17] ,n620);
    nand g2412(n679 ,n4[61] ,n620);
    or g2413(n2126 ,n4[24] ,n2124);
    nand g2414(n1690 ,n1668 ,n3[41]);
    nand g2415(n2107 ,n4[14] ,n2104);
    buf g2416(n7[2] ,n1663);
    nor g2417(n192 ,n64 ,n191);
    dff g2418(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1415), .Q(n5[59]));
    nor g2419(n499 ,n4[0] ,n6[0]);
    not g2420(n423 ,n2[53]);
    dff g2421(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n553), .Q(n9[14]));
    nand g2422(n2087 ,n2073 ,n2086);
    nand g2423(n1990 ,n1684 ,n1678);
    dff g2424(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1353), .Q(n4[13]));
    nand g2425(n918 ,n1832 ,n408);
    xnor g2426(n2002 ,n102 ,n144);
    or g2427(n2164 ,n4[43] ,n2162);
    xor g2428(n1800 ,n2063 ,n6[2]);
    nand g2429(n879 ,n2[6] ,n403);
    not g2430(n320 ,n319);
    not g2431(n1279 ,n1173);
    nand g2432(n593 ,n2[65] ,n6[1]);
    nor g2433(n231 ,n82 ,n230);
    nand g2434(n1486 ,n791 ,n1020);
    not g2435(n1555 ,n1514);
    nand g2436(n1446 ,n1198 ,n954);
    nand g2437(n1750 ,n1668 ,n3[32]);
    nand g2438(n1687 ,n1668 ,n3[58]);
    nand g2439(n1164 ,n777 ,n776);
    nand g2440(n1674 ,n1668 ,n3[39]);
    not g2441(n1403 ,n1376);
    nand g2442(n586 ,n4[2] ,n6[2]);
    nand g2443(n1158 ,n5[47] ,n732);
    nand g2444(n1611 ,n897 ,n1315);
    xnor g2445(n78 ,n2[28] ,n2[92]);
    nor g2446(n154 ,n26 ,n153);
    dff g2447(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1599), .Q(n3[31]));
    nand g2448(n2272 ,n2256 ,n2268);
    nand g2449(n1746 ,n2046 ,n1665);
    nor g2450(n620 ,n1 ,n615);
    nand g2451(n1683 ,n2015 ,n1666);
    xnor g2452(n1875 ,n1943 ,n289);
    nand g2453(n272 ,n1987 ,n1986);
    nor g2454(n235 ,n99 ,n234);
    nand g2455(n595 ,n4[0] ,n6[0]);
    dff g2456(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1559), .Q(n3[7]));
    dff g2457(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1457), .Q(n5[22]));
    nand g2458(n1699 ,n1668 ,n3[53]);
    nand g2459(n1157 ,n799 ,n795);
    xnor g2460(n114 ,n2[61] ,n2[125]);
    or g2461(n2138 ,n4[30] ,n2136);
    nor g2462(n49 ,n2[62] ,n2[126]);
    nand g2463(n317 ,n1958 ,n316);
    nand g2464(n1302 ,n971 ,n1231);
    nand g2465(n1497 ,n804 ,n1046);
    nor g2466(n237 ,n110 ,n236);
    not g2467(n429 ,n2[87]);
    nand g2468(n1161 ,n749 ,n785);
    nor g2469(n234 ,n18 ,n233);
    nor g2470(n532 ,n459 ,n1);
    xnor g2471(n85 ,n2[44] ,n2[108]);
    nand g2472(n1022 ,n2[50] ,n730);
    nand g2473(n1313 ,n913 ,n1242);
    nand g2474(n1300 ,n848 ,n1229);
    nor g2475(n191 ,n80 ,n190);
    not g2476(n391 ,n390);
    xnor g2477(n122 ,n2[15] ,n2[79]);
    nand g2478(n1825 ,n2117 ,n2116);
    nand g2479(n2275 ,n2263 ,n2267);
    nand g2480(n2099 ,n4[10] ,n2096);
    nor g2481(n214 ,n63 ,n213);
    not g2482(n308 ,n307);
    nand g2483(n2244 ,n9[20] ,n2208);
    nand g2484(n1571 ,n1011 ,n1529);
    nand g2485(n1484 ,n790 ,n1017);
    nor g2486(n1636 ,n485 ,n1298);
    nand g2487(n909 ,n1871 ,n729);
    nand g2488(n2085 ,n2078 ,n2084);
    nand g2489(n850 ,n2[18] ,n403);
    nand g2490(n1016 ,n1828 ,n729);
    xnor g2491(n2022 ,n87 ,n184);
    nor g2492(n199 ,n84 ,n198);
    dff g2493(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1574), .Q(n3[51]));
    nor g2494(n47 ,n2[41] ,n2[105]);
    nand g2495(n1467 ,n779 ,n986);
    nand g2496(n1764 ,n1669 ,n3[16]);
    nor g2497(n212 ,n31 ,n211);
    nor g2498(n566 ,n478 ,n1);
    nand g2499(n1733 ,n1668 ,n3[21]);
    not g2500(n1535 ,n1490);
    not g2501(n1937 ,n1747);
    nand g2502(n1320 ,n902 ,n1248);
    nand g2503(n914 ,n1838 ,n729);
    xnor g2504(n126 ,n2[8] ,n2[72]);
    nand g2505(n959 ,n1807 ,n409);
    xnor g2506(n110 ,n2[50] ,n2[114]);
    nand g2507(n861 ,n1884 ,n410);
    nand g2508(n1385 ,n675 ,n881);
    nand g2509(n934 ,n1872 ,n409);
    or g2510(n2160 ,n4[41] ,n2158);
    nand g2511(n1427 ,n1158 ,n922);
    nand g2512(n783 ,n3[59] ,n621);
    nand g2513(n295 ,n1945 ,n294);
    nand g2514(n1822 ,n2111 ,n2110);
    or g2515(n1641 ,n1608 ,n1607);
    nand g2516(n1223 ,n5[9] ,n400);
    nand g2517(n1169 ,n5[42] ,n400);
    nor g2518(n196 ,n13 ,n195);
    nand g2519(n1074 ,n1902 ,n408);
    dff g2520(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n526), .Q(n9[12]));
    nand g2521(n1146 ,n5[52] ,n400);
    dff g2522(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1644), .Q(n4[2]));
    nand g2523(n740 ,n2[88] ,n629);
    nand g2524(n994 ,n1881 ,n405);
    nor g2525(n554 ,n431 ,n1);
    nor g2526(n1290 ,n504 ,n1031);
    nand g2527(n1482 ,n789 ,n1013);
    nand g2528(n1676 ,n2013 ,n1665);
    not g2529(n1406 ,n1379);
    xnor g2530(n604 ,n411 ,n485);
    nand g2531(n1591 ,n1060 ,n1545);
    nand g2532(n1844 ,n2155 ,n2154);
    nand g2533(n1632 ,n842 ,n1395);
    nor g2534(n2269 ,n2252 ,n2251);
    dff g2535(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1362), .Q(n4[4]));
    nand g2536(n1498 ,n805 ,n1049);
    not g2537(n1549 ,n1508);
    nand g2538(n1200 ,n593 ,n638);
    nand g2539(n1684 ,n1668 ,n3[52]);
    nand g2540(n1472 ,n1221 ,n994);
    nand g2541(n1790 ,n2049 ,n1666);
    nand g2542(n930 ,n1822 ,n409);
    nand g2543(n1367 ,n650 ,n839);
endmodule
