module top (n0, n1, n2, n3, n4, n7, n8, n5, n6, n9, n11, n12, n13, n10);
    input n0, n1, n2, n3, n4, n5, n6;
    input [1:0] n7;
    input [7:0] n8;
    output [7:0] n9, n10;
    output n11, n12, n13;
    wire n0, n1, n2, n3, n4, n5, n6;
    wire [1:0] n7;
    wire [7:0] n8;
    wire [7:0] n9, n10;
    wire n11, n12, n13;
    wire n14, n15, n16, n17, n18, n19, n20, n21;
    wire n22, n23, n24, n25, n26, n27, n28, n29;
    wire n30, n31, n32, n33, n34, n35, n36, n37;
    wire n38, n39, n40, n41, n42, n43, n44, n45;
    wire n46, n47, n48, n49, n50, n51, n52, n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146;
    dff g0(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n118), .Q(n9[4]));
    nand g1(n144 ,n44 ,n142);
    buf g2(n10[2], n9[2]);
    nand g3(n73 ,n27 ,n61);
    not g4(n20 ,n1);
    nand g5(n85 ,n9[6] ,n88);
    nand g6(n50 ,n5 ,n6);
    nand g7(n94 ,n9[0] ,n88);
    not g8(n113 ,n112);
    nand g9(n87 ,n9[7] ,n88);
    nand g10(n115 ,n121 ,n114);
    nor g11(n48 ,n126 ,n35);
    nand g12(n25 ,n4 ,n8[6]);
    nand g13(n82 ,n9[3] ,n88);
    nor g14(n140 ,n109 ,n138);
    nor g15(n70 ,n54 ,n69);
    or g16(n142 ,n110 ,n141);
    nor g17(n129 ,n128 ,n115);
    nand g18(n102 ,n106 ,n128);
    nand g19(n47 ,n9[7] ,n45);
    or g20(n130 ,n31 ,n121);
    nand g21(n120 ,n41 ,n99);
    nor g22(n88 ,n4 ,n67);
    nand g23(n81 ,n9[1] ,n88);
    not g24(n17 ,n2);
    nand g25(n72 ,n24 ,n59);
    buf g26(n10[3], n9[3]);
    nand g27(n104 ,n84 ,n90);
    nor g28(n126 ,n30 ,n7[1]);
    buf g29(n10[1], n9[1]);
    nand g30(n26 ,n4 ,n8[0]);
    nor g31(n80 ,n68 ,n78);
    nand g32(n99 ,n106 ,n100);
    nor g33(n49 ,n15 ,n53);
    nor g34(n95 ,n70 ,n77);
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n122), .Q(n9[2]));
    nor g36(n93 ,n55 ,n74);
    nand g37(n79 ,n25 ,n64);
    nand g38(n107 ,n106 ,n105);
    nor g39(n137 ,n111 ,n133);
    not g40(n136 ,n132);
    nand g41(n61 ,n9[6] ,n60);
    not g42(n18 ,n9[7]);
    not g43(n69 ,n63);
    nor g44(n90 ,n71 ,n73);
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n125), .Q(n9[3]));
    nand g46(n29 ,n4 ,n8[3]);
    nand g47(n65 ,n9[1] ,n60);
    nand g48(n117 ,n106 ,n97);
    nor g49(n98 ,n105 ,n97);
    nand g50(n57 ,n9[1] ,n63);
    nand g51(n111 ,n100 ,n103);
    not g52(n16 ,n9[4]);
    nand g53(n96 ,n51 ,n87);
    nor g54(n68 ,n50 ,n69);
    nand g55(n27 ,n4 ,n8[5]);
    nor g56(n55 ,n54 ,n53);
    nor g57(n114 ,n17 ,n104);
    nand g58(n143 ,n98 ,n140);
    nand g59(n77 ,n29 ,n58);
    nand g60(n62 ,n9[3] ,n63);
    or g61(n146 ,n33 ,n145);
    nand g62(n110 ,n109 ,n105);
    nand g63(n109 ,n82 ,n95);
    nand g64(n86 ,n9[4] ,n88);
    nand g65(n43 ,n9[0] ,n45);
    nand g66(n58 ,n9[4] ,n60);
    nand g67(n124 ,n43 ,n112);
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n124), .Q(n9[0]));
    nand g69(n64 ,n9[5] ,n63);
    nand g70(n66 ,n9[0] ,n63);
    nand g71(n118 ,n38 ,n117);
    nand g72(n76 ,n28 ,n62);
    nor g73(n131 ,n126 ,n130);
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n134), .Q(n9[7]));
    nand g75(n46 ,n11 ,n45);
    nor g76(n101 ,n100 ,n103);
    not g77(n19 ,n9[3]);
    nor g78(n33 ,n14 ,n2);
    not g79(n32 ,n3);
    nor g80(n63 ,n37 ,n34);
    nand g81(n42 ,n9[6] ,n45);
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n136), .Q(n9[5]));
    nand g83(n132 ,n1 ,n116);
    buf g84(n10[7], n9[7]);
    nand g85(n34 ,n7[1] ,n30);
    buf g86(n10[0], n9[0]);
    nor g87(n56 ,n18 ,n53);
    not g88(n37 ,n36);
    nand g89(n39 ,n9[2] ,n45);
    nor g90(n121 ,n72 ,n96);
    or g91(n139 ,n131 ,n135);
    nand g92(n133 ,n128 ,n123);
    nand g93(n41 ,n9[1] ,n45);
    nor g94(n91 ,n49 ,n76);
    nor g95(n83 ,n56 ,n79);
    nand g96(n31 ,n1 ,n2);
    nor g97(n67 ,n32 ,n48);
    nand g98(n24 ,n4 ,n8[7]);
    buf g99(n10[4], n9[4]);
    nor g100(n52 ,n19 ,n53);
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n146), .Q(n12));
    nand g102(n134 ,n47 ,n130);
    nand g103(n119 ,n42 ,n102);
    nor g104(n36 ,n32 ,n4);
    nor g105(n71 ,n16 ,n69);
    nand g106(n21 ,n4 ,n8[2]);
    nand g107(n100 ,n81 ,n93);
    nand g108(n122 ,n39 ,n107);
    not g109(n106 ,n31);
    nand g110(n138 ,n101 ,n129);
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n120), .Q(n9[1]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n144), .Q(n13));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n119), .Q(n9[6]));
    not g114(n60 ,n53);
    nand g115(n145 ,n1 ,n143);
    not g116(n54 ,n9[2]);
    not g117(n30 ,n7[0]);
    nand g118(n75 ,n21 ,n57);
    nand g119(n44 ,n13 ,n45);
    nand g120(n22 ,n4 ,n8[1]);
    nand g121(n97 ,n86 ,n91);
    nor g122(n23 ,n9[5] ,n2);
    nor g123(n123 ,n121 ,n117);
    nand g124(n108 ,n106 ,n109);
    nand g125(n28 ,n4 ,n8[4]);
    or g126(n51 ,n50 ,n53);
    nand g127(n125 ,n40 ,n108);
    buf g128(n10[6], n9[6]);
    nand g129(n89 ,n9[2] ,n88);
    nand g130(n40 ,n9[3] ,n45);
    nand g131(n127 ,n126 ,n113);
    nand g132(n38 ,n9[4] ,n45);
    nand g133(n141 ,n104 ,n137);
    nor g134(n45 ,n20 ,n2);
    nand g135(n78 ,n26 ,n65);
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n139), .Q(n11));
    nand g137(n128 ,n85 ,n83);
    nand g138(n53 ,n36 ,n126);
    nand g139(n135 ,n46 ,n127);
    nand g140(n105 ,n89 ,n92);
    not g141(n35 ,n34);
    buf g142(n10[5], n9[5]);
    nand g143(n112 ,n106 ,n103);
    nor g144(n92 ,n52 ,n75);
    not g145(n15 ,n9[5]);
    nand g146(n103 ,n94 ,n80);
    not g147(n14 ,n12);
    nand g148(n59 ,n9[6] ,n63);
    nor g149(n116 ,n23 ,n114);
    nand g150(n84 ,n9[5] ,n88);
    nand g151(n74 ,n22 ,n66);
endmodule
