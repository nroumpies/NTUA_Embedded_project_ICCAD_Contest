module top (n0, n1, n4, n5, n2, n3, n9, n6, n7, n8, n15, n16, n10, n11, n12, n13, n14, n17, n18);
    input n0, n1, n2, n3;
    input [31:0] n4, n5;
    input [3:0] n6;
    input [1:0] n7;
    input [7:0] n8;
    output [31:0] n9, n10, n11, n12, n13, n14;
    output [7:0] n15;
    output [3:0] n16;
    output [15:0] n17, n18;
    wire n0, n1, n2, n3;
    wire [31:0] n4, n5;
    wire [3:0] n6;
    wire [1:0] n7;
    wire [7:0] n8;
    wire [31:0] n9, n10, n11, n12, n13, n14;
    wire [7:0] n15;
    wire [3:0] n16;
    wire [15:0] n17, n18;
    wire [31:0] n19;
    wire [31:0] n20;
    wire [7:0] n21;
    wire [31:0] n22;
    wire [3:0] n23;
    wire [31:0] n24;
    wire [31:0] n25;
    wire [3:0] n26;
    wire [7:0] n27;
    wire [31:0] n28;
    wire [7:0] n29;
    wire [31:0] n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
    wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
    wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
    wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
    wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
    wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
    wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
    wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
    wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
    wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
    wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
    wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
    wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
    wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
    wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
    wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
    wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
    wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
    wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
    wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
    wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
    wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
    wire n1735, n1736, n1737, n1738, n1739, n1740, n1741;
    not g0(n1707 ,n24[20]);
    nand g1(n373 ,n24[27] ,n73);
    nand g2(n354 ,n24[19] ,n69);
    or g3(n1629 ,n1409 ,n1575);
    dff g4(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1701), .Q(n29[1]));
    dff g5(.RN(n1685), .SN(1'b1), .CK(n0), .D(n919), .Q(n15[3]));
    nand g6(n421 ,n25[4] ,n83);
    nand g7(n677 ,n5[11] ,n220);
    nand g8(n1063 ,n22[0] ,n946);
    nand g9(n1540 ,n1282 ,n1129);
    nand g10(n621 ,n22[11] ,n84);
    nand g11(n1578 ,n133 ,n1421);
    or g12(n1649 ,n1402 ,n1612);
    nor g13(n147 ,n87 ,n4[2]);
    dff g14(.RN(n1685), .SN(1'b1), .CK(n0), .D(n854), .Q(n10[21]));
    nand g15(n1544 ,n1287 ,n1133);
    dff g16(.RN(n1685), .SN(1'b1), .CK(n0), .D(n727), .Q(n13[14]));
    dff g17(.RN(n1685), .SN(1'b1), .CK(n0), .D(n842), .Q(n14[1]));
    nand g18(n428 ,n25[15] ,n83);
    dff g19(.RN(n1685), .SN(1'b1), .CK(n0), .D(n814), .Q(n24[2]));
    not g20(n92 ,n25[8]);
    nand g21(n649 ,n20[11] ,n80);
    buf g22(n11[31], n10[31]);
    nand g23(n1495 ,n1279 ,n1176);
    nor g24(n265 ,n217 ,n194);
    or g25(n1168 ,n686 ,n1089);
    nand g26(n601 ,n14[0] ,n214);
    nand g27(n672 ,n5[6] ,n220);
    nand g28(n1356 ,n977 ,n1051);
    nand g29(n1066 ,n22[14] ,n946);
    dff g30(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1551), .Q(n28[16]));
    dff g31(.RN(n1685), .SN(1'b1), .CK(n0), .D(n732), .Q(n13[9]));
    nand g32(n497 ,n12[20] ,n214);
    nand g33(n815 ,n312 ,n448);
    nand g34(n43 ,n27[5] ,n42);
    nand g35(n1409 ,n963 ,n1011);
    nor g36(n71 ,n227 ,n228);
    or g37(n1151 ,n668 ,n1019);
    nand g38(n314 ,n24[4] ,n216);
    nand g39(n1328 ,n962 ,n1008);
    nand g40(n1202 ,n30[20] ,n1089);
    nand g41(n922 ,n222 ,n770);
    nand g42(n1196 ,n25[25] ,n1021);
    not g43(n77 ,n76);
    nor g44(n209 ,n169 ,n111);
    dff g45(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1502), .Q(n30[1]));
    or g46(n1117 ,n675 ,n77);
    not g47(n1424 ,n1341);
    nand g48(n691 ,n5[25] ,n220);
    nand g49(n1224 ,n25[4] ,n1021);
    nor g50(n242 ,n217 ,n181);
    buf g51(n11[21], n10[21]);
    nand g52(n399 ,n13[0] ,n214);
    dff g53(.RN(n1685), .SN(1'b1), .CK(n0), .D(n823), .Q(n11[12]));
    nand g54(n1731 ,n1720 ,n1713);
    nand g55(n367 ,n24[20] ,n73);
    nand g56(n341 ,n8[0] ,n80);
    buf g57(n14[25], n10[21]);
    nor g58(n1465 ,n296 ,n1206);
    nand g59(n1364 ,n981 ,n1065);
    or g60(n1131 ,n692 ,n75);
    nand g61(n132 ,n9[17] ,n85);
    nand g62(n1051 ,n28[4] ,n947);
    nand g63(n1273 ,n30[3] ,n79);
    nand g64(n442 ,n25[6] ,n83);
    nand g65(n130 ,n9[7] ,n85);
    nand g66(n1186 ,n30[24] ,n79);
    dff g67(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1661), .Q(n25[17]));
    dff g68(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1624), .Q(n9[22]));
    nand g69(n597 ,n20[8] ,n73);
    nor g70(n303 ,n21[3] ,n172);
    dff g71(.RN(n1685), .SN(1'b1), .CK(n0), .D(n768), .Q(n24[24]));
    nand g72(n581 ,n20[14] ,n80);
    dff g73(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1536), .Q(n28[31]));
    nand g74(n988 ,n25[24] ,n948);
    nand g75(n1298 ,n28[13] ,n75);
    nand g76(n47 ,n27[1] ,n27[0]);
    nand g77(n921 ,n222 ,n809);
    nand g78(n1515 ,n1235 ,n1106);
    nor g79(n268 ,n233 ,n179);
    nand g80(n1222 ,n22[27] ,n1020);
    nand g81(n440 ,n25[7] ,n83);
    or g82(n1140 ,n697 ,n75);
    or g83(n1624 ,n1320 ,n1570);
    nand g84(n513 ,n6[0] ,n83);
    dff g85(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1638), .Q(n9[8]));
    or g86(n1639 ,n1350 ,n1585);
    or g87(n1630 ,n1332 ,n1576);
    buf g88(n17[3], n14[7]);
    nand g89(n150 ,n9[29] ,n85);
    nand g90(n685 ,n5[19] ,n220);
    nand g91(n736 ,n491 ,n291);
    dff g92(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1509), .Q(n22[26]));
    nand g93(n414 ,n10[9] ,n214);
    nand g94(n722 ,n467 ,n301);
    nand g95(n943 ,n3 ,n939);
    nand g96(n863 ,n373 ,n479);
    or g97(n1106 ,n686 ,n1020);
    nand g98(n869 ,n222 ,n606);
    nand g99(n778 ,n356 ,n422);
    nand g100(n1286 ,n28[24] ,n1019);
    nand g101(n874 ,n625 ,n326);
    nand g102(n358 ,n26[1] ,n69);
    not g103(n1437 ,n1367);
    xnor g104(n191 ,n24[10] ,n20[10]);
    dff g105(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1684), .Q(n9[27]));
    nand g106(n547 ,n20[24] ,n73);
    nand g107(n360 ,n24[13] ,n69);
    nand g108(n802 ,n258 ,n290);
    nand g109(n1064 ,n25[0] ,n948);
    nor g110(n1023 ,n136 ,n953);
    nand g111(n163 ,n9[9] ,n85);
    dff g112(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1653), .Q(n25[30]));
    not g113(n1439 ,n1369);
    not g114(n1620 ,n1618);
    not g115(n1447 ,n1386);
    nand g116(n740 ,n416 ,n300);
    nand g117(n938 ,n71 ,n929);
    nand g118(n395 ,n11[0] ,n214);
    dff g119(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1504), .Q(n22[31]));
    nand g120(n1518 ,n1237 ,n1109);
    nand g121(n730 ,n481 ,n286);
    nor g122(n952 ,n88 ,n937);
    nand g123(n1255 ,n22[1] ,n77);
    nand g124(n1335 ,n1066 ,n984);
    nand g125(n349 ,n24[3] ,n73);
    dff g126(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1640), .Q(n9[6]));
    dff g127(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1554), .Q(n28[14]));
    nand g128(n831 ,n569 ,n462);
    nand g129(n1059 ,n28[2] ,n947);
    nand g130(n1563 ,n1308 ,n1149);
    dff g131(.RN(n1685), .SN(1'b1), .CK(n0), .D(n784), .Q(n27[2]));
    or g132(n292 ,n215 ,n195);
    or g133(n1143 ,n677 ,n75);
    not g134(n1416 ,n1327);
    not g135(n91 ,n25[11]);
    nand g136(n1365 ,n5[31] ,n1023);
    nand g137(n520 ,n10[0] ,n82);
    not g138(n1410 ,n1315);
    dff g139(.RN(n1685), .SN(1'b1), .CK(n0), .D(n733), .Q(n13[8]));
    nor g140(n32 ,n29[3] ,n29[2]);
    nor g141(n243 ,n217 ,n173);
    dff g142(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1646), .Q(n9[0]));
    nand g143(n168 ,n9[16] ,n85);
    nand g144(n374 ,n24[22] ,n69);
    nand g145(n711 ,n598 ,n270);
    or g146(n1137 ,n685 ,n1019);
    nor g147(n1713 ,n24[1] ,n24[0]);
    dff g148(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1563), .Q(n28[4]));
    nand g149(n424 ,n10[1] ,n82);
    dff g150(.RN(n1685), .SN(1'b1), .CK(n0), .D(n756), .Q(n24[31]));
    dff g151(.RN(n1685), .SN(1'b1), .CK(n0), .D(n713), .Q(n13[28]));
    nand g152(n1484 ,n1262 ,n1169);
    nand g153(n540 ,n20[8] ,n216);
    nand g154(n1304 ,n28[8] ,n75);
    or g155(n238 ,n215 ,n184);
    nand g156(n1610 ,n148 ,n1453);
    nand g157(n329 ,n24[18] ,n81);
    nor g158(n1462 ,n249 ,n1199);
    nand g159(n207 ,n147 ,n72);
    nand g160(n1407 ,n1082 ,n1083);
    xnor g161(n180 ,n24[31] ,n20[31]);
    nand g162(n518 ,n10[24] ,n215);
    nor g163(n939 ,n252 ,n927);
    nand g164(n776 ,n354 ,n419);
    buf g165(n14[20], n10[16]);
    dff g166(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1650), .Q(n9[28]));
    dff g167(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1673), .Q(n25[21]));
    dff g168(.RN(n1685), .SN(1'b1), .CK(n0), .D(n780), .Q(n24[17]));
    nand g169(n523 ,n27[5] ,n217);
    nand g170(n619 ,n10[7] ,n215);
    not g171(n140 ,n139);
    dff g172(.RN(n1685), .SN(1'b1), .CK(n0), .D(n899), .Q(n14[4]));
    or g173(n1643 ,n1358 ,n1589);
    or g174(n1645 ,n1362 ,n1591);
    nor g175(n109 ,n6[1] ,n6[0]);
    dff g176(.RN(n1685), .SN(1'b1), .CK(n0), .D(n855), .Q(n20[2]));
    dff g177(.RN(n1685), .SN(1'b1), .CK(n0), .D(n710), .Q(n13[31]));
    nand g178(n806 ,n357 ,n431);
    xnor g179(n190 ,n24[12] ,n20[12]);
    nand g180(n966 ,n30[19] ,n949);
    or g181(n1647 ,n1399 ,n1610);
    nor g182(n107 ,n4[23] ,n4[22]);
    not g183(n1420 ,n1333);
    nand g184(n206 ,n105 ,n119);
    nand g185(n1549 ,n1292 ,n1138);
    not g186(n1423 ,n1339);
    buf g187(n12[5], n10[5]);
    nand g188(n1530 ,n1249 ,n1121);
    nand g189(n307 ,n229 ,n178);
    nand g190(n143 ,n9[19] ,n85);
    nand g191(n448 ,n25[1] ,n84);
    nand g192(n1558 ,n1302 ,n1250);
    dff g193(.RN(n1685), .SN(1'b1), .CK(n0), .D(n935), .Q(n23[2]));
    nor g194(n52 ,n45 ,n51);
    nand g195(n971 ,n30[10] ,n949);
    nand g196(n660 ,n20[17] ,n80);
    nand g197(n473 ,n13[15] ,n215);
    nand g198(n1229 ,n22[24] ,n77);
    or g199(n944 ,n708 ,n936);
    nand g200(n1519 ,n1239 ,n1110);
    dff g201(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1485), .Q(n30[16]));
    nand g202(n1590 ,n134 ,n1433);
    nand g203(n514 ,n10[31] ,n215);
    dff g204(.RN(n1685), .SN(1'b1), .CK(n0), .D(n882), .Q(n10[7]));
    nand g205(n386 ,n13[25] ,n214);
    nand g206(n1405 ,n1080 ,n1079);
    buf g207(n18[4], n14[4]);
    dff g208(.RN(n1685), .SN(1'b1), .CK(n0), .D(n857), .Q(n12[31]));
    nand g209(n1231 ,n22[23] ,n77);
    nand g210(n406 ,n25[26] ,n83);
    nand g211(n708 ,n453 ,n235);
    nand g212(n793 ,n365 ,n665);
    nand g213(n743 ,n395 ,n310);
    nand g214(n690 ,n5[24] ,n220);
    nand g215(n927 ,n209 ,n924);
    nand g216(n1478 ,n1259 ,n1154);
    nand g217(n443 ,n14[1] ,n82);
    or g218(n274 ,n214 ,n197);
    nand g219(n872 ,n611 ,n327);
    buf g220(n18[9], 1'b0);
    dff g221(.RN(n1685), .SN(1'b1), .CK(n0), .D(n908), .Q(n27[1]));
    nand g222(n728 ,n476 ,n284);
    or g223(n935 ,n234 ,n931);
    dff g224(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1547), .Q(n28[20]));
    nand g225(n980 ,n30[1] ,n949);
    nor g226(n305 ,n15[0] ,n201);
    buf g227(n12[11], n10[11]);
    nand g228(n368 ,n24[21] ,n73);
    or g229(n1127 ,n681 ,n1019);
    nand g230(n998 ,n22[21] ,n946);
    nand g231(n1308 ,n28[4] ,n1019);
    not g232(n75 ,n74);
    nand g233(n352 ,n24[23] ,n69);
    or g234(n276 ,n215 ,n198);
    nand g235(n503 ,n12[22] ,n215);
    dff g236(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1527), .Q(n22[8]));
    xnor g237(n183 ,n24[13] ,n20[13]);
    nand g238(n213 ,n108 ,n109);
    nand g239(n894 ,n483 ,n645);
    not g240(n1432 ,n1357);
    dff g241(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1657), .Q(n25[26]));
    nand g242(n670 ,n5[4] ,n220);
    nand g243(n560 ,n20[17] ,n69);
    dff g244(.RN(n1685), .SN(1'b1), .CK(n0), .D(n730), .Q(n13[11]));
    nand g245(n1079 ,n25[27] ,n948);
    nor g246(n1459 ,n237 ,n1189);
    dff g247(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1480), .Q(n30[23]));
    nor g248(n53 ,n27[5] ,n52);
    nand g249(n772 ,n435 ,n595);
    dff g250(.RN(n1685), .SN(1'b1), .CK(n0), .D(n815), .Q(n24[1]));
    or g251(n1171 ,n682 ,n79);
    dff g252(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1700), .Q(n29[2]));
    or g253(n1627 ,n1326 ,n1573);
    nor g254(n121 ,n4[21] ,n4[20]);
    dff g255(.RN(n1685), .SN(1'b1), .CK(n0), .D(n800), .Q(n27[3]));
    nand g256(n1474 ,n1257 ,n1155);
    nor g257(n1701 ,n60 ,n58);
    nand g258(n852 ,n615 ,n466);
    nand g259(n1406 ,n986 ,n1081);
    dff g260(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1698), .Q(n29[4]));
    dff g261(.RN(n1685), .SN(1'b1), .CK(n0), .D(n775), .Q(n20[26]));
    or g262(n1100 ,n692 ,n77);
    nor g263(n40 ,n27[2] ,n27[0]);
    buf g264(n14[14], n10[10]);
    nand g265(n729 ,n478 ,n285);
    dff g266(.RN(n1685), .SN(1'b1), .CK(n0), .D(n719), .Q(n13[22]));
    nand g267(n310 ,n24[0] ,n216);
    or g268(n70 ,n226 ,n802);
    xnor g269(n233 ,n19[0] ,n24[0]);
    dff g270(.RN(n1685), .SN(1'b1), .CK(n0), .D(n859), .Q(n12[21]));
    nor g271(n1207 ,n102 ,n1022);
    nand g272(n1473 ,n1313 ,n1161);
    nand g273(n1655 ,n1194 ,n1596);
    dff g274(.RN(n1685), .SN(1'b1), .CK(n0), .D(n744), .Q(n11[10]));
    buf g275(n14[21], n10[17]);
    nand g276(n149 ,n9[20] ,n85);
    buf g277(n11[25], n10[25]);
    nand g278(n1027 ,n25[12] ,n948);
    dff g279(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1508), .Q(n22[27]));
    or g280(n1646 ,n1364 ,n1592);
    nand g281(n735 ,n489 ,n241);
    nand g282(n624 ,n19[1] ,n69);
    nand g283(n1340 ,n969 ,n1029);
    not g284(n1710 ,n24[25]);
    nand g285(n1359 ,n1057 ,n1058);
    nand g286(n1323 ,n1001 ,n1000);
    nand g287(n537 ,n21[1] ,n69);
    nand g288(n688 ,n5[22] ,n220);
    nand g289(n824 ,n570 ,n457);
    nand g290(n1489 ,n1303 ,n1172);
    or g291(n1159 ,n681 ,n79);
    nand g292(n573 ,n13[22] ,n215);
    dff g293(.RN(n1685), .SN(1'b1), .CK(n0), .D(n822), .Q(n21[1]));
    nand g294(n154 ,n9[10] ,n85);
    nand g295(n1487 ,n1263 ,n1157);
    not g296(n38 ,n27[7]);
    nand g297(n1509 ,n1225 ,n1100);
    nand g298(n787 ,n550 ,n429);
    nor g299(n116 ,n4[9] ,n4[8]);
    or g300(n1096 ,n695 ,n77);
    nand g301(n850 ,n607 ,n584);
    nand g302(n1556 ,n1300 ,n1143);
    nand g303(n784 ,n433 ,n551);
    nand g304(n1674 ,n1376 ,n1463);
    nand g305(n1039 ,n25[8] ,n948);
    nand g306(n1194 ,n25[27] ,n1021);
    nand g307(n372 ,n24[17] ,n73);
    nand g308(n1502 ,n1275 ,n1160);
    or g309(n283 ,n214 ,n191);
    nand g310(n1331 ,n1013 ,n1012);
    not g311(n60 ,n59);
    nand g312(n654 ,n20[3] ,n80);
    or g313(n1169 ,n685 ,n79);
    nand g314(n1721 ,n24[23] ,n1704);
    nand g315(n645 ,n21[3] ,n80);
    nand g316(n362 ,n24[12] ,n73);
    nand g317(n546 ,n20[27] ,n81);
    nand g318(n438 ,n25[10] ,n84);
    nand g319(n821 ,n367 ,n417);
    nor g320(n1199 ,n93 ,n1022);
    nand g321(n1022 ,n135 ,n953);
    nand g322(n661 ,n20[20] ,n69);
    buf g323(n11[20], n10[20]);
    nand g324(n551 ,n1693 ,n218);
    nand g325(n392 ,n11[3] ,n215);
    nand g326(n1232 ,n22[22] ,n1020);
    buf g327(n18[5], n14[5]);
    nand g328(n598 ,n13[30] ,n214);
    nand g329(n862 ,n503 ,n337);
    dff g330(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1473), .Q(n30[30]));
    dff g331(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1474), .Q(n30[29]));
    nor g332(n1717 ,n1703 ,n24[18]);
    nand g333(n1541 ,n1283 ,n1131);
    or g334(n1130 ,n694 ,n75);
    not g335(n1428 ,n1349);
    nand g336(n435 ,n10[10] ,n82);
    or g337(n1108 ,n684 ,n1020);
    nand g338(n169 ,n4[3] ,n4[2]);
    nand g339(n836 ,n580 ,n511);
    buf g340(n12[7], n10[7]);
    nand g341(n632 ,n21[0] ,n216);
    nor g342(n1724 ,n1710 ,n24[24]);
    nor g343(n246 ,n217 ,n197);
    dff g344(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1525), .Q(n22[10]));
    nand g345(n694 ,n5[28] ,n220);
    nor g346(n1715 ,n24[29] ,n24[28]);
    dff g347(.RN(n1685), .SN(1'b1), .CK(n0), .D(n818), .Q(n24[0]));
    dff g348(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1488), .Q(n30[15]));
    nand g349(n1398 ,n1071 ,n1070);
    dff g350(.RN(n1685), .SN(1'b1), .CK(n0), .D(n846), .Q(n15[6]));
    nand g351(n1725 ,n24[13] ,n24[12]);
    or g352(n1628 ,n1328 ,n1574);
    nand g353(n712 ,n596 ,n271);
    nand g354(n337 ,n24[22] ,n216);
    nand g355(n477 ,n22[3] ,n84);
    nand g356(n335 ,n24[24] ,n81);
    dff g357(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1484), .Q(n30[19]));
    dff g358(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1626), .Q(n9[20]));
    nor g359(n1736 ,n1734 ,n1731);
    nand g360(n1003 ,n25[19] ,n948);
    nand g361(n1391 ,n5[5] ,n1023);
    nand g362(n769 ,n544 ,n579);
    nand g363(n1488 ,n1265 ,n1156);
    nand g364(n795 ,n541 ,n420);
    buf g365(n17[14], n10[6]);
    or g366(n1735 ,n1730 ,n1732);
    nand g367(n554 ,n1689 ,n218);
    nand g368(n1043 ,n22[7] ,n946);
    nand g369(n1050 ,n28[5] ,n947);
    dff g370(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1697), .Q(n29[5]));
    or g371(n300 ,n82 ,n212);
    dff g372(.RN(n1685), .SN(1'b1), .CK(n0), .D(n808), .Q(n26[0]));
    nand g373(n1025 ,n22[13] ,n946);
    dff g374(.RN(n1685), .SN(1'b1), .CK(n0), .D(n850), .Q(n20[6]));
    nand g375(n158 ,n9[13] ,n85);
    nand g376(n644 ,n20[29] ,n73);
    nand g377(n716 ,n386 ,n274);
    or g378(n1644 ,n1360 ,n1590);
    nand g379(n542 ,n21[0] ,n69);
    nand g380(n1376 ,n5[20] ,n1023);
    nand g381(n1381 ,n5[15] ,n1023);
    or g382(n288 ,n214 ,n192);
    nand g383(n1226 ,n22[25] ,n1020);
    nand g384(n1192 ,n25[28] ,n1021);
    dff g385(.RN(n1685), .SN(1'b1), .CK(n0), .D(n894), .Q(n14[7]));
    nand g386(n1580 ,n142 ,n1423);
    nand g387(n1575 ,n132 ,n1417);
    nand g388(n1346 ,n972 ,n1036);
    nand g389(n847 ,n587 ,n600);
    nand g390(n1045 ,n22[6] ,n946);
    nand g391(n432 ,n25[13] ,n83);
    nand g392(n1570 ,n144 ,n1412);
    nand g393(n866 ,n498 ,n634);
    nand g394(n164 ,n9[4] ,n85);
    not g395(n93 ,n25[22]);
    nand g396(n1714 ,n24[14] ,n1705);
    xnor g397(n1692 ,n27[3] ,n49);
    nand g398(n720 ,n571 ,n278);
    nand g399(n498 ,n18[3] ,n215);
    nand g400(n1246 ,n22[9] ,n77);
    nand g401(n1349 ,n1043 ,n1042);
    dff g402(.RN(n1685), .SN(1'b1), .CK(n0), .D(n886), .Q(n10[5]));
    dff g403(.RN(n1685), .SN(1'b1), .CK(n0), .D(n825), .Q(n21[2]));
    nand g404(n502 ,n12[27] ,n82);
    dff g405(.RN(n1685), .SN(1'b1), .CK(n0), .D(n813), .Q(n24[3]));
    nor g406(n1208 ,n96 ,n1022);
    dff g407(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1493), .Q(n30[10]));
    dff g408(.RN(n1685), .SN(1'b1), .CK(n0), .D(n798), .Q(n24[7]));
    nand g409(n823 ,n534 ,n328);
    nand g410(n512 ,n10[22] ,n82);
    nor g411(n911 ,n267 ,n705);
    not g412(n1426 ,n1344);
    nand g413(n816 ,n459 ,n561);
    nand g414(n1493 ,n1285 ,n1175);
    nand g415(n1005 ,n28[19] ,n947);
    dff g416(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1629), .Q(n9[17]));
    nand g417(n1361 ,n1061 ,n1060);
    nand g418(n887 ,n521 ,n313);
    buf g419(n17[6], 1'b0);
    nand g420(n884 ,n516 ,n651);
    nand g421(n724 ,n471 ,n297);
    nand g422(n1317 ,n992 ,n991);
    or g423(n289 ,n82 ,n193);
    nand g424(n429 ,n22[23] ,n83);
    nor g425(n934 ,n202 ,n70);
    buf g426(n17[12], n10[4]);
    nand g427(n817 ,n559 ,n410);
    nand g428(n536 ,n11[11] ,n214);
    dff g429(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1496), .Q(n30[7]));
    nand g430(n1235 ,n22[20] ,n1020);
    nand g431(n865 ,n527 ,n343);
    buf g432(n14[3], 1'b0);
    nand g433(n1277 ,n28[31] ,n75);
    not g434(n1414 ,n1323);
    nand g435(n160 ,n9[8] ,n85);
    nand g436(n42 ,n40 ,n41);
    nand g437(n877 ,n613 ,n635);
    dff g438(.RN(n1685), .SN(1'b1), .CK(n0), .D(n801), .Q(n27[0]));
    buf g439(n17[1], n14[5]);
    nand g440(n439 ,n22[20] ,n84);
    or g441(n1125 ,n666 ,n1020);
    nor g442(n251 ,n217 ,n199);
    nand g443(n848 ,n594 ,n329);
    nor g444(n249 ,n217 ,n198);
    dff g445(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1475), .Q(n30[28]));
    or g446(n1178 ,n672 ,n1089);
    nand g447(n901 ,n379 ,n535);
    dff g448(.RN(n1685), .SN(1'b1), .CK(n0), .D(n763), .Q(n20[16]));
    nand g449(n1071 ,n22[30] ,n946);
    nand g450(n446 ,n25[2] ,n84);
    nand g451(n1270 ,n30[6] ,n79);
    nand g452(n1058 ,n25[2] ,n948);
    dff g453(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1683), .Q(n25[2]));
    nand g454(n1481 ,n1218 ,n1167);
    or g455(n1622 ,n1316 ,n1568);
    buf g456(n12[15], n10[15]);
    not g457(n1413 ,n1321);
    or g458(n114 ,n15[2] ,n15[3]);
    nor g459(n1609 ,n912 ,n1452);
    nand g460(n1248 ,n22[7] ,n77);
    nand g461(n68 ,n29[6] ,n67);
    nand g462(n553 ,n20[21] ,n69);
    nand g463(n1565 ,n1310 ,n1151);
    dff g464(.RN(n1685), .SN(1'b1), .CK(n0), .D(n833), .Q(n10[15]));
    nand g465(n975 ,n30[6] ,n949);
    nand g466(n749 ,n390 ,n331);
    dff g467(.RN(n1685), .SN(1'b1), .CK(n0), .D(n723), .Q(n13[18]));
    nand g468(n697 ,n5[15] ,n220);
    xnor g469(n212 ,n20[1] ,n24[1]);
    nand g470(n34 ,n32 ,n31);
    dff g471(.RN(n1685), .SN(1'b1), .CK(n0), .D(n817), .Q(n20[18]));
    nand g472(n646 ,n20[30] ,n80);
    nand g473(n427 ,n22[31] ,n83);
    nand g474(n35 ,n29[4] ,n34);
    nand g475(n1501 ,n1274 ,n1182);
    nand g476(n1337 ,n1025 ,n1024);
    nor g477(n1197 ,n89 ,n1022);
    nand g478(n574 ,n22[5] ,n83);
    nand g479(n431 ,n25[5] ,n83);
    nand g480(n1536 ,n1277 ,n1127);
    xnor g481(n192 ,n24[8] ,n20[8]);
    nand g482(n674 ,n5[8] ,n220);
    nand g483(n745 ,n385 ,n319);
    dff g484(.RN(n1685), .SN(1'b1), .CK(n0), .D(n751), .Q(n11[3]));
    nand g485(n489 ,n13[6] ,n214);
    dff g486(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1636), .Q(n9[10]));
    dff g487(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1482), .Q(n30[21]));
    buf g488(n18[6], n14[6]);
    xnor g489(n179 ,n21[0] ,n26[0]);
    nor g490(n1596 ,n240 ,n1439);
    dff g491(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1630), .Q(n9[16]));
    nand g492(n777 ,n547 ,n423);
    nand g493(n1037 ,n25[9] ,n948);
    dff g494(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1550), .Q(n28[17]));
    nand g495(n1035 ,n28[10] ,n947);
    nand g496(n1491 ,n1294 ,n1173);
    nand g497(n689 ,n5[23] ,n220);
    nand g498(n974 ,n30[7] ,n949);
    nand g499(n1533 ,n1254 ,n1124);
    nand g500(n737 ,n492 ,n292);
    nand g501(n1329 ,n1010 ,n1009);
    nand g502(n605 ,n10[18] ,n215);
    nand g503(n1213 ,n22[30] ,n1020);
    dff g504(.RN(n1685), .SN(1'b1), .CK(n0), .D(n860), .Q(n12[29]));
    nand g505(n751 ,n392 ,n325);
    nor g506(n464 ,n225 ,n219);
    nand g507(n1342 ,n970 ,n1032);
    nand g508(n1215 ,n22[29] ,n1020);
    nand g509(n1520 ,n1240 ,n1111);
    nand g510(n595 ,n20[10] ,n80);
    dff g511(.RN(n1685), .SN(1'b1), .CK(n0), .D(n871), .Q(n15[4]));
    nand g512(n695 ,n5[29] ,n220);
    or g513(n287 ,n214 ,n175);
    dff g514(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1664), .Q(n25[10]));
    nor g515(n200 ,n23[0] ,n137);
    not g516(n100 ,n25[20]);
    nand g517(n956 ,n30[25] ,n949);
    nand g518(n1472 ,n1256 ,n1159);
    nand g519(n733 ,n487 ,n288);
    or g520(n1145 ,n674 ,n1019);
    nand g521(n1727 ,n1716 ,n1724);
    dff g522(.RN(n1685), .SN(1'b1), .CK(n0), .D(n774), .Q(n10[6]));
    not g523(n85 ,n3);
    nand g524(n635 ,n8[1] ,n80);
    nand g525(n1550 ,n1293 ,n1098);
    dff g526(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1534), .Q(n22[1]));
    nand g527(n1616 ,n146 ,n1418);
    nor g528(n948 ,n85 ,n941);
    or g529(n1129 ,n693 ,n75);
    dff g530(.RN(n1685), .SN(1'b1), .CK(n0), .D(n881), .Q(n12[24]));
    nand g531(n1053 ,n22[4] ,n946);
    nand g532(n994 ,n22[22] ,n946);
    nand g533(n562 ,n20[25] ,n69);
    nand g534(n1499 ,n1272 ,n1180);
    dff g535(.RN(n1685), .SN(1'b1), .CK(n0), .D(n841), .Q(n20[10]));
    nand g536(n1209 ,n25[13] ,n1021);
    nand g537(n804 ,n627 ,n486);
    not g538(n94 ,n23[0]);
    dff g539(.RN(n1685), .SN(1'b1), .CK(n0), .D(n779), .Q(n10[9]));
    or g540(n1123 ,n669 ,n1020);
    or g541(n1637 ,n1346 ,n1583);
    nand g542(n347 ,n26[0] ,n218);
    xor g543(n172 ,n24[3] ,n20[3]);
    not g544(n96 ,n25[14]);
    nand g545(n768 ,n369 ,n409);
    not g546(n1685 ,n1);
    nor g547(n247 ,n217 ,n184);
    nand g548(n764 ,n350 ,n406);
    dff g549(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1544), .Q(n28[23]));
    nor g550(n264 ,n217 ,n193);
    nand g551(n1400 ,n1018 ,n1072);
    nand g552(n826 ,n617 ,n340);
    buf g553(n17[11], n10[3]);
    nand g554(n1320 ,n959 ,n996);
    xor g555(n171 ,n24[2] ,n20[2]);
    nand g556(n328 ,n24[12] ,n80);
    nand g557(n1251 ,n22[4] ,n77);
    dff g558(.RN(n1685), .SN(1'b1), .CK(n0), .D(n835), .Q(n14[6]));
    nand g559(n332 ,n24[13] ,n216);
    not g560(n79 ,n78);
    or g561(n1155 ,n695 ,n79);
    nand g562(n1195 ,n25[26] ,n1021);
    nand g563(n548 ,n20[31] ,n80);
    not g564(n89 ,n25[24]);
    nand g565(n885 ,n447 ,n316);
    nand g566(n451 ,n10[6] ,n214);
    nand g567(n331 ,n24[5] ,n81);
    dff g568(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1512), .Q(n22[23]));
    nand g569(n1589 ,n165 ,n1432);
    dff g570(.RN(n1685), .SN(1'b1), .CK(n0), .D(n905), .Q(n11[14]));
    nor g571(n1697 ,n65 ,n67);
    nand g572(n142 ,n9[12] ,n85);
    nand g573(n1665 ,n1220 ,n1605);
    nand g574(n466 ,n22[4] ,n84);
    nand g575(n1571 ,n161 ,n1413);
    nand g576(n859 ,n500 ,n333);
    dff g577(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1531), .Q(n22[4]));
    nand g578(n1740 ,n1729 ,n1739);
    nand g579(n617 ,n12[30] ,n214);
    nand g580(n131 ,n9[18] ,n85);
    nand g581(n471 ,n13[17] ,n214);
    nand g582(n1618 ,n917 ,n1228);
    nand g583(n370 ,n24[25] ,n73);
    nand g584(n521 ,n12[26] ,n215);
    dff g585(.RN(n1685), .SN(1'b1), .CK(n0), .D(n820), .Q(n20[17]));
    nand g586(n967 ,n30[14] ,n949);
    nor g587(n1230 ,n101 ,n1022);
    buf g588(n12[13], n10[13]);
    nand g589(n336 ,n24[15] ,n216);
    nand g590(n721 ,n465 ,n279);
    dff g591(.RN(n1685), .SN(1'b1), .CK(n0), .D(n752), .Q(n11[2]));
    nand g592(n1504 ,n1210 ,n1094);
    nand g593(n312 ,n24[1] ,n69);
    nand g594(n148 ,n9[31] ,n85);
    nand g595(n941 ,n71 ,n934);
    nand g596(n919 ,n629 ,n910);
    nand g597(n139 ,n23[2] ,n94);
    nand g598(n986 ,n30[27] ,n949);
    dff g599(.RN(n1685), .SN(1'b1), .CK(n0), .D(n787), .Q(n20[23]));
    nand g600(n1485 ,n1264 ,n1171);
    buf g601(n18[14], n10[2]);
    nand g602(n1353 ,n1049 ,n1048);
    dff g603(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1519), .Q(n22[16]));
    nor g604(n162 ,n86 ,n4[3]);
    dff g605(.RN(n1685), .SN(1'b1), .CK(n0), .D(n840), .Q(n20[11]));
    nand g606(n1397 ,n1068 ,n1067);
    nand g607(n1652 ,n1395 ,n1471);
    dff g608(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1675), .Q(n25[19]));
    nand g609(n1033 ,n22[10] ,n946);
    nor g610(n1603 ,n302 ,n1446);
    nand g611(n313 ,n24[26] ,n81);
    nand g612(n662 ,n1690 ,n218);
    nand g613(n747 ,n401 ,n321);
    nand g614(n1373 ,n5[23] ,n1023);
    nand g615(n161 ,n9[21] ,n85);
    nand g616(n1297 ,n28[14] ,n75);
    or g617(n1179 ,n671 ,n1089);
    nand g618(n727 ,n475 ,n282);
    dff g619(.RN(n1685), .SN(1'b1), .CK(n0), .D(n866), .Q(n18[3]));
    nand g620(n1327 ,n1006 ,n1007);
    buf g621(n17[0], n14[4]);
    or g622(n239 ,n214 ,n182);
    nand g623(n992 ,n22[23] ,n946);
    dff g624(.RN(n1685), .SN(1'b1), .CK(n0), .D(n804), .Q(n19[0]));
    nand g625(n170 ,n9[26] ,n85);
    not g626(n50 ,n49);
    nand g627(n896 ,n507 ,n655);
    not g628(n1452 ,n1396);
    dff g629(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1639), .Q(n9[7]));
    dff g630(.RN(n1685), .SN(1'b1), .CK(n0), .D(n781), .Q(n24[15]));
    nand g631(n1245 ,n22[10] ,n77);
    dff g632(.RN(n1685), .SN(1'b1), .CK(n0), .D(n749), .Q(n11[5]));
    dff g633(.RN(n1685), .SN(1'b1), .CK(n0), .D(n737), .Q(n13[4]));
    nand g634(n1586 ,n159 ,n1429);
    dff g635(.RN(n1685), .SN(1'b1), .CK(n0), .D(n716), .Q(n13[25]));
    nand g636(n800 ,n530 ,n555);
    not g637(n101 ,n25[1]);
    dff g638(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1537), .Q(n28[28]));
    nand g639(n544 ,n20[27] ,n69);
    nand g640(n491 ,n13[5] ,n215);
    nand g641(n1679 ,n1385 ,n1468);
    nand g642(n827 ,n519 ,n565);
    or g643(n1154 ,n691 ,n79);
    nand g644(n353 ,n24[4] ,n69);
    nand g645(n888 ,n387 ,n659);
    nand g646(n220 ,n23[2] ,n136);
    nand g647(n1611 ,n152 ,n1454);
    nand g648(n1557 ,n1301 ,n1144);
    nand g649(n734 ,n488 ,n289);
    dff g650(.RN(n1685), .SN(1'b1), .CK(n0), .D(n903), .Q(n10[16]));
    nor g651(n1201 ,n100 ,n1022);
    nand g652(n612 ,n22[10] ,n83);
    dff g653(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1532), .Q(n22[3]));
    nand g654(n411 ,n25[3] ,n83);
    nand g655(n485 ,n22[22] ,n83);
    nand g656(n510 ,n25[28] ,n84);
    nor g657(n1466 ,n256 ,n1207);
    nand g658(n567 ,n15[0] ,n223);
    nand g659(n717 ,n425 ,n238);
    dff g660(.RN(n1685), .SN(1'b1), .CK(n0), .D(n858), .Q(n11[15]));
    nand g661(n528 ,n11[15] ,n82);
    or g662(n275 ,n214 ,n232);
    nor g663(n1594 ,n243 ,n1437);
    dff g664(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1497), .Q(n30[6]));
    nand g665(n987 ,n30[26] ,n949);
    nand g666(n797 ,n523 ,n662);
    dff g667(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1644), .Q(n9[2]));
    nand g668(n54 ,n27[5] ,n52);
    dff g669(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1699), .Q(n29[3]));
    dff g670(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1559), .Q(n28[8]));
    nand g671(n1301 ,n28[10] ,n75);
    nand g672(n834 ,n496 ,n646);
    nand g673(n628 ,n21[3] ,n73);
    nand g674(n1220 ,n25[7] ,n1021);
    not g675(n1433 ,n1359);
    dff g676(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1656), .Q(n25[28]));
    nand g677(n1566 ,n1311 ,n1152);
    nand g678(n402 ,n25[30] ,n83);
    or g679(n1621 ,n1314 ,n1616);
    nand g680(n1573 ,n143 ,n1415);
    or g681(n39 ,n27[4] ,n27[3]);
    nor g682(n106 ,n4[17] ,n4[16]);
    dff g683(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1628), .Q(n9[18]));
    nand g684(n665 ,n25[9] ,n84);
    nand g685(n640 ,n16[0] ,n216);
    buf g686(n11[28], n10[28]);
    nand g687(n1055 ,n28[14] ,n947);
    dff g688(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1495), .Q(n30[8]));
    nand g689(n1306 ,n28[6] ,n1019);
    or g690(n236 ,n82 ,n211);
    nand g691(n596 ,n13[29] ,n82);
    dff g692(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1564), .Q(n28[3]));
    nand g693(n561 ,n20[12] ,n81);
    nand g694(n1188 ,n30[28] ,n1089);
    nand g695(n541 ,n20[19] ,n73);
    dff g696(.RN(n1685), .SN(1'b1), .CK(n0), .D(n767), .Q(n24[23]));
    buf g697(n14[12], n10[8]);
    dff g698(.RN(n1685), .SN(1'b1), .CK(n0), .D(n740), .Q(n13[1]));
    not g699(n1430 ,n1353);
    nand g700(n456 ,n10[14] ,n214);
    nand g701(n981 ,n30[0] ,n949);
    nand g702(n506 ,n10[16] ,n215);
    nand g703(n1564 ,n1309 ,n1150);
    dff g704(.RN(n1685), .SN(1'b1), .CK(n0), .D(n849), .Q(n20[7]));
    buf g705(n11[24], n10[24]);
    xnor g706(n1698 ,n29[4] ,n63);
    buf g707(n17[13], n10[5]);
    dff g708(.RN(n1685), .SN(1'b1), .CK(n0), .D(n757), .Q(n20[30]));
    dff g709(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1513), .Q(n22[22]));
    nand g710(n989 ,n22[24] ,n946);
    nand g711(n957 ,n30[24] ,n949);
    dff g712(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1659), .Q(n25[23]));
    not g713(n219 ,n220);
    nand g714(n1009 ,n25[17] ,n948);
    dff g715(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1654), .Q(n25[29]));
    nand g716(n1513 ,n1232 ,n1104);
    dff g717(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1521), .Q(n22[14]));
    dff g718(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1555), .Q(n28[12]));
    or g719(n1097 ,n694 ,n1020);
    nand g720(n496 ,n10[30] ,n215);
    nor g721(n1690 ,n53 ,n55);
    nor g722(n37 ,n29[7] ,n36);
    nand g723(n586 ,n13[26] ,n215);
    dff g724(.RN(n1685), .SN(1'b1), .CK(n0), .D(n907), .Q(n11[11]));
    dff g725(.RN(n1685), .SN(1'b1), .CK(n0), .D(n722), .Q(n13[19]));
    nand g726(n669 ,n5[3] ,n220);
    dff g727(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1506), .Q(n22[29]));
    nand g728(n634 ,n8[3] ,n81);
    dff g729(.RN(n1685), .SN(1'b1), .CK(n0), .D(n877), .Q(n18[1]));
    not g730(n84 ,n69);
    nand g731(n571 ,n13[21] ,n215);
    or g732(n272 ,n214 ,n187);
    nand g733(n557 ,n8[2] ,n225);
    nand g734(n141 ,n9[0] ,n85);
    or g735(n273 ,n82 ,n196);
    or g736(n1166 ,n689 ,n1089);
    dff g737(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1677), .Q(n25[15]));
    nand g738(n1382 ,n5[14] ,n1023);
    dff g739(.RN(n1685), .SN(1'b1), .CK(n0), .D(n738), .Q(n13[3]));
    nand g740(n879 ,n222 ,n567);
    not g741(n1451 ,n1392);
    nand g742(n1234 ,n25[0] ,n1021);
    nand g743(n671 ,n5[5] ,n220);
    or g744(n1111 ,n697 ,n77);
    nand g745(n151 ,n9[11] ,n85);
    nand g746(n470 ,n18[2] ,n82);
    nand g747(n851 ,n608 ,n574);
    nor g748(n253 ,n217 ,n230);
    nand g749(n796 ,n525 ,n554);
    nand g750(n1503 ,n1276 ,n1183);
    nand g751(n704 ,n361 ,n442);
    nor g752(n1605 ,n264 ,n1448);
    nand g753(n1584 ,n160 ,n1427);
    nand g754(n1088 ,n22[3] ,n946);
    dff g755(.RN(n1685), .SN(1'b1), .CK(n0), .D(n704), .Q(n24[6]));
    nand g756(n610 ,n15[6] ,n223);
    nand g757(n639 ,n20[15] ,n80);
    nand g758(n663 ,n20[6] ,n80);
    dff g759(.RN(n1685), .SN(1'b1), .CK(n0), .D(n793), .Q(n24[9]));
    nand g760(n472 ,n13[16] ,n214);
    dff g761(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1672), .Q(n25[22]));
    not g762(n1429 ,n1351);
    nand g763(n765 ,n370 ,n407);
    xnor g764(n231 ,n24[18] ,n20[18]);
    not g765(n221 ,n222);
    nand g766(n1568 ,n145 ,n1410);
    dff g767(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1627), .Q(n9[19]));
    nand g768(n1332 ,n964 ,n1014);
    or g769(n1625 ,n1322 ,n1571);
    nand g770(n398 ,n25[31] ,n83);
    nand g771(n1087 ,n22[25] ,n946);
    nand g772(n227 ,n117 ,n116);
    nand g773(n1319 ,n994 ,n995);
    or g774(n301 ,n214 ,n230);
    nand g775(n1315 ,n989 ,n988);
    nand g776(n1054 ,n25[3] ,n948);
    nand g777(n1543 ,n1286 ,n1132);
    dff g778(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1520), .Q(n22[15]));
    dff g779(.RN(n1685), .SN(1'b1), .CK(n0), .D(n824), .Q(n20[14]));
    or g780(n1161 ,n696 ,n79);
    not g781(n1418 ,n1330);
    nand g782(n965 ,n30[15] ,n949);
    dff g783(.RN(n1685), .SN(1'b1), .CK(n0), .D(n852), .Q(n20[4]));
    not g784(n80 ,n82);
    or g785(n1109 ,n683 ,n1020);
    or g786(n1157 ,n683 ,n79);
    nand g787(n1613 ,n156 ,n1456);
    nand g788(n1016 ,n22[15] ,n946);
    nand g789(n1534 ,n1255 ,n1126);
    dff g790(.RN(n1685), .SN(1'b1), .CK(n0), .D(n717), .Q(n13[24]));
    dff g791(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1558), .Q(n28[9]));
    dff g792(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1548), .Q(n28[19]));
    or g793(n1121 ,n671 ,n77);
    xnor g794(n199 ,n24[20] ,n20[20]);
    nor g795(n1460 ,n247 ,n1197);
    nand g796(n1408 ,n987 ,n1084);
    xnor g797(n195 ,n24[4] ,n20[4]);
    nand g798(n973 ,n30[8] ,n949);
    nand g799(n1592 ,n141 ,n1435);
    nand g800(n773 ,n368 ,n515);
    nand g801(n407 ,n25[25] ,n83);
    or g802(n1094 ,n681 ,n1020);
    dff g803(.RN(n1685), .SN(1'b1), .CK(n0), .D(n789), .Q(n10[28]));
    dff g804(.RN(n1685), .SN(1'b1), .CK(n0), .D(n887), .Q(n12[26]));
    nand g805(n673 ,n5[7] ,n220);
    nand g806(n294 ,n216 ,n171);
    nand g807(n61 ,n29[2] ,n60);
    nand g808(n955 ,n933 ,n945);
    nand g809(n898 ,n526 ,n664);
    dff g810(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1543), .Q(n28[24]));
    nand g811(n1732 ,n1712 ,n1715);
    or g812(n928 ,n701 ,n922);
    dff g813(.RN(n1685), .SN(1'b1), .CK(n0), .D(n783), .Q(n20[25]));
    buf g814(n18[13], n10[1]);
    nand g815(n1559 ,n1304 ,n1145);
    nand g816(n1483 ,n1202 ,n1168);
    nor g817(n1723 ,n1706 ,n24[17]);
    dff g818(.RN(n1685), .SN(1'b1), .CK(n0), .D(n728), .Q(n13[13]));
    nand g819(n338 ,n24[20] ,n80);
    nand g820(n144 ,n9[22] ,n85);
    dff g821(.RN(n1685), .SN(1'b1), .CK(n0), .D(n712), .Q(n13[29]));
    nand g822(n725 ,n472 ,n299);
    buf g823(n18[8], 1'b0);
    nor g824(n699 ,n217 ,n303);
    nand g825(n1547 ,n1290 ,n1136);
    nand g826(n1362 ,n980 ,n1062);
    buf g827(n14[30], n10[26]);
    nand g828(n1281 ,n28[28] ,n1019);
    buf g829(n18[15], n10[3]);
    nor g830(n64 ,n57 ,n63);
    nand g831(n678 ,n5[12] ,n220);
    nand g832(n522 ,n10[21] ,n215);
    nand g833(n582 ,n25[11] ,n83);
    buf g834(n14[11], 1'b0);
    nand g835(n1531 ,n1251 ,n1122);
    nand g836(n1193 ,n30[18] ,n1089);
    nand g837(n715 ,n586 ,n273);
    or g838(n241 ,n215 ,n194);
    dff g839(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1647), .Q(n9[31]));
    nand g840(n350 ,n24[26] ,n69);
    dff g841(.RN(n1685), .SN(1'b1), .CK(n0), .D(n709), .Q(n13[0]));
    nand g842(n908 ,n434 ,n556);
    nand g843(n449 ,n25[0] ,n84);
    buf g844(n14[28], n10[24]);
    dff g845(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1529), .Q(n22[6]));
    or g846(n1144 ,n676 ,n1019);
    nor g847(n1604 ,n261 ,n1447);
    nand g848(n552 ,n20[5] ,n80);
    nand g849(n1243 ,n22[12] ,n77);
    nand g850(n593 ,n15[3] ,n223);
    nand g851(n1011 ,n28[17] ,n947);
    nor g852(n33 ,n29[6] ,n29[5]);
    nand g853(n1554 ,n1297 ,n1141);
    or g854(n1174 ,n677 ,n79);
    nand g855(n1588 ,n164 ,n1431);
    nand g856(n940 ,n380 ,n932);
    nand g857(n564 ,n20[16] ,n73);
    nand g858(n1083 ,n25[26] ,n948);
    buf g859(n11[18], n10[18]);
    not g860(n217 ,n218);
    buf g861(n14[16], n10[12]);
    nand g862(n1733 ,n1711 ,n1718);
    not g863(n99 ,n25[16]);
    nand g864(n1497 ,n1270 ,n1178);
    nand g865(n702 ,n129 ,n304);
    or g866(n1124 ,n668 ,n1020);
    nor g867(n216 ,n23[1] ,n139);
    nand g868(n1004 ,n22[19] ,n946);
    nand g869(n1265 ,n30[15] ,n79);
    not g870(n949 ,n943);
    nand g871(n1654 ,n1191 ,n1594);
    nand g872(n434 ,n27[1] ,n217);
    nand g873(n1372 ,n5[24] ,n1023);
    xnor g874(n1693 ,n27[2] ,n47);
    nand g875(n1506 ,n1215 ,n1096);
    nand g876(n838 ,n509 ,n642);
    nand g877(n1338 ,n968 ,n1026);
    nand g878(n782 ,n371 ,n501);
    dff g879(.RN(n1685), .SN(1'b1), .CK(n0), .D(n753), .Q(n11[1]));
    dff g880(.RN(n1685), .SN(1'b1), .CK(n0), .D(n739), .Q(n13[2]));
    nand g881(n611 ,n12[17] ,n215);
    or g882(n1148 ,n671 ,n1019);
    dff g883(.RN(n1685), .SN(1'b1), .CK(n0), .D(n725), .Q(n13[16]));
    dff g884(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1492), .Q(n30[11]));
    dff g885(.RN(n1685), .SN(1'b1), .CK(n0), .D(n766), .Q(n20[28]));
    nand g886(n1366 ,n5[30] ,n1023);
    nand g887(n1384 ,n5[12] ,n1023);
    nand g888(n844 ,n591 ,n604);
    nand g889(n1085 ,n28[25] ,n947);
    nand g890(n413 ,n25[22] ,n83);
    nand g891(n682 ,n5[16] ,n220);
    or g892(n1632 ,n1336 ,n1578);
    nor g893(n1468 ,n260 ,n1212);
    nand g894(n1017 ,n28[15] ,n947);
    not g895(n1453 ,n1397);
    nand g896(n683 ,n5[17] ,n220);
    nand g897(n380 ,n200 ,n213);
    dff g898(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1477), .Q(n30[26]));
    nand g899(n578 ,n13[23] ,n82);
    nand g900(n589 ,n20[18] ,n80);
    nand g901(n657 ,n21[2] ,n80);
    nand g902(n1719 ,n24[21] ,n1707);
    or g903(n1156 ,n697 ,n1089);
    nand g904(n997 ,n25[21] ,n948);
    nand g905(n741 ,n568 ,n255);
    not g906(n62 ,n61);
    nand g907(n319 ,n24[8] ,n81);
    nand g908(n320 ,n24[28] ,n80);
    buf g909(n14[18], n10[14]);
    nand g910(n524 ,n22[16] ,n83);
    or g911(n1138 ,n684 ,n75);
    nand g912(n762 ,n644 ,n400);
    nand g913(n342 ,n24[31] ,n80);
    nand g914(n1517 ,n1238 ,n1108);
    nand g915(n1344 ,n1038 ,n1037);
    dff g916(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1557), .Q(n28[10]));
    nand g917(n1394 ,n5[2] ,n1023);
    buf g918(n14[23], n10[19]);
    nand g919(n1357 ,n1088 ,n1054);
    nand g920(n509 ,n10[13] ,n215);
    not g921(n1441 ,n1371);
    nand g922(n1238 ,n22[18] ,n77);
    nand g923(n1191 ,n25[29] ,n1021);
    dff g924(.RN(n1685), .SN(1'b1), .CK(n0), .D(n807), .Q(n26[1]));
    nand g925(n843 ,n601 ,n315);
    nand g926(n1529 ,n1090 ,n1120);
    or g927(n1183 ,n666 ,n1089);
    nand g928(n419 ,n25[19] ,n83);
    xnor g929(n193 ,n24[7] ,n20[7]);
    or g930(n1150 ,n669 ,n1019);
    nand g931(n202 ,n123 ,n72);
    xnor g932(n181 ,n24[30] ,n20[30]);
    xnor g933(n184 ,n24[24] ,n20[24]);
    nand g934(n870 ,n470 ,n631);
    nand g935(n1015 ,n25[15] ,n948);
    nand g936(n1676 ,n1380 ,n1465);
    nand g937(n616 ,n20[3] ,n73);
    nand g938(n771 ,n374 ,n413);
    dff g939(.RN(n1685), .SN(1'b1), .CK(n0), .D(n821), .Q(n24[20]));
    dff g940(.RN(n1685), .SN(1'b1), .CK(n0), .D(n788), .Q(n24[12]));
    dff g941(.RN(n1685), .SN(1'b1), .CK(n0), .D(n729), .Q(n13[12]));
    dff g942(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1530), .Q(n22[5]));
    nand g943(n890 ,n454 ,n654);
    or g944(n1142 ,n679 ,n1019);
    nand g945(n1479 ,n1186 ,n1165);
    nor g946(n123 ,n4[3] ,n4[2]);
    nand g947(n1738 ,n1736 ,n1737);
    dff g948(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1660), .Q(n25[18]));
    nand g949(n1211 ,n25[12] ,n1021);
    dff g950(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1486), .Q(n30[18]));
    nand g951(n382 ,n22[30] ,n83);
    nand g952(n488 ,n13[7] ,n82);
    nor g953(n1469 ,n262 ,n1216);
    nand g954(n880 ,n508 ,n341);
    dff g955(.RN(n1685), .SN(1'b1), .CK(n0), .D(n889), .Q(n10[0]));
    nand g956(n1581 ,n151 ,n1424);
    nand g957(n494 ,n13[2] ,n214);
    nand g958(n1567 ,n1312 ,n1153);
    or g959(n281 ,n82 ,n188);
    nand g960(n1274 ,n30[2] ,n1089);
    nand g961(n159 ,n9[6] ,n85);
    nand g962(n559 ,n20[18] ,n73);
    nand g963(n1348 ,n973 ,n1041);
    not g964(n1415 ,n1325);
    not g965(n1021 ,n1022);
    dff g966(.RN(n1685), .SN(1'b1), .CK(n0), .D(n896), .Q(n10[20]));
    nand g967(n422 ,n25[18] ,n83);
    nand g968(n343 ,n24[23] ,n81);
    nand g969(n1492 ,n1267 ,n1174);
    nor g970(n258 ,n208 ,n206);
    nand g971(n752 ,n393 ,n330);
    not g972(n1442 ,n1373);
    nand g973(n1225 ,n22[26] ,n1020);
    nand g974(n1300 ,n28[11] ,n75);
    nand g975(n583 ,n16[1] ,n80);
    nand g976(n810 ,n353 ,n421);
    dff g977(.RN(n1685), .SN(1'b1), .CK(n0), .D(n750), .Q(n11[4]));
    buf g978(n14[2], 1'b0);
    nand g979(n1537 ,n1281 ,n1130);
    nand g980(n1662 ,n1209 ,n1602);
    nand g981(n330 ,n24[2] ,n80);
    dff g982(.RN(n1685), .SN(1'b1), .CK(n0), .D(n928), .Q(n16[2]));
    or g983(n252 ,n227 ,n228);
    nand g984(n351 ,n24[2] ,n69);
    or g985(n1651 ,n1408 ,n1615);
    nand g986(n664 ,n1688 ,n218);
    buf g987(n14[27], n10[23]);
    nand g988(n882 ,n619 ,n641);
    nand g989(n710 ,n599 ,n269);
    or g990(n1641 ,n1354 ,n1587);
    nand g991(n459 ,n10[12] ,n82);
    nand g992(n507 ,n10[20] ,n214);
    nand g993(n1269 ,n30[7] ,n79);
    dff g994(.RN(n1685), .SN(1'b1), .CK(n0), .D(n718), .Q(n13[23]));
    nand g995(n1223 ,n25[5] ,n1021);
    nand g996(n538 ,n20[31] ,n69);
    dff g997(.RN(n1685), .SN(1'b1), .CK(n0), .D(n791), .Q(n24[10]));
    nand g998(n1084 ,n28[26] ,n947);
    xnor g999(n1689 ,n27[6] ,n54);
    nor g1000(n1741 ,n1735 ,n1740);
    nand g1001(n889 ,n520 ,n647);
    nor g1002(n58 ,n29[1] ,n29[0]);
    nand g1003(n311 ,n24[0] ,n69);
    nand g1004(n226 ,n127 ,n124);
    nand g1005(n968 ,n30[13] ,n949);
    not g1006(n1708 ,n24[6]);
    xnor g1007(n174 ,n24[5] ,n20[5]);
    or g1008(n201 ,n15[1] ,n114);
    dff g1009(.RN(n1685), .SN(1'b1), .CK(n0), .D(n748), .Q(n21[0]));
    buf g1010(n11[27], n10[27]);
    not g1011(n102 ,n25[15]);
    nand g1012(n1374 ,n5[22] ,n1023);
    nand g1013(n1330 ,n1087 ,n1086);
    not g1014(n87 ,n4[3]);
    or g1015(n277 ,n140 ,n223);
    nand g1016(n755 ,n538 ,n427);
    nand g1017(n1326 ,n966 ,n1005);
    dff g1018(.RN(n1685), .SN(1'b1), .CK(n0), .D(n834), .Q(n10[30]));
    nand g1019(n1490 ,n1266 ,n1185);
    nand g1020(n526 ,n27[7] ,n217);
    nand g1021(n705 ,n218 ,n307);
    not g1022(n1703 ,n24[19]);
    not g1023(n1446 ,n1384);
    nand g1024(n738 ,n493 ,n293);
    nand g1025(n468 ,n14[6] ,n214);
    dff g1026(.RN(n1685), .SN(1'b1), .CK(n0), .D(n103), .Q(n29[0]));
    nand g1027(n390 ,n11[5] ,n82);
    dff g1028(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1648), .Q(n9[30]));
    nand g1029(n829 ,n456 ,n581);
    buf g1030(n12[0], n10[0]);
    nand g1031(n450 ,n12[24] ,n82);
    nand g1032(n1388 ,n5[8] ,n1023);
    nor g1033(n1718 ,n24[9] ,n24[8]);
    dff g1034(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1632), .Q(n9[14]));
    nor g1035(n119 ,n4[25] ,n4[24]);
    nand g1036(n363 ,n24[11] ,n69);
    nand g1037(n66 ,n29[5] ,n64);
    nor g1038(n125 ,n15[6] ,n15[7]);
    nor g1039(n929 ,n210 ,n70);
    nand g1040(n1576 ,n168 ,n1419);
    nand g1041(n1280 ,n28[29] ,n1019);
    nand g1042(n403 ,n25[29] ,n83);
    nand g1043(n166 ,n9[15] ,n85);
    nand g1044(n693 ,n5[27] ,n220);
    nand g1045(n1077 ,n22[28] ,n946);
    xnor g1046(n178 ,n21[1] ,n26[1]);
    nand g1047(n936 ,n933 ,n932);
    nand g1048(n761 ,n405 ,n577);
    nand g1049(n1385 ,n5[11] ,n1023);
    nand g1050(n1010 ,n22[17] ,n946);
    nand g1051(n1290 ,n28[20] ,n75);
    nand g1052(n480 ,n22[2] ,n84);
    buf g1053(n11[23], n10[23]);
    nand g1054(n1073 ,n25[29] ,n948);
    nor g1055(n1595 ,n244 ,n1438);
    nand g1056(n1062 ,n28[1] ,n947);
    or g1057(n1095 ,n696 ,n1020);
    nand g1058(n607 ,n20[6] ,n69);
    dff g1059(.RN(n1685), .SN(1'b1), .CK(n0), .D(n773), .Q(n24[21]));
    dff g1060(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1549), .Q(n28[18]));
    nor g1061(n124 ,n4[13] ,n4[12]);
    not g1062(n103 ,n29[0]);
    or g1063(n1650 ,n1404 ,n1613);
    dff g1064(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1528), .Q(n22[7]));
    or g1065(n926 ,n698 ,n923);
    dff g1066(.RN(n1685), .SN(1'b1), .CK(n0), .D(n743), .Q(n11[0]));
    dff g1067(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1545), .Q(n28[22]));
    dff g1068(.RN(n1685), .SN(1'b1), .CK(n0), .D(n782), .Q(n24[16]));
    nand g1069(n447 ,n12[25] ,n82);
    nand g1070(n585 ,n20[11] ,n73);
    nand g1071(n770 ,n16[2] ,n464);
    not g1072(n88 ,n2);
    not g1073(n1449 ,n1390);
    nand g1074(n858 ,n528 ,n336);
    nor g1075(n1200 ,n97 ,n1022);
    not g1076(n98 ,n25[9]);
    dff g1077(.RN(n1685), .SN(1'b1), .CK(n0), .D(n863), .Q(n24[27]));
    nand g1078(n531 ,n11[14] ,n215);
    nand g1079(n1258 ,n30[27] ,n79);
    or g1080(n203 ,n8[1] ,n110);
    dff g1081(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1526), .Q(n22[9]));
    or g1082(n1734 ,n1722 ,n1726);
    nand g1083(n873 ,n222 ,n593);
    or g1084(n1134 ,n688 ,n75);
    or g1085(n1162 ,n694 ,n79);
    nor g1086(n126 ,n4[29] ,n4[28]);
    buf g1087(n14[29], n10[25]);
    nand g1088(n223 ,n138 ,n137);
    nor g1089(n1461 ,n250 ,n1200);
    nand g1090(n853 ,n616 ,n477);
    nand g1091(n1347 ,n1040 ,n1039);
    nand g1092(n718 ,n578 ,n275);
    nand g1093(n500 ,n12[21] ,n214);
    dff g1094(.RN(n1685), .SN(1'b1), .CK(n0), .D(n898), .Q(n27[7]));
    or g1095(n1631 ,n1334 ,n1577);
    nor g1096(n267 ,n229 ,n178);
    nand g1097(n758 ,n377 ,n402);
    buf g1098(n17[4], 1'b0);
    nand g1099(n1379 ,n5[17] ,n1023);
    nand g1100(n566 ,n20[15] ,n69);
    nand g1101(n1377 ,n5[19] ,n1023);
    nand g1102(n588 ,n20[10] ,n69);
    nand g1103(n1371 ,n5[25] ,n1023);
    nand g1104(n959 ,n30[22] ,n949);
    nor g1105(n65 ,n29[5] ,n64);
    nand g1106(n1498 ,n1271 ,n1179);
    dff g1107(.RN(n1685), .SN(1'b1), .CK(n0), .D(n827), .Q(n10[25]));
    dff g1108(.RN(n1685), .SN(1'b1), .CK(n0), .D(n711), .Q(n13[30]));
    nand g1109(n465 ,n13[20] ,n215);
    nand g1110(n532 ,n14[4] ,n82);
    or g1111(n1182 ,n668 ,n1089);
    dff g1112(.RN(n1685), .SN(1'b1), .CK(n0), .D(n746), .Q(n11[7]));
    nand g1113(n318 ,n26[1] ,n80);
    not g1114(n1425 ,n1343);
    dff g1115(.RN(n1685), .SN(1'b1), .CK(n0), .D(n745), .Q(n11[8]));
    nand g1116(n857 ,n426 ,n342);
    or g1117(n1098 ,n683 ,n75);
    nand g1118(n636 ,n15[5] ,n223);
    nand g1119(n309 ,n24[1] ,n81);
    nand g1120(n388 ,n11[7] ,n214);
    dff g1121(.RN(n1685), .SN(1'b1), .CK(n0), .D(n755), .Q(n20[31]));
    or g1122(n1152 ,n667 ,n1019);
    nand g1123(n1577 ,n166 ,n1420);
    dff g1124(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1635), .Q(n9[11]));
    nand g1125(n1052 ,n25[4] ,n948);
    dff g1126(.RN(n1685), .SN(1'b1), .CK(n0), .D(n914), .Q(n15[0]));
    not g1127(n1457 ,n1405);
    buf g1128(n14[19], n10[15]);
    nand g1129(n555 ,n1692 ,n218);
    nand g1130(n569 ,n20[13] ,n73);
    nand g1131(n572 ,n15[1] ,n223);
    nand g1132(n790 ,n363 ,n582);
    nand g1133(n1040 ,n22[8] ,n946);
    not g1134(n136 ,n135);
    dff g1135(.RN(n1685), .SN(1'b1), .CK(n0), .D(n921), .Q(n16[3]));
    nand g1136(n1355 ,n1053 ,n1052);
    nand g1137(n1666 ,n1221 ,n1606);
    dff g1138(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1637), .Q(n9[9]));
    not g1139(n1417 ,n1329);
    nor g1140(n1711 ,n24[11] ,n24[10]);
    nand g1141(n1333 ,n1016 ,n1015);
    dff g1142(.RN(n1685), .SN(1'b1), .CK(n0), .D(n920), .Q(n15[2]));
    xnor g1143(n188 ,n24[15] ,n20[15]);
    nand g1144(n808 ,n355 ,n445);
    not g1145(n78 ,n1089);
    nand g1146(n1552 ,n1296 ,n1140);
    not g1147(n48 ,n47);
    nand g1148(n1392 ,n5[4] ,n1023);
    nand g1149(n1266 ,n30[13] ,n79);
    not g1150(n954 ,n951);
    nand g1151(n1279 ,n30[8] ,n1089);
    nand g1152(n530 ,n27[3] ,n217);
    nand g1153(n1562 ,n1307 ,n1148);
    or g1154(n1634 ,n1340 ,n1580);
    nand g1155(n1482 ,n1261 ,n1158);
    nand g1156(n452 ,n22[17] ,n84);
    dff g1157(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1665), .Q(n25[7]));
    dff g1158(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1490), .Q(n30[13]));
    dff g1159(.RN(n1685), .SN(1'b1), .CK(n0), .D(n795), .Q(n20[19]));
    xnor g1160(n189 ,n24[14] ,n20[14]);
    nand g1161(n1070 ,n25[30] ,n948);
    nand g1162(n781 ,n359 ,n428);
    nor g1163(n260 ,n217 ,n177);
    dff g1164(.RN(n1685), .SN(1'b1), .CK(n0), .D(n864), .Q(n21[3]));
    xnor g1165(n198 ,n24[22] ,n20[22]);
    nand g1166(n565 ,n20[25] ,n81);
    nand g1167(n1572 ,n149 ,n1414);
    dff g1168(.RN(n1685), .SN(1'b1), .CK(n0), .D(n806), .Q(n24[5]));
    or g1169(n1633 ,n1338 ,n1579);
    nand g1170(n1579 ,n158 ,n1422);
    xnor g1171(n175 ,n24[9] ,n20[9]);
    nand g1172(n1006 ,n22[18] ,n946);
    dff g1173(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1498), .Q(n30[5]));
    nand g1174(n322 ,n24[11] ,n80);
    nand g1175(n881 ,n450 ,n335);
    nand g1176(n978 ,n30[3] ,n949);
    dff g1177(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1623), .Q(n9[23]));
    dff g1178(.RN(n1685), .SN(1'b1), .CK(n0), .D(n832), .Q(n11[9]));
    nand g1179(n457 ,n22[14] ,n84);
    nand g1180(n1551 ,n1295 ,n1139);
    nand g1181(n609 ,n25[23] ,n84);
    nand g1182(n623 ,n22[21] ,n84);
    or g1183(n1728 ,n1725 ,n1714);
    dff g1184(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1566), .Q(n28[1]));
    nand g1185(n1614 ,n157 ,n1457);
    nand g1186(n750 ,n391 ,n314);
    nand g1187(n953 ,n2 ,n942);
    or g1188(n118 ,n8[1] ,n8[0]);
    nand g1189(n1527 ,n1247 ,n1118);
    or g1190(n1115 ,n677 ,n77);
    xnor g1191(n1700 ,n29[2] ,n59);
    nor g1192(n701 ,n118 ,n557);
    nand g1193(n680 ,n5[14] ,n220);
    nand g1194(n535 ,n25[8] ,n84);
    nand g1195(n1067 ,n25[31] ,n948);
    dff g1196(.RN(n1685), .SN(1'b1), .CK(n0), .D(n829), .Q(n10[14]));
    or g1197(n137 ,n23[1] ,n23[2]);
    nand g1198(n789 ,n517 ,n563);
    dff g1199(.RN(n1685), .SN(1'b1), .CK(n0), .D(n720), .Q(n13[21]));
    nor g1200(n700 ,n217 ,n306);
    not g1201(n1444 ,n1379);
    xnor g1202(n229 ,n19[1] ,n24[1]);
    nand g1203(n1007 ,n25[18] ,n948);
    buf g1204(n14[13], n10[9]);
    xnor g1205(n1696 ,n29[6] ,n66);
    nand g1206(n1360 ,n979 ,n1059);
    nand g1207(n916 ,n618 ,n699);
    nand g1208(n1001 ,n22[20] ,n946);
    dff g1209(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1622), .Q(n9[24]));
    nor g1210(n1212 ,n91 ,n1022);
    nor g1211(n122 ,n4[5] ,n4[4]);
    dff g1212(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1681), .Q(n25[8]));
    nand g1213(n731 ,n482 ,n283);
    nand g1214(n854 ,n522 ,n643);
    not g1215(n910 ,n873);
    dff g1216(.RN(n1685), .SN(1'b1), .CK(n0), .D(n918), .Q(n16[0]));
    dff g1217(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1507), .Q(n22[28]));
    nand g1218(n799 ,n441 ,n656);
    dff g1219(.RN(n1685), .SN(1'b1), .CK(n0), .D(n892), .Q(n10[1]));
    nand g1220(n767 ,n352 ,n609);
    nand g1221(n1305 ,n28[7] ,n1019);
    nand g1222(n1252 ,n22[3] ,n1020);
    nor g1223(n250 ,n217 ,n176);
    dff g1224(.RN(n1685), .SN(1'b1), .CK(n0), .D(n778), .Q(n24[18]));
    buf g1225(n18[12], n10[0]);
    dff g1226(.RN(n1685), .SN(1'b1), .CK(n0), .D(n715), .Q(n13[26]));
    nand g1227(n1272 ,n30[4] ,n79);
    nand g1228(n1008 ,n28[18] ,n947);
    nor g1229(n947 ,n85 ,n937);
    dff g1230(.RN(n1685), .SN(1'b1), .CK(n0), .D(n851), .Q(n20[5]));
    nand g1231(n441 ,n27[4] ,n217);
    nand g1232(n608 ,n20[5] ,n69);
    nand g1233(n614 ,n21[2] ,n171);
    or g1234(n1103 ,n689 ,n1020);
    buf g1235(n14[15], n10[11]);
    nand g1236(n515 ,n25[21] ,n83);
    nor g1237(n304 ,n8[0] ,n203);
    nand g1238(n809 ,n16[3] ,n464);
    nand g1239(n1028 ,n22[12] ,n946);
    nand g1240(n603 ,n22[8] ,n84);
    nand g1241(n469 ,n13[18] ,n214);
    nor g1242(n1716 ,n1709 ,n24[26]);
    buf g1243(n17[5], 1'b0);
    or g1244(n1184 ,n675 ,n1089);
    xnor g1245(n232 ,n24[23] ,n20[23]);
    nand g1246(n1523 ,n1243 ,n1114);
    not g1247(n1427 ,n1347);
    nand g1248(n791 ,n364 ,n438);
    nor g1249(n240 ,n217 ,n187);
    nand g1250(n1663 ,n1211 ,n1603);
    dff g1251(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1669), .Q(n25[0]));
    nand g1252(n1242 ,n22[13] ,n77);
    dff g1253(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1522), .Q(n22[13]));
    nand g1254(n985 ,n30[28] ,n949);
    nand g1255(n760 ,n375 ,n510);
    nand g1256(n357 ,n24[5] ,n73);
    nand g1257(n622 ,n20[2] ,n69);
    nand g1258(n156 ,n9[28] ,n85);
    nand g1259(n920 ,n576 ,n909);
    or g1260(n291 ,n214 ,n174);
    nand g1261(n1322 ,n960 ,n999);
    dff g1262(.RN(n1685), .SN(1'b1), .CK(n0), .D(n869), .Q(n15[7]));
    or g1263(n285 ,n215 ,n190);
    nand g1264(n487 ,n13[8] ,n214);
    xnor g1265(n176 ,n24[21] ,n20[21]);
    not g1266(n90 ,n25[19]);
    nand g1267(n652 ,n20[22] ,n216);
    nand g1268(n1494 ,n1268 ,n1184);
    nand g1269(n1615 ,n170 ,n1458);
    buf g1270(n18[11], 1'b0);
    nand g1271(n210 ,n162 ,n72);
    nand g1272(n653 ,n21[2] ,n73);
    or g1273(n1165 ,n690 ,n79);
    dff g1274(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1472), .Q(n30[31]));
    not g1275(n57 ,n29[4]);
    or g1276(n286 ,n215 ,n177);
    or g1277(n299 ,n82 ,n186);
    not g1278(n224 ,n225);
    nand g1279(n323 ,n24[29] ,n216);
    dff g1280(.RN(n1685), .SN(1'b1), .CK(n0), .D(n777), .Q(n20[24]));
    nand g1281(n1024 ,n25[13] ,n948);
    nand g1282(n825 ,n653 ,n529);
    not g1283(n36 ,n35);
    buf g1284(n14[9], 1'b0);
    nand g1285(n723 ,n469 ,n280);
    nand g1286(n543 ,n20[9] ,n80);
    or g1287(n1146 ,n673 ,n1019);
    dff g1288(.RN(n1685), .SN(1'b1), .CK(n0), .D(n902), .Q(n10[31]));
    nand g1289(n1538 ,n1278 ,n1128);
    xnor g1290(n1688 ,n27[7] ,n56);
    dff g1291(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1680), .Q(n25[9]));
    nand g1292(n1233 ,n22[21] ,n77);
    nand g1293(n1086 ,n25[25] ,n948);
    dff g1294(.RN(n1685), .SN(1'b1), .CK(n0), .D(n810), .Q(n24[4]));
    nand g1295(n1312 ,n28[0] ,n1019);
    nand g1296(n1283 ,n28[26] ,n1019);
    nand g1297(n1228 ,n25[2] ,n1021);
    nor g1298(n930 ,n207 ,n70);
    nand g1299(n839 ,n222 ,n638);
    nand g1300(n1352 ,n975 ,n1047);
    nand g1301(n1268 ,n30[9] ,n79);
    nand g1302(n1321 ,n998 ,n997);
    or g1303(n1684 ,n1406 ,n1614);
    or g1304(n113 ,n8[5] ,n8[4]);
    nand g1305(n918 ,n812 ,n803);
    dff g1306(.RN(n1685), .SN(1'b1), .CK(n0), .D(n926), .Q(n16[1]));
    not g1307(n95 ,n25[31]);
    nand g1308(n44 ,n38 ,n43);
    nand g1309(n539 ,n20[30] ,n73);
    buf g1310(n12[12], n10[12]);
    nor g1311(n1608 ,n266 ,n1451);
    nand g1312(n798 ,n378 ,n440);
    dff g1313(.RN(n1685), .SN(1'b1), .CK(n0), .D(n726), .Q(n13[15]));
    nand g1314(n626 ,n10[17] ,n214);
    dff g1315(.RN(n1685), .SN(1'b1), .CK(n0), .D(n758), .Q(n24[30]));
    dff g1316(.RN(n1685), .SN(1'b1), .CK(n0), .D(n853), .Q(n20[3]));
    dff g1317(.RN(n1685), .SN(1'b1), .CK(n0), .D(n904), .Q(n14[5]));
    or g1318(n914 ,n879 ,n878);
    nand g1319(n1339 ,n1028 ,n1027);
    xnor g1320(n182 ,n24[28] ,n20[28]);
    nand g1321(n478 ,n13[12] ,n82);
    dff g1322(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1695), .Q(n29[7]));
    buf g1323(n17[7], 1'b0);
    nand g1324(n982 ,n30[29] ,n949);
    not g1325(n1705 ,n24[15]);
    nand g1326(n1546 ,n1289 ,n1135);
    nand g1327(n1295 ,n28[16] ,n75);
    buf g1328(n12[8], n10[8]);
    nand g1329(n1673 ,n1375 ,n1461);
    nand g1330(n828 ,n397 ,n320);
    nand g1331(n1014 ,n28[16] ,n947);
    dff g1332(.RN(n1685), .SN(1'b1), .CK(n0), .D(n759), .Q(n24[29]));
    nor g1333(n1737 ,n1728 ,n1733);
    nand g1334(n1399 ,n983 ,n1069);
    nand g1335(n204 ,n112 ,n106);
    not g1336(n97 ,n25[21]);
    nand g1337(n1476 ,n1258 ,n1163);
    nand g1338(n904 ,n504 ,n658);
    nand g1339(n348 ,n24[31] ,n69);
    nand g1340(n868 ,n495 ,n339);
    nand g1341(n397 ,n12[28] ,n214);
    or g1342(n1092 ,n691 ,n75);
    dff g1343(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1649), .Q(n9[29]));
    dff g1344(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1541), .Q(n28[26]));
    nand g1345(n604 ,n22[9] ,n84);
    nand g1346(n709 ,n399 ,n236);
    not g1347(n74 ,n1019);
    nand g1348(n1730 ,n1717 ,n1723);
    nand g1349(n996 ,n28[22] ,n947);
    dff g1350(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1633), .Q(n9[13]));
    or g1351(n278 ,n82 ,n176);
    nand g1352(n138 ,n23[0] ,n23[1]);
    or g1353(n1104 ,n688 ,n77);
    nand g1354(n763 ,n564 ,n524);
    dff g1355(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1655), .Q(n25[27]));
    nand g1356(n483 ,n14[7] ,n215);
    dff g1357(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1645), .Q(n9[1]));
    xnor g1358(n187 ,n24[27] ,n20[27]);
    nand g1359(n1038 ,n22[9] ,n946);
    nand g1360(n366 ,n24[14] ,n69);
    dff g1361(.RN(n1685), .SN(1'b1), .CK(n0), .D(n805), .Q(n20[20]));
    dff g1362(.RN(n1685), .SN(1'b1), .CK(n0), .D(n776), .Q(n24[19]));
    nand g1363(n780 ,n372 ,n505);
    nand g1364(n1190 ,n25[30] ,n1021);
    or g1365(n1640 ,n1352 ,n1586);
    nand g1366(n875 ,n346 ,n583);
    dff g1367(.RN(n1685), .SN(1'b1), .CK(n0), .D(n900), .Q(n10[17]));
    not g1368(n1434 ,n1361);
    or g1369(n1139 ,n682 ,n75);
    nor g1370(n108 ,n6[3] ,n6[2]);
    nand g1371(n1336 ,n967 ,n1055);
    not g1372(n1455 ,n1401);
    nand g1373(n871 ,n222 ,n637);
    nand g1374(n1046 ,n25[6] ,n948);
    dff g1375(.RN(n1685), .SN(1'b1), .CK(n0), .D(n893), .Q(n10[22]));
    nand g1376(n324 ,n24[27] ,n80);
    nand g1377(n1072 ,n28[30] ,n947);
    nand g1378(n779 ,n414 ,n543);
    nor g1379(n257 ,n217 ,n189);
    nand g1380(n883 ,n461 ,n649);
    nand g1381(n1687 ,n33 ,n37);
    nand g1382(n860 ,n458 ,n323);
    nand g1383(n1358 ,n978 ,n1056);
    nand g1384(n748 ,n542 ,n513);
    dff g1385(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1643), .Q(n9[3]));
    nand g1386(n963 ,n30[17] ,n949);
    or g1387(n110 ,n8[3] ,n8[2]);
    nor g1388(n263 ,n217 ,n192);
    not g1389(n1445 ,n1383);
    dff g1390(.RN(n1685), .SN(1'b1), .CK(n0), .D(n901), .Q(n24[8]));
    nand g1391(n811 ,n16[1] ,n464);
    or g1392(n1185 ,n679 ,n79);
    nand g1393(n361 ,n24[6] ,n69);
    nand g1394(n1334 ,n965 ,n1017);
    nand g1395(n753 ,n394 ,n309);
    dff g1396(.RN(n1685), .SN(1'b1), .CK(n0), .D(n721), .Q(n13[20]));
    nand g1397(n686 ,n5[20] ,n220);
    nand g1398(n864 ,n628 ,n533);
    nor g1399(n950 ,n88 ,n938);
    or g1400(n1686 ,n27[6] ,n44);
    nand g1401(n732 ,n484 ,n287);
    dff g1402(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1542), .Q(n28[25]));
    nand g1403(n1512 ,n1231 ,n1103);
    nand g1404(n1555 ,n1299 ,n1093);
    nand g1405(n1267 ,n30[11] ,n79);
    nand g1406(n1524 ,n1244 ,n1115);
    nor g1407(n1712 ,n24[31] ,n24[30]);
    nor g1408(n1599 ,n248 ,n1442);
    nand g1409(n453 ,n1687 ,n84);
    nand g1410(n1514 ,n1233 ,n1105);
    nand g1411(n391 ,n11[4] ,n215);
    nor g1412(n112 ,n4[19] ,n4[18]);
    nand g1413(n1031 ,n22[11] ,n946);
    nor g1414(n244 ,n217 ,n182);
    nand g1415(n746 ,n388 ,n317);
    or g1416(n1623 ,n1318 ,n1569);
    nand g1417(n1535 ,n1253 ,n1125);
    nand g1418(n1276 ,n30[0] ,n1089);
    or g1419(n279 ,n82 ,n199);
    xnor g1420(n230 ,n24[19] ,n20[19]);
    nand g1421(n445 ,n7[0] ,n84);
    nand g1422(n499 ,n11[13] ,n214);
    nand g1423(n1221 ,n25[6] ,n1021);
    nand g1424(n675 ,n5[9] ,n220);
    or g1425(n1167 ,n688 ,n1089);
    nand g1426(n1076 ,n25[28] ,n948);
    nand g1427(n631 ,n8[2] ,n81);
    nand g1428(n1480 ,n1260 ,n1166);
    or g1429(n1635 ,n1342 ,n1581);
    dff g1430(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1696), .Q(n29[6]));
    nand g1431(n972 ,n30[9] ,n949);
    nand g1432(n1585 ,n130 ,n1428);
    nand g1433(n861 ,n502 ,n324);
    dff g1434(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1516), .Q(n22[19]));
    nand g1435(n146 ,n9[25] ,n85);
    nand g1436(n1477 ,n1187 ,n1164);
    not g1437(n909 ,n839);
    dff g1438(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1487), .Q(n30[17]));
    nor g1439(n266 ,n217 ,n195);
    buf g1440(n17[10], n10[2]);
    dff g1441(.RN(n1685), .SN(1'b1), .CK(n0), .D(n874), .Q(n12[16]));
    xnor g1442(n186 ,n24[16] ,n20[16]);
    nand g1443(n410 ,n22[18] ,n83);
    dff g1444(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1634), .Q(n9[12]));
    dff g1445(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1642), .Q(n9[4]));
    nor g1446(n245 ,n217 ,n196);
    or g1447(n284 ,n215 ,n183);
    not g1448(n803 ,n707);
    nor g1449(n1203 ,n90 ,n1022);
    nor g1450(n225 ,n23[2] ,n138);
    nand g1451(n59 ,n29[1] ,n29[0]);
    nand g1452(n983 ,n30[31] ,n949);
    dff g1453(.RN(n1685), .SN(1'b1), .CK(n0), .D(n862), .Q(n12[22]));
    nand g1454(n1000 ,n25[20] ,n948);
    nand g1455(n668 ,n5[2] ,n220);
    nand g1456(n1678 ,n1382 ,n1467);
    nand g1457(n1617 ,n916 ,n1393);
    nand g1458(n545 ,n20[26] ,n73);
    nand g1459(n759 ,n376 ,n403);
    dff g1460(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1565), .Q(n28[2]));
    nand g1461(n713 ,n408 ,n239);
    nand g1462(n899 ,n532 ,n632);
    dff g1463(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1674), .Q(n25[20]));
    nand g1464(n766 ,n630 ,n404);
    nand g1465(n383 ,n11[10] ,n214);
    nand g1466(n401 ,n11[6] ,n214);
    nand g1467(n618 ,n21[3] ,n172);
    nand g1468(n893 ,n512 ,n652);
    dff g1469(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1682), .Q(n25[3]));
    nand g1470(n165 ,n9[3] ,n85);
    nand g1471(n744 ,n383 ,n345);
    buf g1472(n11[26], n10[26]);
    nand g1473(n346 ,n26[1] ,n218);
    dff g1474(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1510), .Q(n22[25]));
    nor g1475(n256 ,n217 ,n188);
    nand g1476(n1683 ,n1394 ,n1620);
    nand g1477(n365 ,n24[9] ,n69);
    dff g1478(.RN(n1685), .SN(1'b1), .CK(n0), .D(n819), .Q(n10[29]));
    nand g1479(n1239 ,n22[16] ,n77);
    or g1480(n1164 ,n692 ,n1089);
    dff g1481(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1561), .Q(n28[6]));
    nand g1482(n63 ,n29[3] ,n62);
    dff g1483(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1625), .Q(n9[21]));
    not g1484(n67 ,n66);
    buf g1485(n14[17], n10[13]);
    nand g1486(n1047 ,n28[6] ,n947);
    not g1487(n1419 ,n1331);
    dff g1488(.RN(n1685), .SN(1'b1), .CK(n0), .D(n868), .Q(n12[19]));
    not g1489(n86 ,n4[2]);
    nor g1490(n298 ,n217 ,n185);
    nand g1491(n961 ,n30[20] ,n949);
    dff g1492(.RN(n1685), .SN(1'b1), .CK(n0), .D(n955), .Q(n23[0]));
    nand g1493(n577 ,n20[2] ,n216);
    nand g1494(n393 ,n11[2] ,n214);
    dff g1495(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1489), .Q(n30[14]));
    dff g1496(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1503), .Q(n30[0]));
    nand g1497(n1318 ,n958 ,n993);
    nand g1498(n1074 ,n22[29] ,n946);
    not g1499(n1450 ,n1391);
    nand g1500(n819 ,n474 ,n650);
    nand g1501(n376 ,n24[29] ,n73);
    buf g1502(n12[4], n10[4]);
    buf g1503(n17[9], n10[1]);
    nand g1504(n627 ,n19[0] ,n73);
    nand g1505(n835 ,n468 ,n657);
    nand g1506(n460 ,n6[1] ,n83);
    nor g1507(n41 ,n27[1] ,n39);
    or g1508(n1160 ,n667 ,n79);
    nand g1509(n1285 ,n30[10] ,n1089);
    nand g1510(n234 ,n222 ,n214);
    nor g1511(n1463 ,n251 ,n1201);
    nand g1512(n1378 ,n5[18] ,n1023);
    nand g1513(n591 ,n20[9] ,n73);
    nand g1514(n387 ,n10[4] ,n82);
    nand g1515(n1303 ,n30[14] ,n79);
    or g1516(n20[1] ,n19[1] ,n1741);
    nand g1517(n822 ,n537 ,n460);
    nand g1518(n937 ,n71 ,n930);
    xnor g1519(n197 ,n24[25] ,n20[25]);
    nor g1520(n259 ,n217 ,n183);
    nand g1521(n49 ,n27[2] ,n48);
    dff g1522(.RN(n1685), .SN(1'b1), .CK(n0), .D(n870), .Q(n18[2]));
    nand g1523(n1061 ,n22[1] ,n946);
    or g1524(n1110 ,n682 ,n1020);
    nand g1525(n508 ,n18[0] ,n215);
    or g1526(n915 ,n115 ,n703);
    nor g1527(n1216 ,n98 ,n1022);
    buf g1528(n12[1], n10[1]);
    nor g1529(n1607 ,n295 ,n1450);
    nand g1530(n152 ,n9[30] ,n85);
    buf g1531(n18[7], n14[7]);
    nand g1532(n805 ,n661 ,n439);
    nand g1533(n317 ,n24[7] ,n216);
    nand g1534(n832 ,n384 ,n344);
    nand g1535(n1271 ,n30[5] ,n79);
    dff g1536(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1518), .Q(n22[17]));
    nor g1537(n1600 ,n254 ,n1443);
    dff g1538(.RN(n1685), .SN(1'b1), .CK(n0), .D(n865), .Q(n12[23]));
    nor g1539(n1739 ,n1727 ,n1738);
    dff g1540(.RN(n1685), .SN(1'b1), .CK(n0), .D(n836), .Q(n20[12]));
    not g1541(n81 ,n82);
    nand g1542(n405 ,n10[2] ,n214);
    nand g1543(n1310 ,n28[2] ,n75);
    nand g1544(n1292 ,n28[18] ,n1019);
    nand g1545(n1311 ,n28[1] ,n75);
    not g1546(n1436 ,n1366);
    nand g1547(n650 ,n20[29] ,n81);
    nand g1548(n625 ,n12[16] ,n82);
    dff g1549(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1553), .Q(n28[13]));
    dff g1550(.RN(n1685), .SN(1'b1), .CK(n0), .D(n731), .Q(n13[10]));
    nand g1551(n587 ,n10[19] ,n82);
    dff g1552(.RN(n1685), .SN(1'b1), .CK(n0), .D(n872), .Q(n12[17]));
    nand g1553(n895 ,n518 ,n648);
    nand g1554(n1080 ,n22[27] ,n946);
    buf g1555(n11[16], n10[16]);
    nand g1556(n613 ,n18[1] ,n214);
    nand g1557(n1259 ,n30[25] ,n79);
    nand g1558(n1542 ,n1284 ,n1092);
    nand g1559(n742 ,n636 ,n277);
    nand g1560(n51 ,n27[3] ,n50);
    nor g1561(n290 ,n205 ,n204);
    nand g1562(n707 ,n222 ,n381);
    nand g1563(n599 ,n13[31] ,n214);
    nand g1564(n1325 ,n1004 ,n1003);
    nand g1565(n458 ,n12[29] ,n215);
    nand g1566(n479 ,n25[27] ,n84);
    not g1567(n1709 ,n24[27]);
    nor g1568(n698 ,n8[0] ,n558);
    nand g1569(n754 ,n396 ,n575);
    nand g1570(n517 ,n10[28] ,n82);
    nand g1571(n481 ,n13[11] ,n82);
    nand g1572(n1505 ,n1213 ,n1095);
    xnor g1573(n196 ,n24[26] ,n20[26]);
    buf g1574(n14[22], n10[18]);
    nand g1575(n1553 ,n1298 ,n1142);
    nand g1576(n1548 ,n1291 ,n1137);
    or g1577(n1116 ,n676 ,n1020);
    dff g1578(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1667), .Q(n25[5]));
    nand g1579(n726 ,n473 ,n281);
    buf g1580(n12[6], n10[6]);
    dff g1581(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1546), .Q(n28[21]));
    nand g1582(n1218 ,n30[22] ,n1089);
    or g1583(n1136 ,n686 ,n1019);
    dff g1584(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1641), .Q(n9[5]));
    dff g1585(.RN(n1685), .SN(1'b1), .CK(n0), .D(n890), .Q(n10[3]));
    nand g1586(n1351 ,n1045 ,n1046);
    nand g1587(n1370 ,n5[26] ,n1023);
    nand g1588(n1680 ,n1387 ,n1469);
    dff g1589(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1658), .Q(n25[25]));
    dff g1590(.RN(n1685), .SN(1'b1), .CK(n0), .D(n828), .Q(n12[28]));
    nor g1591(n1729 ,n1721 ,n1719);
    dff g1592(.RN(n1685), .SN(1'b1), .CK(n0), .D(n762), .Q(n20[29]));
    nor g1593(n1694 ,n48 ,n46);
    buf g1594(n18[10], 1'b0);
    nand g1595(n692 ,n5[26] ,n220);
    nand g1596(n923 ,n222 ,n811);
    or g1597(n1250 ,n675 ,n75);
    nand g1598(n979 ,n30[2] ,n949);
    xnor g1599(n211 ,n20[0] ,n24[0]);
    nand g1600(n905 ,n531 ,n334);
    nand g1601(n492 ,n13[4] ,n215);
    nand g1602(n1350 ,n974 ,n1044);
    not g1603(n45 ,n27[4]);
    nand g1604(n1041 ,n28[8] ,n947);
    nand g1605(n900 ,n626 ,n660);
    nand g1606(n1658 ,n1196 ,n1598);
    nand g1607(n344 ,n24[9] ,n81);
    not g1608(n83 ,n73);
    nand g1609(n1240 ,n22[15] ,n77);
    nand g1610(n437 ,n22[25] ,n84);
    nand g1611(n706 ,n218 ,n308);
    dff g1612(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1552), .Q(n28[15]));
    nand g1613(n962 ,n30[18] ,n949);
    nand g1614(n475 ,n13[14] ,n82);
    nor g1615(n1020 ,n219 ,n950);
    nand g1616(n1309 ,n28[3] ,n1019);
    nand g1617(n1368 ,n5[28] ,n1023);
    nand g1618(n379 ,n24[8] ,n73);
    nand g1619(n1291 ,n28[19] ,n1019);
    nand g1620(n504 ,n14[5] ,n214);
    nand g1621(n316 ,n24[25] ,n80);
    nand g1622(n556 ,n1694 ,n218);
    nand g1623(n840 ,n585 ,n621);
    not g1624(n1435 ,n1363);
    nand g1625(n696 ,n5[30] ,n220);
    dff g1626(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1491), .Q(n30[12]));
    nand g1627(n845 ,n597 ,n603);
    nand g1628(n375 ,n24[28] ,n73);
    buf g1629(n11[17], n10[17]);
    nand g1630(n633 ,n20[16] ,n80);
    nand g1631(n1532 ,n1252 ,n1123);
    nand g1632(n814 ,n351 ,n446);
    nand g1633(n1002 ,n28[20] ,n947);
    nand g1634(n1296 ,n28[15] ,n75);
    nand g1635(n1667 ,n1223 ,n1607);
    nand g1636(n425 ,n13[24] ,n82);
    dff g1637(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1514), .Q(n22[21]));
    nand g1638(n1386 ,n5[10] ,n1023);
    nor g1639(n1597 ,n245 ,n1440);
    nand g1640(n1681 ,n1388 ,n1470);
    dff g1641(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1567), .Q(n28[0]));
    dff g1642(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1560), .Q(n28[7]));
    nor g1643(n1606 ,n265 ,n1449);
    nand g1644(n293 ,n81 ,n172);
    nand g1645(n1263 ,n30[17] ,n1089);
    nand g1646(n417 ,n25[20] ,n83);
    nand g1647(n476 ,n13[13] ,n215);
    dff g1648(.RN(n1685), .SN(1'b1), .CK(n0), .D(n847), .Q(n10[19]));
    nand g1649(n205 ,n107 ,n121);
    not g1650(n1704 ,n24[22]);
    nand g1651(n1669 ,n1234 ,n1609);
    nand g1652(n384 ,n11[9] ,n215);
    nand g1653(n436 ,n25[12] ,n84);
    nor g1654(n262 ,n217 ,n175);
    nand g1655(n1078 ,n28[28] ,n947);
    nand g1656(n519 ,n10[25] ,n215);
    or g1657(n1172 ,n680 ,n79);
    nand g1658(n1018 ,n30[30] ,n949);
    dff g1659(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1476), .Q(n30[27]));
    dff g1660(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1478), .Q(n30[25]));
    or g1661(n1636 ,n1345 ,n1582);
    dff g1662(.RN(n1685), .SN(1'b1), .CK(n0), .D(n790), .Q(n24[11]));
    nand g1663(n1560 ,n1305 ,n1146);
    nand g1664(n970 ,n30[11] ,n949);
    nand g1665(n1256 ,n30[31] ,n1089);
    nand g1666(n484 ,n13[9] ,n215);
    buf g1667(n12[14], n10[14]);
    nand g1668(n1198 ,n25[23] ,n1021);
    nand g1669(n1660 ,n1204 ,n1600);
    nand g1670(n932 ,n225 ,n925);
    or g1671(n1101 ,n691 ,n77);
    nand g1672(n630 ,n20[28] ,n69);
    nand g1673(n892 ,n424 ,n549);
    nand g1674(n958 ,n30[23] ,n949);
    nand g1675(n463 ,n10[15] ,n214);
    dff g1676(.RN(n1685), .SN(1'b1), .CK(n0), .D(n772), .Q(n10[10]));
    nand g1677(n345 ,n24[10] ,n80);
    nand g1678(n867 ,n624 ,n490);
    nor g1679(n1601 ,n298 ,n1444);
    nand g1680(n333 ,n24[21] ,n80);
    nand g1681(n1075 ,n28[29] ,n947);
    nor g1682(n1089 ,n219 ,n954);
    nand g1683(n371 ,n24[16] ,n73);
    dff g1684(.RN(n1685), .SN(1'b1), .CK(n0), .D(n913), .Q(n15[1]));
    or g1685(n270 ,n82 ,n181);
    or g1686(n1112 ,n680 ,n77);
    dff g1687(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1515), .Q(n22[20]));
    nor g1688(n237 ,n217 ,n180);
    nand g1689(n1204 ,n25[18] ,n1021);
    nand g1690(n385 ,n11[8] ,n214);
    nor g1691(n296 ,n217 ,n186);
    nand g1692(n1257 ,n30[29] ,n1089);
    dff g1693(.RN(n1685), .SN(1'b1), .CK(n0), .D(n785), .Q(n24[14]));
    or g1694(n20[0] ,n19[0] ,n1741);
    dff g1695(.RN(n1685), .SN(1'b1), .CK(n0), .D(n888), .Q(n10[4]));
    not g1696(n1421 ,n1335);
    dff g1697(.RN(n1685), .SN(1'b1), .CK(n0), .D(n792), .Q(n20[22]));
    nand g1698(n1682 ,n1227 ,n1619);
    or g1699(n1126 ,n667 ,n77);
    nand g1700(n1069 ,n28[31] ,n947);
    nand g1701(n334 ,n24[14] ,n81);
    not g1702(n942 ,n941);
    not g1703(n1706 ,n24[16]);
    nand g1704(n1661 ,n1205 ,n1601);
    nand g1705(n756 ,n348 ,n398);
    dff g1706(.RN(n1685), .SN(1'b1), .CK(n0), .D(n764), .Q(n24[26]));
    nand g1707(n1249 ,n22[5] ,n1020);
    or g1708(n1648 ,n1400 ,n1611);
    nand g1709(n444 ,n7[1] ,n83);
    or g1710(n1118 ,n674 ,n77);
    nand g1711(n775 ,n545 ,n415);
    nand g1712(n1677 ,n1381 ,n1466);
    nand g1713(n1539 ,n1280 ,n1091);
    nand g1714(n1722 ,n24[5] ,n24[4]);
    dff g1715(.RN(n1685), .SN(1'b1), .CK(n0), .D(n799), .Q(n27[4]));
    dff g1716(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1533), .Q(n22[2]));
    dff g1717(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1671), .Q(n25[24]));
    dff g1718(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1539), .Q(n28[29]));
    xnor g1719(n194 ,n24[6] ,n20[6]);
    nand g1720(n1034 ,n25[10] ,n948);
    or g1721(n1135 ,n687 ,n1019);
    nand g1722(n474 ,n10[29] ,n215);
    nor g1723(n117 ,n4[11] ,n4[10]);
    nand g1724(n153 ,n9[23] ,n85);
    nand g1725(n647 ,n20[0] ,n81);
    nand g1726(n651 ,n20[23] ,n80);
    nand g1727(n580 ,n20[12] ,n73);
    dff g1728(.RN(n1685), .SN(1'b1), .CK(n0), .D(n816), .Q(n10[12]));
    dff g1729(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1666), .Q(n25[6]));
    nand g1730(n1302 ,n28[9] ,n75);
    nand g1731(n467 ,n13[19] ,n214);
    dff g1732(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1631), .Q(n9[15]));
    nand g1733(n1528 ,n1248 ,n1119);
    nand g1734(n426 ,n12[31] ,n82);
    nor g1735(n1598 ,n246 ,n1441);
    buf g1736(n14[8], 1'b0);
    dff g1737(.RN(n1685), .SN(1'b1), .CK(n0), .D(n830), .Q(n20[15]));
    nand g1738(n786 ,n360 ,n432);
    nand g1739(n739 ,n494 ,n294);
    nand g1740(n1475 ,n1188 ,n1162);
    nand g1741(n891 ,n418 ,n546);
    buf g1742(n12[2], n10[2]);
    nand g1743(n886 ,n412 ,n552);
    nand g1744(n655 ,n20[20] ,n216);
    nand g1745(n855 ,n622 ,n480);
    nand g1746(n575 ,n20[26] ,n80);
    nand g1747(n1675 ,n1377 ,n1464);
    nand g1748(n1307 ,n28[5] ,n1019);
    nand g1749(n594 ,n12[18] ,n82);
    nand g1750(n568 ,n1686 ,n218);
    nor g1751(n1471 ,n911 ,n1230);
    nand g1752(n325 ,n24[3] ,n80);
    nand g1753(n1591 ,n167 ,n1434);
    nand g1754(n666 ,n5[0] ,n220);
    dff g1755(.RN(n1685), .SN(1'b1), .CK(n0), .D(n856), .Q(n12[20]));
    nand g1756(n1036 ,n28[9] ,n947);
    nor g1757(n295 ,n217 ,n174);
    nand g1758(n364 ,n24[10] ,n69);
    not g1759(n1438 ,n1368);
    dff g1760(.RN(n1685), .SN(1'b1), .CK(n0), .D(n765), .Q(n24[25]));
    not g1761(n82 ,n216);
    dff g1762(.RN(n1685), .SN(1'b1), .CK(n0), .D(n796), .Q(n27[6]));
    nand g1763(n394 ,n11[1] ,n215);
    nand g1764(n340 ,n24[30] ,n80);
    nand g1765(n1288 ,n28[22] ,n75);
    nand g1766(n656 ,n1691 ,n218);
    nand g1767(n1395 ,n5[1] ,n1023);
    nand g1768(n133 ,n9[14] ,n85);
    not g1769(n1619 ,n1617);
    nand g1770(n1387 ,n5[9] ,n1023);
    buf g1771(n11[30], n10[30]);
    buf g1772(n12[9], n10[9]);
    xnor g1773(n185 ,n24[17] ,n20[17]);
    dff g1774(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1663), .Q(n25[12]));
    nand g1775(n830 ,n566 ,n455);
    nand g1776(n495 ,n12[19] ,n215);
    or g1777(n1120 ,n672 ,n77);
    nor g1778(n945 ,n741 ,n940);
    nand g1779(n222 ,n23[2] ,n128);
    nand g1780(n1363 ,n1063 ,n1064);
    nand g1781(n846 ,n222 ,n610);
    nand g1782(n1065 ,n28[0] ,n947);
    nand g1783(n420 ,n22[19] ,n83);
    or g1784(n1175 ,n676 ,n1089);
    nand g1785(n1032 ,n28[11] ,n947);
    nand g1786(n1244 ,n22[11] ,n1020);
    dff g1787(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1556), .Q(n28[11]));
    nand g1788(n1516 ,n1236 ,n1107);
    not g1789(n1458 ,n1407);
    dff g1790(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1517), .Q(n22[18]));
    nand g1791(n1341 ,n1031 ,n1030);
    dff g1792(.RN(n1685), .SN(1'b1), .CK(n0), .D(n883), .Q(n10[11]));
    nand g1793(n841 ,n588 ,n612);
    nor g1794(n31 ,n29[1] ,n29[0]);
    dff g1795(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1511), .Q(n22[24]));
    nand g1796(n606 ,n15[7] ,n223);
    or g1797(n111 ,n4[1] ,n4[0]);
    nor g1798(n46 ,n27[1] ,n27[0]);
    nand g1799(n1042 ,n25[7] ,n948);
    nand g1800(n327 ,n24[17] ,n216);
    nand g1801(n563 ,n20[28] ,n80);
    nand g1802(n505 ,n25[17] ,n84);
    nand g1803(n1237 ,n22[17] ,n1020);
    nand g1804(n1525 ,n1245 ,n1116);
    nand g1805(n326 ,n24[16] ,n80);
    xnor g1806(n1691 ,n27[4] ,n51);
    nand g1807(n409 ,n25[24] ,n83);
    or g1808(n1642 ,n1356 ,n1588);
    dff g1809(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1483), .Q(n30[20]));
    nand g1810(n1612 ,n150 ,n1455);
    dff g1811(.RN(n1685), .SN(1'b1), .CK(n0), .D(n848), .Q(n12[18]));
    dff g1812(.RN(n1685), .SN(1'b1), .CK(n0), .D(n838), .Q(n10[13]));
    or g1813(n1181 ,n669 ,n1089);
    nor g1814(n925 ,n113 ,n702);
    or g1815(n1173 ,n678 ,n1089);
    nand g1816(n339 ,n24[19] ,n216);
    nand g1817(n590 ,n13[27] ,n215);
    buf g1818(n12[10], n10[10]);
    nand g1819(n1396 ,n5[0] ,n1023);
    xnor g1820(n1699 ,n29[3] ,n61);
    nand g1821(n416 ,n13[1] ,n215);
    nor g1822(n1470 ,n263 ,n1217);
    nand g1823(n525 ,n27[6] ,n217);
    nand g1824(n1264 ,n30[16] ,n79);
    dff g1825(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1538), .Q(n28[30]));
    nand g1826(n1664 ,n1214 ,n1604);
    nor g1827(n129 ,n8[7] ,n8[6]);
    nand g1828(n719 ,n573 ,n276);
    nand g1829(n135 ,n23[1] ,n94);
    nand g1830(n400 ,n22[29] ,n84);
    nand g1831(n1282 ,n28[27] ,n1019);
    nand g1832(n1389 ,n5[7] ,n1023);
    nor g1833(n127 ,n4[15] ,n4[14]);
    nand g1834(n455 ,n22[15] ,n84);
    nor g1835(n1464 ,n253 ,n1203);
    nand g1836(n433 ,n27[2] ,n217);
    nand g1837(n658 ,n21[1] ,n80);
    or g1838(n1147 ,n672 ,n1019);
    nand g1839(n412 ,n10[5] ,n215);
    nand g1840(n969 ,n30[12] ,n949);
    nand g1841(n482 ,n13[10] ,n82);
    dff g1842(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1523), .Q(n22[12]));
    nand g1843(n1656 ,n1192 ,n1595);
    nand g1844(n415 ,n22[26] ,n83);
    nand g1845(n1670 ,n1365 ,n1459);
    nand g1846(n1299 ,n28[12] ,n75);
    nand g1847(n418 ,n10[27] ,n82);
    nand g1848(n1582 ,n154 ,n1425);
    nand g1849(n1508 ,n1222 ,n1099);
    nand g1850(n1068 ,n22[31] ,n946);
    dff g1851(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1479), .Q(n30[24]));
    nor g1852(n1602 ,n259 ,n1445);
    nand g1853(n1369 ,n5[27] ,n1023);
    dff g1854(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1662), .Q(n25[13]));
    nand g1855(n818 ,n311 ,n449);
    nand g1856(n355 ,n26[0] ,n69);
    nand g1857(n676 ,n5[10] ,n220);
    nand g1858(n157 ,n9[27] ,n85);
    nand g1859(n1668 ,n1224 ,n1608);
    nand g1860(n228 ,n104 ,n122);
    nand g1861(n321 ,n24[6] ,n81);
    nand g1862(n620 ,n20[22] ,n69);
    buf g1863(n12[3], n10[3]);
    nand g1864(n1049 ,n22[5] ,n946);
    dff g1865(.RN(n1685), .SN(1'b1), .CK(n0), .D(n735), .Q(n13[6]));
    nor g1866(n1467 ,n257 ,n1208);
    or g1867(n1102 ,n690 ,n77);
    nand g1868(n629 ,n16[3] ,n81);
    nand g1869(n579 ,n22[27] ,n83);
    dff g1870(.RN(n1685), .SN(1'b1), .CK(n0), .D(n843), .Q(n14[0]));
    nand g1871(n984 ,n25[14] ,n948);
    nand g1872(n1404 ,n985 ,n1078);
    nand g1873(n167 ,n9[1] ,n85);
    nand g1874(n1254 ,n22[2] ,n1020);
    nand g1875(n1324 ,n961 ,n1002);
    nand g1876(n308 ,n233 ,n179);
    not g1877(n55 ,n54);
    nand g1878(n757 ,n539 ,n382);
    nand g1879(n1510 ,n1226 ,n1101);
    dff g1880(.RN(n1685), .SN(1'b1), .CK(n0), .D(n897), .Q(n10[18]));
    nand g1881(n381 ,n8[0] ,n225);
    nand g1882(n1082 ,n22[26] ,n946);
    nand g1883(n837 ,n389 ,n540);
    nand g1884(n576 ,n15[2] ,n223);
    nor g1885(n104 ,n4[7] ,n4[6]);
    nand g1886(n359 ,n24[15] ,n69);
    nand g1887(n1496 ,n1269 ,n1177);
    dff g1888(.RN(n1685), .SN(1'b1), .CK(n0), .D(n891), .Q(n10[27]));
    or g1889(n1158 ,n687 ,n1089);
    nand g1890(n783 ,n562 ,n437);
    nand g1891(n1545 ,n1288 ,n1134);
    nand g1892(n1048 ,n25[5] ,n948);
    nand g1893(n1210 ,n22[31] ,n1020);
    nand g1894(n1205 ,n25[17] ,n1021);
    nand g1895(n1657 ,n1195 ,n1597);
    nor g1896(n302 ,n217 ,n190);
    or g1897(n255 ,n1687 ,n69);
    or g1898(n1099 ,n693 ,n77);
    nand g1899(n1287 ,n28[23] ,n75);
    dff g1900(.RN(n1685), .SN(1'b1), .CK(n0), .D(n797), .Q(n27[5]));
    nand g1901(n493 ,n13[3] ,n215);
    dff g1902(.RN(n1685), .SN(1'b1), .CK(n0), .D(n837), .Q(n10[8]));
    dff g1903(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1678), .Q(n25[14]));
    nor g1904(n1206 ,n99 ,n1022);
    nand g1905(n1081 ,n28[27] ,n947);
    nor g1906(n1019 ,n219 ,n952);
    nand g1907(n960 ,n30[21] ,n949);
    not g1908(n76 ,n1020);
    not g1909(n215 ,n216);
    or g1910(n271 ,n214 ,n173);
    nand g1911(n813 ,n349 ,n411);
    nor g1912(n1720 ,n1702 ,n24[2]);
    or g1913(n280 ,n215 ,n231);
    nor g1914(n306 ,n21[2] ,n171);
    nand g1915(n917 ,n614 ,n700);
    dff g1916(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1540), .Q(n28[27]));
    nand g1917(n1214 ,n25[10] ,n1021);
    or g1918(n1153 ,n666 ,n1019);
    nor g1919(n235 ,n221 ,n218);
    nand g1920(n1672 ,n1374 ,n1462);
    nand g1921(n408 ,n13[28] ,n82);
    dff g1922(.RN(n1685), .SN(1'b1), .CK(n0), .D(n724), .Q(n13[17]));
    nand g1923(n1383 ,n5[13] ,n1023);
    nand g1924(n951 ,n2 ,n939);
    nand g1925(n687 ,n5[21] ,n220);
    buf g1926(n11[19], n10[19]);
    or g1927(n282 ,n214 ,n189);
    nand g1928(n1343 ,n1033 ,n1034);
    or g1929(n1091 ,n695 ,n75);
    nand g1930(n684 ,n5[18] ,n220);
    nand g1931(n1486 ,n1193 ,n1170);
    nand g1932(n1671 ,n1372 ,n1460);
    nand g1933(n1044 ,n28[7] ,n947);
    dff g1934(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1621), .Q(n9[25]));
    nand g1935(n1521 ,n1241 ,n1112);
    nand g1936(n1236 ,n22[19] ,n77);
    dff g1937(.RN(n1685), .SN(1'b1), .CK(n0), .D(n895), .Q(n10[24]));
    or g1938(n1093 ,n678 ,n1019);
    nand g1939(n1511 ,n1229 ,n1102);
    dff g1940(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1505), .Q(n22[30]));
    dff g1941(.RN(n1685), .SN(1'b1), .CK(n0), .D(n786), .Q(n24[13]));
    nand g1942(n1390 ,n5[6] ,n1023);
    nand g1943(n1354 ,n976 ,n1050);
    or g1944(n1105 ,n687 ,n77);
    nand g1945(n1227 ,n25[3] ,n1021);
    or g1946(n1163 ,n693 ,n79);
    not g1947(n1456 ,n1403);
    dff g1948(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1676), .Q(n25[16]));
    nand g1949(n792 ,n620 ,n485);
    not g1950(n1440 ,n1370);
    or g1951(n1176 ,n674 ,n1089);
    nand g1952(n208 ,n120 ,n126);
    nand g1953(n389 ,n10[8] ,n215);
    nand g1954(n527 ,n12[23] ,n82);
    nand g1955(n423 ,n22[24] ,n83);
    nand g1956(n1284 ,n28[25] ,n1019);
    nand g1957(n1569 ,n153 ,n1411);
    not g1958(n214 ,n81);
    nand g1959(n703 ,n125 ,n305);
    nand g1960(n404 ,n22[28] ,n83);
    nand g1961(n1345 ,n971 ,n1035);
    or g1962(n1149 ,n670 ,n75);
    nand g1963(n842 ,n443 ,n318);
    nand g1964(n1247 ,n22[8] ,n1020);
    dff g1965(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1500), .Q(n30[3]));
    nand g1966(n876 ,n222 ,n572);
    nand g1967(n1030 ,n25[11] ,n948);
    dff g1968(.RN(n1685), .SN(1'b1), .CK(n0), .D(n861), .Q(n12[27]));
    nand g1969(n659 ,n20[4] ,n80);
    nand g1970(n1726 ,n24[7] ,n1708);
    dff g1971(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1501), .Q(n30[2]));
    or g1972(n1638 ,n1348 ,n1584);
    nand g1973(n1262 ,n30[19] ,n1089);
    dff g1974(.RN(n1685), .SN(1'b1), .CK(n0), .D(n714), .Q(n13[27]));
    nand g1975(n1057 ,n22[2] ,n946);
    nand g1976(n558 ,n8[1] ,n225);
    nand g1977(n501 ,n25[16] ,n84);
    nand g1978(n550 ,n20[23] ,n69);
    nand g1979(n1219 ,n22[28] ,n1020);
    or g1980(n297 ,n82 ,n185);
    nand g1981(n897 ,n605 ,n589);
    nand g1982(n1380 ,n5[16] ,n1023);
    nand g1983(n1375 ,n5[21] ,n1023);
    nor g1984(n1593 ,n242 ,n1436);
    or g1985(n1170 ,n684 ,n79);
    or g1986(n69 ,n94 ,n137);
    nand g1987(n490 ,n22[1] ,n83);
    nand g1988(n356 ,n24[18] ,n73);
    not g1989(n1411 ,n1317);
    nand g1990(n1401 ,n1074 ,n1073);
    nand g1991(n1314 ,n956 ,n1085);
    nand g1992(n977 ,n30[4] ,n949);
    or g1993(n1113 ,n679 ,n1020);
    nand g1994(n1583 ,n163 ,n1426);
    nand g1995(n991 ,n25[23] ,n948);
    nand g1996(n907 ,n536 ,n322);
    buf g1997(n14[10], 1'b0);
    nand g1998(n1653 ,n1190 ,n1593);
    nand g1999(n820 ,n560 ,n452);
    nand g2000(n1241 ,n22[14] ,n77);
    or g2001(n1119 ,n673 ,n1020);
    nand g2002(n134 ,n9[2] ,n85);
    or g2003(n913 ,n876 ,n875);
    dff g2004(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1535), .Q(n22[0]));
    dff g2005(.RN(n1685), .SN(1'b1), .CK(n0), .D(n944), .Q(n23[1]));
    buf g2006(n14[26], n10[22]);
    or g2007(n1122 ,n670 ,n1020);
    nand g2008(n714 ,n590 ,n272);
    nor g2009(n946 ,n85 ,n938);
    dff g2010(.RN(n1685), .SN(1'b1), .CK(n0), .D(n742), .Q(n15[5]));
    nand g2011(n807 ,n358 ,n444);
    nand g2012(n461 ,n10[11] ,n82);
    xnor g2013(n1695 ,n68 ,n29[7]);
    nand g2014(n430 ,n25[14] ,n84);
    dff g2015(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1652), .Q(n25[1]));
    nand g2016(n1289 ,n28[21] ,n1019);
    nor g2017(n105 ,n4[27] ,n4[26]);
    nand g2018(n906 ,n499 ,n332);
    nand g2019(n462 ,n22[13] ,n83);
    nand g2020(n1574 ,n131 ,n1416);
    dff g2021(.RN(n1685), .SN(1'b1), .CK(n0), .D(n760), .Q(n24[28]));
    dff g2022(.RN(n1685), .SN(1'b1), .CK(n0), .D(n771), .Q(n24[22]));
    dff g2023(.RN(n1685), .SN(1'b1), .CK(n0), .D(n754), .Q(n10[26]));
    dff g2024(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1481), .Q(n30[22]));
    nand g2025(n995 ,n25[22] ,n948);
    nand g2026(n1187 ,n30[26] ,n1089);
    dff g2027(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1651), .Q(n9[26]));
    nand g2028(n833 ,n463 ,n639);
    dff g2029(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1499), .Q(n30[4]));
    dff g2030(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1562), .Q(n28[5]));
    nand g2031(n812 ,n16[0] ,n464);
    nand g2032(n856 ,n497 ,n338);
    nor g2033(n912 ,n268 ,n706);
    nand g2034(n155 ,n9[5] ,n85);
    nand g2035(n785 ,n366 ,n430);
    xnor g2036(n173 ,n24[29] ,n20[29]);
    buf g2037(n11[29], n10[29]);
    not g2038(n1454 ,n1398);
    nand g2039(n1260 ,n30[23] ,n1089);
    dff g2040(.RN(n1685), .SN(1'b1), .CK(n0), .D(n761), .Q(n10[2]));
    or g2041(n115 ,n15[4] ,n15[5]);
    nand g2042(n1659 ,n1198 ,n1599);
    nand g2043(n878 ,n347 ,n640);
    nand g2044(n1316 ,n957 ,n990);
    nand g2045(n1561 ,n1306 ,n1147);
    nor g2046(n218 ,n23[2] ,n135);
    nor g2047(n931 ,n224 ,n925);
    or g2048(n1177 ,n673 ,n1089);
    nand g2049(n1526 ,n1246 ,n1117);
    or g2050(n269 ,n215 ,n180);
    nand g2051(n1313 ,n30[30] ,n1089);
    or g2052(n1141 ,n680 ,n75);
    nand g2053(n681 ,n5[31] ,n220);
    or g2054(n1132 ,n690 ,n75);
    nand g2055(n667 ,n5[1] ,n220);
    or g2056(n1133 ,n689 ,n1019);
    dff g2057(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1679), .Q(n25[11]));
    nand g2058(n641 ,n20[7] ,n81);
    nand g2059(n648 ,n20[24] ,n80);
    nand g2060(n903 ,n506 ,n633);
    dff g2061(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1494), .Q(n30[9]));
    nand g2062(n1029 ,n28[12] ,n947);
    or g2063(n1107 ,n685 ,n77);
    not g2064(n73 ,n84);
    nand g2065(n999 ,n28[21] ,n947);
    nand g2066(n990 ,n28[24] ,n947);
    nand g2067(n1587 ,n155 ,n1430);
    not g2068(n1448 ,n1389);
    nor g2069(n1189 ,n95 ,n1022);
    nand g2070(n1367 ,n5[29] ,n1023);
    nand g2071(n145 ,n9[24] ,n85);
    nand g2072(n1013 ,n22[16] ,n946);
    dff g2073(.RN(n1685), .SN(1'b1), .CK(n0), .D(n844), .Q(n20[9]));
    buf g2074(n14[24], n10[20]);
    nor g2075(n1217 ,n92 ,n1022);
    nand g2076(n584 ,n22[6] ,n84);
    not g2077(n1431 ,n1355);
    nor g2078(n72 ,n4[1] ,n4[0]);
    nand g2079(n511 ,n22[12] ,n83);
    nand g2080(n993 ,n28[23] ,n947);
    nand g2081(n679 ,n5[13] ,n220);
    nand g2082(n933 ,n80 ,n915);
    nand g2083(n774 ,n451 ,n663);
    nand g2084(n1275 ,n30[1] ,n1089);
    nand g2085(n592 ,n22[7] ,n84);
    dff g2086(.RN(n1685), .SN(1'b1), .CK(n0), .D(n736), .Q(n13[5]));
    nand g2087(n56 ,n27[6] ,n55);
    nand g2088(n315 ,n26[0] ,n216);
    nand g2089(n902 ,n514 ,n548);
    buf g2090(n17[8], n10[0]);
    dff g2091(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1670), .Q(n25[31]));
    nand g2092(n1060 ,n25[1] ,n948);
    nand g2093(n396 ,n10[26] ,n215);
    nand g2094(n643 ,n20[21] ,n80);
    or g2095(n1128 ,n696 ,n75);
    nand g2096(n1500 ,n1273 ,n1181);
    not g2097(n1422 ,n1337);
    nand g2098(n1507 ,n1219 ,n1097);
    nand g2099(n794 ,n553 ,n623);
    nand g2100(n570 ,n20[14] ,n73);
    buf g2101(n14[31], n10[27]);
    dff g2102(.RN(n1685), .SN(1'b1), .CK(n0), .D(n885), .Q(n12[25]));
    buf g2103(n11[22], n10[22]);
    nor g2104(n261 ,n217 ,n191);
    nor g2105(n120 ,n4[31] ,n4[30]);
    nand g2106(n637 ,n15[4] ,n223);
    dff g2107(.RN(n1685), .SN(1'b1), .CK(n0), .D(n747), .Q(n11[6]));
    not g2108(n1702 ,n24[3]);
    nand g2109(n1293 ,n28[17] ,n75);
    nand g2110(n849 ,n602 ,n592);
    or g2111(n1626 ,n1324 ,n1572);
    nor g2112(n924 ,n226 ,n802);
    dff g2113(.RN(n1685), .SN(1'b1), .CK(n0), .D(n826), .Q(n12[30]));
    or g2114(n1114 ,n678 ,n1020);
    xnor g2115(n177 ,n24[11] ,n20[11]);
    dff g2116(.RN(n1685), .SN(1'b1), .CK(n0), .D(n880), .Q(n18[0]));
    not g2117(n1443 ,n1378);
    nand g2118(n1402 ,n982 ,n1075);
    nand g2119(n615 ,n20[4] ,n73);
    nand g2120(n529 ,n6[2] ,n84);
    nor g2121(n248 ,n217 ,n232);
    nand g2122(n638 ,n16[2] ,n216);
    nand g2123(n1026 ,n28[13] ,n947);
    nand g2124(n788 ,n362 ,n436);
    nand g2125(n976 ,n30[5] ,n949);
    nand g2126(n369 ,n24[24] ,n73);
    nand g2127(n533 ,n6[3] ,n84);
    nand g2128(n1012 ,n25[16] ,n948);
    nand g2129(n549 ,n20[1] ,n216);
    nand g2130(n534 ,n11[12] ,n215);
    or g2131(n1180 ,n670 ,n79);
    nand g2132(n964 ,n30[16] ,n949);
    nand g2133(n378 ,n24[7] ,n69);
    nand g2134(n486 ,n22[0] ,n83);
    nand g2135(n1294 ,n30[12] ,n79);
    not g2136(n1412 ,n1319);
    nand g2137(n1393 ,n5[3] ,n1023);
    nand g2138(n454 ,n10[3] ,n214);
    nand g2139(n1261 ,n30[21] ,n79);
    dff g2140(.RN(n1685), .SN(1'b1), .CK(n0), .D(n867), .Q(n19[1]));
    dff g2141(.RN(n1685), .SN(1'b1), .CK(n0), .D(n845), .Q(n20[8]));
    nand g2142(n1090 ,n22[6] ,n77);
    dff g2143(.RN(n1685), .SN(1'b1), .CK(n0), .D(n769), .Q(n20[27]));
    dff g2144(.RN(n1685), .SN(1'b1), .CK(n0), .D(n734), .Q(n13[7]));
    nand g2145(n1253 ,n22[0] ,n1020);
    nand g2146(n602 ,n20[7] ,n73);
    dff g2147(.RN(n1685), .SN(1'b1), .CK(n0), .D(n906), .Q(n11[13]));
    dff g2148(.RN(n1685), .SN(1'b1), .CK(n0), .D(n831), .Q(n20[13]));
    xnor g2149(n801 ,n217 ,n27[0]);
    dff g2150(.RN(n1685), .SN(1'b1), .CK(n0), .D(n884), .Q(n10[23]));
    nand g2151(n1522 ,n1242 ,n1113);
    nand g2152(n1403 ,n1077 ,n1076);
    nor g2153(n128 ,n94 ,n23[1]);
    buf g2154(n17[2], n14[6]);
    dff g2155(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1668), .Q(n25[4]));
    nand g2156(n1056 ,n28[3] ,n947);
    nand g2157(n642 ,n20[13] ,n80);
    nand g2158(n377 ,n24[30] ,n73);
    dff g2159(.RN(n1685), .SN(1'b1), .CK(n0), .D(n794), .Q(n20[21]));
    buf g2160(n17[15], n10[7]);
    dff g2161(.RN(n1685), .SN(1'b1), .CK(n0), .D(n1524), .Q(n22[11]));
    nor g2162(n254 ,n217 ,n231);
    nand g2163(n516 ,n10[23] ,n82);
    nand g2164(n1278 ,n28[30] ,n1019);
    nand g2165(n600 ,n20[19] ,n216);
endmodule
