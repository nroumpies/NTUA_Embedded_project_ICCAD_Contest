module top (n0, n1, n2, n3, n4, n5, n13, n17, n18, n6, n7, n14, n19, n20, n8, n9, n15, n21, n22, n10, n11, n16, n23, n24, n12, n25, n26, n27, n28, n29, n30, n31, n32, n34, n33);
    input n0, n1;
    input [3:0] n2, n3;
    input [31:0] n4, n5, n6, n7, n8, n9, n10, n11, n12;
    input [15:0] n13, n14, n15, n16;
    input [1:0] n17, n18, n19, n20, n21, n22, n23, n24;
    output [31:0] n25, n26;
    output n27, n28;
    output [3:0] n29, n30;
    output [7:0] n31, n32, n33;
    output [15:0] n34;
    wire n0, n1;
    wire [3:0] n2, n3;
    wire [31:0] n4, n5, n6, n7, n8, n9, n10, n11, n12;
    wire [15:0] n13, n14, n15, n16;
    wire [1:0] n17, n18, n19, n20, n21, n22, n23, n24;
    wire [31:0] n25, n26;
    wire n27, n28;
    wire [3:0] n29, n30;
    wire [7:0] n31, n32, n33;
    wire [15:0] n34;
    wire [3:0] n35;
    wire [3:0] n36;
    wire [3:0] n37;
    wire [3:0] n38;
    wire [3:0] n39;
    wire [31:0] n40;
    wire [15:0] n41;
    wire [31:0] n42;
    wire [2:0] n43;
    wire [1:0] n44;
    wire [2:0] n45;
    wire [31:0] n46;
    wire [31:0] n47;
    wire [31:0] n48;
    wire [31:0] n49;
    wire [15:0] n50;
    wire [15:0] n51;
    wire [15:0] n52;
    wire [15:0] n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171, n172, n173;
    wire n174, n175, n176, n177, n178, n179, n180, n181;
    wire n182, n183, n184, n185, n186, n187, n188, n189;
    wire n190, n191, n192, n193, n194, n195, n196, n197;
    wire n198, n199, n200, n201, n202, n203, n204, n205;
    wire n206, n207, n208, n209, n210, n211, n212, n213;
    wire n214, n215, n216, n217, n218, n219, n220, n221;
    wire n222, n223, n224, n225, n226, n227, n228, n229;
    wire n230, n231, n232, n233, n234, n235, n236, n237;
    wire n238, n239, n240, n241, n242, n243, n244, n245;
    wire n246, n247, n248, n249, n250, n251, n252, n253;
    wire n254, n255, n256, n257, n258, n259, n260, n261;
    wire n262, n263, n264, n265, n266, n267, n268, n269;
    wire n270, n271, n272, n273, n274, n275, n276, n277;
    wire n278, n279, n280, n281, n282, n283, n284, n285;
    wire n286, n287, n288, n289, n290, n291, n292, n293;
    wire n294, n295, n296, n297, n298, n299, n300, n301;
    wire n302, n303, n304, n305, n306, n307, n308, n309;
    wire n310, n311, n312, n313, n314, n315, n316, n317;
    wire n318, n319, n320, n321, n322, n323, n324, n325;
    wire n326, n327, n328, n329, n330, n331, n332, n333;
    wire n334, n335, n336, n337, n338, n339, n340, n341;
    wire n342, n343, n344, n345, n346, n347, n348, n349;
    wire n350, n351, n352, n353, n354, n355, n356, n357;
    wire n358, n359, n360, n361, n362, n363, n364, n365;
    wire n366, n367, n368, n369, n370, n371, n372, n373;
    wire n374, n375, n376, n377, n378, n379, n380, n381;
    wire n382, n383, n384, n385, n386, n387, n388, n389;
    wire n390, n391, n392, n393, n394, n395, n396, n397;
    wire n398, n399, n400, n401, n402, n403, n404, n405;
    wire n406, n407, n408, n409, n410, n411, n412, n413;
    wire n414, n415, n416, n417, n418, n419, n420, n421;
    wire n422, n423, n424, n425, n426, n427, n428, n429;
    wire n430, n431, n432, n433, n434, n435, n436, n437;
    wire n438, n439, n440, n441, n442, n443, n444, n445;
    wire n446, n447, n448, n449, n450, n451, n452, n453;
    wire n454, n455, n456, n457, n458, n459, n460, n461;
    wire n462, n463, n464, n465, n466, n467, n468, n469;
    wire n470, n471, n472, n473, n474, n475, n476, n477;
    wire n478, n479, n480, n481, n482, n483, n484, n485;
    wire n486, n487, n488, n489, n490, n491, n492, n493;
    wire n494, n495, n496, n497, n498, n499, n500, n501;
    wire n502, n503, n504, n505, n506, n507, n508, n509;
    wire n510, n511, n512, n513, n514, n515, n516, n517;
    wire n518, n519, n520, n521, n522, n523, n524, n525;
    wire n526, n527, n528, n529, n530, n531, n532, n533;
    wire n534, n535, n536, n537, n538, n539, n540, n541;
    wire n542, n543, n544, n545, n546, n547, n548, n549;
    wire n550, n551, n552, n553, n554, n555, n556, n557;
    wire n558, n559, n560, n561, n562, n563, n564, n565;
    wire n566, n567, n568, n569, n570, n571, n572, n573;
    wire n574, n575, n576, n577, n578, n579, n580, n581;
    wire n582, n583, n584, n585, n586, n587, n588, n589;
    wire n590, n591, n592, n593, n594, n595, n596, n597;
    wire n598, n599, n600, n601, n602, n603, n604, n605;
    wire n606, n607, n608, n609, n610, n611, n612, n613;
    wire n614, n615, n616, n617, n618, n619, n620, n621;
    wire n622, n623, n624, n625, n626, n627, n628, n629;
    wire n630, n631, n632, n633, n634, n635, n636, n637;
    wire n638, n639, n640, n641, n642, n643, n644, n645;
    wire n646, n647, n648, n649, n650, n651, n652, n653;
    wire n654, n655, n656, n657, n658, n659, n660, n661;
    wire n662, n663, n664, n665, n666, n667, n668, n669;
    wire n670, n671, n672, n673, n674, n675, n676, n677;
    wire n678, n679, n680, n681, n682, n683, n684, n685;
    wire n686, n687, n688, n689, n690, n691, n692, n693;
    wire n694, n695, n696, n697, n698, n699, n700, n701;
    wire n702, n703, n704, n705, n706, n707, n708, n709;
    wire n710, n711, n712, n713, n714, n715, n716, n717;
    wire n718, n719, n720, n721, n722, n723, n724, n725;
    wire n726, n727, n728, n729, n730, n731, n732, n733;
    wire n734, n735, n736, n737, n738, n739, n740, n741;
    wire n742, n743, n744, n745, n746, n747, n748, n749;
    wire n750, n751, n752, n753, n754, n755, n756, n757;
    wire n758, n759, n760, n761, n762, n763, n764, n765;
    wire n766, n767, n768, n769, n770, n771, n772, n773;
    wire n774, n775, n776, n777, n778, n779, n780, n781;
    wire n782, n783, n784, n785, n786, n787, n788, n789;
    wire n790, n791, n792, n793, n794, n795, n796, n797;
    wire n798, n799, n800, n801, n802, n803, n804, n805;
    wire n806, n807, n808, n809, n810, n811, n812, n813;
    wire n814, n815, n816, n817, n818, n819, n820, n821;
    wire n822, n823, n824, n825, n826, n827, n828, n829;
    wire n830, n831, n832, n833, n834, n835, n836, n837;
    wire n838, n839, n840, n841, n842, n843, n844, n845;
    wire n846, n847, n848, n849, n850, n851, n852, n853;
    wire n854, n855, n856, n857, n858, n859, n860, n861;
    wire n862, n863, n864, n865, n866, n867, n868, n869;
    wire n870, n871, n872, n873, n874, n875, n876, n877;
    wire n878, n879, n880, n881, n882, n883, n884, n885;
    wire n886, n887, n888, n889, n890, n891, n892, n893;
    wire n894, n895, n896, n897, n898, n899, n900, n901;
    wire n902, n903, n904, n905, n906, n907, n908, n909;
    wire n910, n911, n912, n913, n914, n915, n916, n917;
    wire n918, n919, n920, n921, n922, n923, n924, n925;
    wire n926, n927, n928, n929, n930, n931, n932, n933;
    wire n934, n935, n936, n937, n938, n939, n940, n941;
    wire n942, n943, n944, n945, n946, n947, n948, n949;
    wire n950, n951, n952, n953, n954, n955, n956, n957;
    wire n958, n959, n960, n961, n962, n963, n964, n965;
    wire n966, n967, n968, n969, n970, n971, n972, n973;
    wire n974, n975, n976, n977, n978, n979, n980, n981;
    wire n982, n983, n984, n985, n986, n987, n988, n989;
    wire n990, n991, n992, n993, n994, n995, n996, n997;
    wire n998, n999, n1000, n1001, n1002, n1003, n1004, n1005;
    wire n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013;
    wire n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
    wire n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
    wire n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
    wire n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;
    wire n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053;
    wire n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061;
    wire n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069;
    wire n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077;
    wire n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085;
    wire n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093;
    wire n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101;
    wire n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109;
    wire n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117;
    wire n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125;
    wire n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133;
    wire n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141;
    wire n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149;
    wire n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157;
    wire n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165;
    wire n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173;
    wire n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181;
    wire n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189;
    wire n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197;
    wire n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205;
    wire n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
    wire n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221;
    wire n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229;
    wire n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237;
    wire n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245;
    wire n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253;
    wire n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261;
    wire n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269;
    wire n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277;
    wire n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285;
    wire n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293;
    wire n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301;
    wire n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309;
    wire n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;
    wire n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325;
    wire n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333;
    wire n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;
    wire n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349;
    wire n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;
    wire n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365;
    wire n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373;
    wire n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381;
    wire n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389;
    wire n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397;
    wire n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405;
    wire n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413;
    wire n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421;
    wire n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429;
    wire n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437;
    wire n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445;
    wire n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453;
    wire n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461;
    wire n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469;
    wire n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477;
    wire n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485;
    wire n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493;
    wire n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501;
    wire n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509;
    wire n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517;
    wire n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525;
    wire n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533;
    wire n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541;
    wire n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
    wire n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557;
    wire n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565;
    wire n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573;
    wire n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581;
    wire n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589;
    wire n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597;
    wire n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605;
    wire n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613;
    wire n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621;
    wire n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629;
    wire n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637;
    wire n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645;
    wire n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653;
    wire n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661;
    wire n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669;
    wire n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677;
    wire n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685;
    wire n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693;
    wire n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701;
    wire n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709;
    wire n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717;
    wire n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725;
    wire n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733;
    wire n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741;
    wire n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749;
    wire n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757;
    wire n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765;
    wire n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773;
    wire n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781;
    wire n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789;
    wire n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797;
    wire n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805;
    wire n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813;
    wire n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821;
    wire n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829;
    wire n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837;
    wire n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845;
    wire n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853;
    wire n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861;
    wire n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869;
    wire n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877;
    wire n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885;
    wire n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893;
    wire n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901;
    wire n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909;
    wire n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917;
    wire n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925;
    wire n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933;
    wire n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941;
    wire n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949;
    wire n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957;
    wire n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965;
    wire n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973;
    wire n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981;
    wire n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989;
    wire n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997;
    wire n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005;
    wire n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013;
    wire n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021;
    wire n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029;
    wire n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037;
    wire n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045;
    wire n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053;
    wire n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061;
    wire n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069;
    wire n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077;
    wire n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085;
    wire n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093;
    wire n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101;
    wire n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109;
    wire n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117;
    wire n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125;
    wire n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133;
    wire n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141;
    wire n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149;
    wire n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157;
    wire n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165;
    wire n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173;
    wire n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181;
    wire n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189;
    wire n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197;
    wire n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205;
    wire n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213;
    wire n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221;
    wire n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229;
    wire n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237;
    wire n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245;
    wire n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253;
    wire n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261;
    wire n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269;
    wire n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277;
    wire n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285;
    wire n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293;
    wire n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301;
    wire n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309;
    wire n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317;
    wire n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325;
    wire n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333;
    wire n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341;
    wire n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349;
    wire n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357;
    wire n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365;
    wire n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373;
    wire n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381;
    wire n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389;
    wire n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397;
    wire n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405;
    wire n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413;
    wire n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421;
    wire n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429;
    wire n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437;
    wire n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445;
    wire n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453;
    wire n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461;
    wire n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469;
    wire n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477;
    wire n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485;
    wire n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493;
    wire n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501;
    wire n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509;
    wire n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517;
    wire n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525;
    wire n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533;
    wire n2534, n2535;
    or g0(n402 ,n323 ,n52[11]);
    nand g1(n2278 ,n1979 ,n2100);
    dff g2(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2336), .Q(n50[12]));
    xnor g3(n2517 ,n34[15] ,n288);
    nand g4(n1106 ,n818 ,n786);
    nor g5(n2418 ,n2396 ,n2408);
    nand g6(n655 ,n2529 ,n523);
    xnor g7(n2510 ,n50[10] ,n107);
    nand g8(n1509 ,n953 ,n1034);
    not g9(n2150 ,n2037);
    nor g10(n1696 ,n670 ,n1398);
    nand g11(n710 ,n2447 ,n528);
    nand g12(n1092 ,n7[7] ,n295);
    nand g13(n93 ,n50[1] ,n50[0]);
    nand g14(n1742 ,n1135 ,n1382);
    not g15(n339 ,n47[0]);
    not g16(n119 ,n51[12]);
    nand g17(n1323 ,n37[0] ,n1142);
    nand g18(n1436 ,n42[5] ,n292);
    nand g19(n1367 ,n1119 ,n1010);
    nand g20(n607 ,n339 ,n526);
    not g21(n1147 ,n1099);
    nand g22(n1656 ,n1132 ,n1421);
    nand g23(n1494 ,n944 ,n1238);
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n896), .Q(n47[6]));
    not g25(n146 ,n52[8]);
    nand g26(n102 ,n50[6] ,n101);
    nand g27(n2061 ,n2484 ,n1696);
    nand g28(n1720 ,n42[27] ,n289);
    nand g29(n1429 ,n42[9] ,n1139);
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2363), .Q(n52[2]));
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1587), .Q(n30[0]));
    nand g32(n1136 ,n8[26] ,n300);
    nand g33(n1505 ,n1261 ,n1036);
    nor g34(n394 ,n327 ,n53[7]);
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n888), .Q(n48[5]));
    nand g36(n2366 ,n2061 ,n2303);
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2228), .Q(n26[30]));
    nand g38(n1797 ,n1204 ,n1466);
    nor g39(n55 ,n54 ,n2419);
    nand g40(n652 ,n47[2] ,n587);
    not g41(n115 ,n114);
    xnor g42(n2446 ,n47[9] ,n230);
    nand g43(n2217 ,n50[10] ,n1992);
    nand g44(n2054 ,n2493 ,n1701);
    nor g45(n526 ,n2533 ,n487);
    nand g46(n2118 ,n27 ,n1704);
    xnor g47(n2499 ,n51[14] ,n142);
    nor g48(n134 ,n51[9] ,n133);
    xnor g49(n2428 ,n49[9] ,n260);
    or g50(n1899 ,n1797 ,n1821);
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2211), .Q(n26[0]));
    nand g52(n1301 ,n41[15] ,n1139);
    nand g53(n228 ,n47[7] ,n226);
    nand g54(n1808 ,n1234 ,n1489);
    nand g55(n1990 ,n25[6] ,n1693);
    nor g56(n381 ,n314 ,n52[5]);
    nand g57(n2053 ,n1643 ,n1642);
    nor g58(n382 ,n320 ,n51[15]);
    nor g59(n127 ,n51[5] ,n126);
    nor g60(n1361 ,n2407 ,n1156);
    nand g61(n1334 ,n40[11] ,n292);
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1883), .Q(n41[13]));
    xnor g63(n2421 ,n49[2] ,n248);
    nand g64(n2105 ,n12[12] ,n1694);
    nand g65(n2351 ,n1994 ,n2288);
    nand g66(n579 ,n441 ,n416);
    nor g67(n494 ,n361 ,n398);
    nand g68(n1332 ,n40[12] ,n1139);
    not g69(n1540 ,n1458);
    nand g70(n1498 ,n40[15] ,n1139);
    nand g71(n1711 ,n40[31] ,n291);
    nand g72(n2066 ,n2479 ,n1696);
    nand g73(n1732 ,n1110 ,n1358);
    nand g74(n1282 ,n8[22] ,n299);
    not g75(n2146 ,n2028);
    nand g76(n752 ,n34[7] ,n524);
    or g77(n362 ,n332 ,n41[0]);
    nand g78(n1100 ,n813 ,n781);
    nand g79(n747 ,n2430 ,n530);
    nand g80(n2099 ,n12[18] ,n1694);
    nand g81(n650 ,n47[4] ,n587);
    nand g82(n1643 ,n40[2] ,n291);
    nand g83(n1706 ,n1235 ,n1555);
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2227), .Q(n26[31]));
    nor g85(n422 ,n336 ,n41[3]);
    not g86(n2134 ,n2003);
    nand g87(n2378 ,n2059 ,n2316);
    nand g88(n792 ,n638 ,n604);
    xnor g89(n2484 ,n52[14] ,n170);
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n891), .Q(n48[3]));
    nand g91(n1241 ,n8[2] ,n299);
    nor g92(n2381 ,n1398 ,n2380);
    nand g93(n1492 ,n40[18] ,n292);
    nand g94(n1942 ,n2463 ,n1698);
    nor g95(n284 ,n263 ,n283);
    nand g96(n626 ,n479 ,n542);
    nand g97(n426 ,n50[8] ,n319);
    nand g98(n2055 ,n1644 ,n1645);
    nand g99(n1691 ,n914 ,n1540);
    nand g100(n1709 ,n950 ,n1560);
    nand g101(n1777 ,n1083 ,n1443);
    nand g102(n1449 ,n1223 ,n1064);
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2361), .Q(n53[4]));
    nand g104(n2202 ,n2039 ,n2151);
    nand g105(n1743 ,n1137 ,n1384);
    or g106(n1902 ,n1803 ,n1818);
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1899), .Q(n40[30]));
    nor g108(n527 ,n2407 ,n476);
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2271), .Q(n25[10]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1929), .Q(n36[1]));
    nand g111(n1105 ,n817 ,n785);
    nand g112(n608 ,n38[0] ,n532);
    nor g113(n353 ,n43[0] ,n43[1]);
    not g114(n1829 ,n1737);
    nor g115(n84 ,n49[4] ,n49[3]);
    not g116(n124 ,n123);
    nand g117(n2035 ,n26[11] ,n1695);
    nand g118(n555 ,n463 ,n373);
    nand g119(n1629 ,n42[8] ,n289);
    nand g120(n1632 ,n40[7] ,n1397);
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2179), .Q(n40[7]));
    nor g122(n538 ,n38[2] ,n479);
    nand g123(n940 ,n11[21] ,n294);
    or g124(n379 ,n326 ,n50[12]);
    nand g125(n1768 ,n35[3] ,n1399);
    nand g126(n2275 ,n1982 ,n2103);
    nand g127(n639 ,n38[3] ,n532);
    or g128(n1568 ,n1317 ,n974);
    nand g129(n1297 ,n985 ,n984);
    nor g130(n595 ,n575 ,n581);
    not g131(n321 ,n41[10]);
    nand g132(n2215 ,n50[12] ,n1992);
    not g133(n261 ,n34[4]);
    nand g134(n1686 ,n1167 ,n1535);
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2354), .Q(n53[11]));
    nand g136(n495 ,n360 ,n399);
    nand g137(n203 ,n46[1] ,n46[0]);
    nand g138(n1291 ,n308 ,n973);
    nor g139(n519 ,n348 ,n346);
    nor g140(n386 ,n323 ,n50[11]);
    nor g141(n408 ,n328 ,n51[1]);
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2338), .Q(n50[9]));
    nand g143(n2328 ,n2019 ,n2242);
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1892), .Q(n42[4]));
    not g145(n971 ,n934);
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1850), .Q(n40[2]));
    nand g147(n1218 ,n7[26] ,n295);
    nand g148(n1427 ,n1211 ,n1037);
    nand g149(n2283 ,n1882 ,n2182);
    nand g150(n1988 ,n25[8] ,n1693);
    nand g151(n149 ,n52[1] ,n52[0]);
    not g152(n299 ,n305);
    nand g153(n2287 ,n53[15] ,n2259);
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n459), .Q(n43[2]));
    nand g155(n1989 ,n25[7] ,n1693);
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2205), .Q(n26[6]));
    nand g157(n1734 ,n827 ,n1321);
    nand g158(n2333 ,n1950 ,n2213);
    not g159(n968 ,n927);
    nand g160(n2088 ,n2495 ,n1701);
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1763), .Q(n30[2]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2321), .Q(n51[9]));
    not g163(n282 ,n281);
    nand g164(n1387 ,n838 ,n1020);
    nand g165(n104 ,n50[7] ,n103);
    nand g166(n1755 ,n1276 ,n1521);
    not g167(n1524 ,n1433);
    nand g168(n2067 ,n2478 ,n1696);
    nand g169(n628 ,n423 ,n493);
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2203), .Q(n26[8]));
    nand g171(n931 ,n11[28] ,n294);
    nand g172(n1299 ,n505 ,n988);
    not g173(n1550 ,n1481);
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n625), .Q(n39[2]));
    nor g175(n271 ,n34[5] ,n270);
    nor g176(n624 ,n2407 ,n561);
    nand g177(n1285 ,n6[23] ,n295);
    nand g178(n881 ,n16[13] ,n293);
    nand g179(n880 ,n657 ,n741);
    xnor g180(n2529 ,n34[3] ,n267);
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2229), .Q(n26[29]));
    nand g182(n1467 ,n40[29] ,n1139);
    nand g183(n1391 ,n1284 ,n1285);
    nand g184(n1338 ,n1087 ,n998);
    nand g185(n464 ,n52[6] ,n324);
    nor g186(n609 ,n577 ,n546);
    nand g187(n1281 ,n8[21] ,n299);
    nand g188(n2124 ,n26[29] ,n1695);
    nand g189(n871 ,n10[1] ,n293);
    nand g190(n702 ,n48[6] ,n527);
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n892), .Q(n48[2]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n619), .Q(n33[3]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n469), .Q(n43[1]));
    or g194(n1844 ,n1725 ,n1613);
    nand g195(n874 ,n659 ,n718);
    nand g196(n2132 ,n2470 ,n1698);
    nand g197(n1012 ,n17[0] ,n848);
    nand g198(n1013 ,n4[31] ,n297);
    nand g199(n950 ,n11[13] ,n664);
    nand g200(n2393 ,n1472 ,n2385);
    nand g201(n70 ,n46[6] ,n46[5]);
    nand g202(n2298 ,n53[4] ,n2259);
    nand g203(n121 ,n51[1] ,n51[0]);
    buf g204(n33[1], 1'b0);
    nand g205(n2198 ,n2031 ,n2147);
    nor g206(n364 ,n317 ,n50[0]);
    nand g207(n1479 ,n1221 ,n1065);
    nand g208(n2074 ,n2500 ,n1701);
    nor g209(n126 ,n117 ,n125);
    nor g210(n98 ,n89 ,n97);
    nand g211(n466 ,n50[12] ,n326);
    nand g212(n1451 ,n1163 ,n1024);
    or g213(n992 ,n580 ,n765);
    nand g214(n2052 ,n26[2] ,n1695);
    nand g215(n210 ,n46[5] ,n209);
    not g216(n314 ,n41[5]);
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2352), .Q(n53[13]));
    nand g218(n803 ,n10[2] ,n294);
    nand g219(n675 ,n2409 ,n592);
    nand g220(n1345 ,n40[6] ,n292);
    nor g221(n395 ,n326 ,n53[12]);
    nand g222(n151 ,n52[2] ,n150);
    nand g223(n1705 ,n1233 ,n1554);
    nand g224(n1817 ,n938 ,n1550);
    nand g225(n1442 ,n1097 ,n1251);
    or g226(n2173 ,n1442 ,n1948);
    nand g227(n1216 ,n7[27] ,n295);
    xnor g228(n2473 ,n52[3] ,n151);
    or g229(n365 ,n334 ,n41[0]);
    nand g230(n1490 ,n942 ,n1070);
    or g231(n1901 ,n1800 ,n1819);
    nand g232(n1063 ,n5[25] ,n297);
    nor g233(n391 ,n320 ,n50[15]);
    nor g234(n1160 ,n301 ,n958);
    not g235(n1150 ,n1102);
    not g236(n311 ,n38[0]);
    nand g237(n1681 ,n876 ,n1530);
    or g238(n1869 ,n1767 ,n1670);
    nand g239(n911 ,n643 ,n720);
    nand g240(n363 ,n41[0] ,n332);
    nand g241(n1140 ,n669 ,n853);
    nand g242(n678 ,n34[1] ,n524);
    not g243(n306 ,n1139);
    nand g244(n1432 ,n802 ,n1004);
    nand g245(n1169 ,n15[9] ,n300);
    not g246(n964 ,n922);
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n880), .Q(n49[5]));
    nand g248(n1610 ,n42[16] ,n289);
    buf g249(n33[0], 1'b0);
    nand g250(n191 ,n53[9] ,n189);
    nand g251(n1639 ,n40[3] ,n1397);
    dff g252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1585), .Q(n35[1]));
    nand g253(n1599 ,n40[21] ,n1397);
    xnor g254(n2455 ,n46[9] ,n215);
    nor g255(n1208 ,n2407 ,n970);
    nand g256(n2205 ,n2045 ,n2154);
    nand g257(n462 ,n50[5] ,n314);
    not g258(n1155 ,n1108);
    nand g259(n2188 ,n2009 ,n2137);
    nand g260(n230 ,n47[8] ,n229);
    not g261(n665 ,n666);
    nand g262(n1176 ,n8[5] ,n300);
    nor g263(n212 ,n46[7] ,n211);
    nand g264(n2223 ,n50[4] ,n1992);
    nor g265(n242 ,n48[7] ,n241);
    nand g266(n1672 ,n1212 ,n1522);
    xnor g267(n496 ,n41[3] ,n52[3]);
    nand g268(n653 ,n49[6] ,n588);
    nand g269(n2234 ,n51[12] ,n1991);
    dff g270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n906), .Q(n46[5]));
    not g271(n2155 ,n2046);
    nand g272(n2360 ,n1940 ,n2297);
    xnor g273(n779 ,n523 ,n34[0]);
    nand g274(n780 ,n37[3] ,n665);
    or g275(n1866 ,n1759 ,n1666);
    nand g276(n2103 ,n12[14] ,n1694);
    nand g277(n637 ,n331 ,n573);
    nand g278(n2352 ,n1996 ,n2289);
    nand g279(n2241 ,n51[5] ,n1991);
    nand g280(n461 ,n38[0] ,n3[1]);
    nand g281(n751 ,n34[12] ,n524);
    or g282(n1890 ,n1790 ,n1712);
    dff g283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2347), .Q(n53[0]));
    not g284(n185 ,n184);
    nand g285(n218 ,n47[1] ,n47[0]);
    nand g286(n111 ,n50[11] ,n110);
    nor g287(n1695 ,n671 ,n1397);
    nor g288(n120 ,n51[1] ,n51[0]);
    nor g289(n1194 ,n2407 ,n962);
    nand g290(n1233 ,n9[19] ,n849);
    nand g291(n954 ,n10[14] ,n293);
    nand g292(n2345 ,n1962 ,n2224);
    nand g293(n1446 ,n42[8] ,n1139);
    nand g294(n1611 ,n40[16] ,n291);
    nand g295(n1962 ,n2503 ,n1700);
    nand g296(n643 ,n49[3] ,n588);
    nand g297(n2184 ,n2001 ,n2133);
    nand g298(n2299 ,n53[3] ,n2259);
    dff g299(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2358), .Q(n53[8]));
    nand g300(n440 ,n38[3] ,n331);
    nand g301(n2197 ,n2029 ,n2146);
    not g302(n2154 ,n2044);
    xnor g303(n2443 ,n47[6] ,n225);
    nand g304(n240 ,n48[5] ,n239);
    dff g305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2248), .Q(n25[29]));
    dff g306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1359), .Q(n31[4]));
    xnor g307(n2526 ,n34[6] ,n272);
    nand g308(n2399 ,n20[1] ,n2397);
    not g309(n1548 ,n1473);
    not g310(n1411 ,n1341);
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n792), .Q(n49[0]));
    nand g312(n1138 ,n8[25] ,n300);
    nor g313(n1320 ,n579 ,n980);
    nor g314(n2453 ,n212 ,n214);
    nand g315(n2387 ,n45[2] ,n2383);
    nand g316(n2268 ,n1989 ,n2110);
    or g317(n1861 ,n1752 ,n1661);
    not g318(n1151 ,n1104);
    nor g319(n1577 ,n1298 ,n1297);
    not g320(n1834 ,n1773);
    dff g321(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2198), .Q(n26[13]));
    nand g322(n1243 ,n6[8] ,n296);
    nand g323(n566 ,n449 ,n402);
    dff g324(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2328), .Q(n51[4]));
    nand g325(n1585 ,n303 ,n1328);
    nor g326(n1352 ,n2407 ,n1150);
    nand g327(n223 ,n47[4] ,n222);
    nand g328(n923 ,n753 ,n679);
    not g329(n1410 ,n1340);
    nand g330(n485 ,n44[0] ,n44[1]);
    dff g331(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1870), .Q(n42[9]));
    nor g332(n1207 ,n2407 ,n969);
    nor g333(n616 ,n2407 ,n517);
    nand g334(n1213 ,n9[28] ,n299);
    dff g335(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2366), .Q(n52[14]));
    dff g336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n846), .Q(n47[0]));
    dff g337(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1194), .Q(n34[14]));
    xnor g338(n2477 ,n52[7] ,n158);
    nor g339(n2464 ,n190 ,n192);
    nand g340(n1726 ,n1088 ,n1339);
    dff g341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2174), .Q(n40[29]));
    not g342(n266 ,n265);
    xnor g343(n510 ,n41[10] ,n52[10]);
    nand g344(n2318 ,n2075 ,n2232);
    nand g345(n1716 ,n42[29] ,n289);
    nand g346(n1388 ,n37[2] ,n1141);
    not g347(n1526 ,n1435);
    not g348(n199 ,n198);
    nand g349(n1814 ,n1231 ,n1553);
    not g350(n1699 ,n1700);
    not g351(n1541 ,n1459);
    nor g352(n403 ,n328 ,n52[1]);
    dff g353(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2272), .Q(n25[11]));
    dff g354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2199), .Q(n26[12]));
    nand g355(n1650 ,n1109 ,n1415);
    nand g356(n2005 ,n26[25] ,n1695);
    nand g357(n2321 ,n2079 ,n2237);
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2253), .Q(n25[22]));
    nand g359(n1236 ,n7[18] ,n847);
    nand g360(n1437 ,n42[7] ,n1139);
    nand g361(n1110 ,n7[3] ,n295);
    nand g362(n1671 ,n1243 ,n1529);
    nand g363(n443 ,n50[7] ,n327);
    dff g364(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2191), .Q(n26[20]));
    nor g365(n613 ,n557 ,n489);
    nand g366(n1316 ,n41[0] ,n1139);
    nand g367(n724 ,n48[7] ,n527);
    nor g368(n241 ,n232 ,n240);
    not g369(n2395 ,n18[1]);
    nor g370(n285 ,n34[13] ,n284);
    nand g371(n1821 ,n925 ,n1546);
    nor g372(n197 ,n53[13] ,n196);
    nand g373(n1219 ,n9[25] ,n299);
    nand g374(n1128 ,n8[30] ,n299);
    nand g375(n2340 ,n1957 ,n2220);
    nand g376(n1370 ,n44[0] ,n292);
    nand g377(n78 ,n47[7] ,n77);
    nand g378(n1264 ,n6[13] ,n296);
    nor g379(n77 ,n76 ,n74);
    nand g380(n1003 ,n5[6] ,n297);
    dff g381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2317), .Q(n51[15]));
    nand g382(n1097 ,n8[3] ,n299);
    not g383(n1405 ,n1331);
    nand g384(n2384 ,n1291 ,n2382);
    nand g385(n1822 ,n1197 ,n1545);
    or g386(n593 ,n311 ,n484);
    not g387(n319 ,n41[8]);
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2206), .Q(n26[5]));
    dff g389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2190), .Q(n26[21]));
    dff g390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2355), .Q(n53[10]));
    nand g391(n1330 ,n40[13] ,n292);
    not g392(n324 ,n41[6]);
    nor g393(n378 ,n313 ,n51[9]);
    nand g394(n283 ,n34[11] ,n282);
    nand g395(n1448 ,n1258 ,n1038);
    nor g396(n518 ,n350 ,n352);
    nand g397(n1029 ,n4[18] ,n298);
    nand g398(n1053 ,n13[2] ,n297);
    nand g399(n2339 ,n1956 ,n2219);
    nand g400(n982 ,n507 ,n773);
    nand g401(n1806 ,n1230 ,n1486);
    nand g402(n1112 ,n823 ,n789);
    nand g403(n843 ,n10[19] ,n293);
    nor g404(n161 ,n146 ,n160);
    xnor g405(n2496 ,n51[11] ,n137);
    not g406(n150 ,n149);
    not g407(n2152 ,n2040);
    dff g408(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2342), .Q(n50[5]));
    nand g409(n712 ,n2444 ,n526);
    nor g410(n667 ,n410 ,n539);
    dff g411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1866), .Q(n42[16]));
    nand g412(n245 ,n48[8] ,n244);
    nor g413(n227 ,n47[7] ,n226);
    nand g414(n62 ,n22[0] ,n61);
    nand g415(n1931 ,n1267 ,n1832);
    nand g416(n2025 ,n26[16] ,n1695);
    not g417(n1144 ,n1143);
    dff g418(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2329), .Q(n51[3]));
    nand g419(n1269 ,n8[15] ,n299);
    nand g420(n1600 ,n42[21] ,n289);
    not g421(n1558 ,n1499);
    dff g422(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2276), .Q(n25[15]));
    nand g423(n1256 ,n8[7] ,n299);
    or g424(n1867 ,n1760 ,n1667);
    nand g425(n2296 ,n53[6] ,n2259);
    nand g426(n1597 ,n42[22] ,n289);
    not g427(n294 ,n302);
    dff g428(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2208), .Q(n26[3]));
    nand g429(n1655 ,n833 ,n1420);
    nand g430(n1089 ,n9[8] ,n299);
    nand g431(n753 ,n34[9] ,n524);
    or g432(n1848 ,n1730 ,n1647);
    nand g433(n429 ,n50[11] ,n323);
    nand g434(n837 ,n10[25] ,n294);
    nand g435(n2006 ,n1593 ,n1592);
    xnor g436(n2424 ,n49[5] ,n253);
    nand g437(n1087 ,n9[9] ,n299);
    nand g438(n1279 ,n8[20] ,n849);
    nor g439(n1350 ,n2407 ,n1149);
    not g440(n969 ,n928);
    nand g441(n290 ,n671 ,n1146);
    nor g442(n854 ,n540 ,n671);
    xor g443(n2429 ,n48[1] ,n48[0]);
    nand g444(n1099 ,n811 ,n780);
    nand g445(n1511 ,n954 ,n1266);
    nor g446(n1360 ,n2407 ,n1155);
    nand g447(n2049 ,n26[4] ,n1695);
    nand g448(n1271 ,n8[16] ,n849);
    nand g449(n740 ,n2455 ,n528);
    nand g450(n757 ,n312 ,n610);
    nand g451(n181 ,n53[3] ,n180);
    nor g452(n257 ,n49[7] ,n256);
    nand g453(n804 ,n11[9] ,n293);
    nand g454(n1636 ,n40[5] ,n1397);
    nand g455(n785 ,n36[2] ,n665);
    nor g456(n517 ,n351 ,n355);
    nand g457(n2323 ,n2088 ,n2236);
    nand g458(n1094 ,n9[6] ,n300);
    nand g459(n1604 ,n42[19] ,n289);
    nand g460(n952 ,n10[12] ,n293);
    not g461(n338 ,n49[0]);
    nand g462(n906 ,n690 ,n735);
    or g463(n1892 ,n1776 ,n1677);
    nand g464(n1070 ,n5[19] ,n297);
    nand g465(n862 ,n10[11] ,n664);
    nand g466(n693 ,n2427 ,n525);
    nand g467(n1129 ,n6[30] ,n296);
    nand g468(n132 ,n51[7] ,n131);
    dff g469(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2319), .Q(n51[13]));
    nor g470(n2533 ,n75 ,n78);
    not g471(n1157 ,n1112);
    nand g472(n630 ,n455 ,n496);
    nor g473(n2259 ,n612 ,n1840);
    nand g474(n71 ,n46[9] ,n46[8]);
    nand g475(n904 ,n692 ,n695);
    nand g476(n1476 ,n936 ,n1220);
    nand g477(n1179 ,n14[5] ,n296);
    nand g478(n791 ,n2408 ,n676);
    nand g479(n1231 ,n9[20] ,n300);
    nand g480(n1481 ,n1224 ,n1066);
    nand g481(n265 ,n34[1] ,n34[0]);
    nand g482(n1664 ,n844 ,n1566);
    dff g483(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1935), .Q(n35[3]));
    nand g484(n2307 ,n52[10] ,n2260);
    nor g485(n525 ,n2535 ,n486);
    nand g486(n2120 ,n26[31] ,n1695);
    nand g487(n1485 ,n1229 ,n1068);
    or g488(n1904 ,n1805 ,n1816);
    dff g489(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1871), .Q(n42[8]));
    nand g490(n834 ,n10[28] ,n664);
    nand g491(n2058 ,n26[0] ,n1695);
    nand g492(n912 ,n10[3] ,n664);
    or g493(n351 ,n35[1] ,n35[2]);
    nand g494(n2114 ,n12[3] ,n1694);
    nor g495(n405 ,n320 ,n53[15]);
    nand g496(n1226 ,n9[22] ,n849);
    or g497(n989 ,n556 ,n770);
    dff g498(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n806), .Q(n46[8]));
    dff g499(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2343), .Q(n50[1]));
    not g500(n325 ,n41[2]);
    or g501(n1900 ,n1799 ,n1820);
    nand g502(n1121 ,n19[0] ,n295);
    xnor g503(n2472 ,n52[2] ,n149);
    xnor g504(n2458 ,n53[3] ,n179);
    nor g505(n1198 ,n2407 ,n960);
    nand g506(n615 ,n43[0] ,n537);
    nand g507(n2398 ,n20[0] ,n2397);
    nor g508(n377 ,n318 ,n52[14]);
    nand g509(n872 ,n10[23] ,n293);
    nand g510(n457 ,n53[12] ,n326);
    nand g511(n1803 ,n937 ,n1480);
    dff g512(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2265), .Q(n25[4]));
    nand g513(n1376 ,n42[30] ,n1139);
    nand g514(n553 ,n432 ,n392);
    nand g515(n1212 ,n6[10] ,n847);
    or g516(n468 ,n324 ,n51[6]);
    dff g517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1868), .Q(n42[13]));
    nand g518(n186 ,n53[6] ,n185);
    nand g519(n2372 ,n2067 ,n2309);
    nor g520(n586 ,n2[0] ,n356);
    xnor g521(n508 ,n41[1] ,n53[1]);
    nand g522(n918 ,n16[1] ,n664);
    nand g523(n1996 ,n2468 ,n1698);
    not g524(n209 ,n208);
    not g525(n676 ,n675);
    nand g526(n1280 ,n6[21] ,n847);
    dff g527(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2362), .Q(n53[3]));
    nand g528(n705 ,n2437 ,n530);
    nand g529(n1145 ,n672 ,n775);
    nand g530(n1973 ,n25[23] ,n1693);
    not g531(n1421 ,n1379);
    nand g532(n465 ,n50[9] ,n313);
    not g533(n342 ,n45[0]);
    nand g534(n1728 ,n1342 ,n1001);
    dff g535(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n411), .Q(n33[7]));
    nand g536(n1772 ,n1254 ,n1431);
    nand g537(n1512 ,n42[14] ,n1139);
    nor g538(n1363 ,n2407 ,n1157);
    nor g539(n389 ,n316 ,n52[4]);
    nand g540(n2102 ,n12[15] ,n1694);
    nand g541(n648 ,n2530 ,n523);
    not g542(n1423 ,n1383);
    dff g543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1878), .Q(n42[2]));
    or g544(n1896 ,n1794 ,n1824);
    or g545(n2172 ,n1367 ,n1921);
    nand g546(n1292 ,n1277 ,n1028);
    nand g547(n1259 ,n6[9] ,n847);
    not g548(n960 ,n917);
    not g549(n194 ,n193);
    nand g550(n1660 ,n1287 ,n1425);
    nand g551(n81 ,n48[9] ,n48[8]);
    dff g552(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1586), .Q(n37[0]));
    not g553(n252 ,n251);
    or g554(n1891 ,n1789 ,n1690);
    nand g555(n701 ,n2433 ,n530);
    nand g556(n1445 ,n42[1] ,n1139);
    not g557(n2159 ,n2055);
    nand g558(n1997 ,n1219 ,n1838);
    nand g559(n1920 ,n1091 ,n1826);
    nand g560(n2073 ,n2472 ,n1696);
    nand g561(n897 ,n16[9] ,n293);
    nand g562(n763 ,n492 ,n609);
    dff g563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1861), .Q(n42[21]));
    xnor g564(n2522 ,n34[10] ,n279);
    nand g565(n1938 ,n2462 ,n1698);
    not g566(n178 ,n177);
    xnor g567(n2528 ,n34[4] ,n269);
    nand g568(n2063 ,n2482 ,n1696);
    nor g569(n501 ,n390 ,n406);
    nand g570(n1079 ,n7[12] ,n296);
    nand g571(n1465 ,n1202 ,n1058);
    or g572(n774 ,n396 ,n629);
    or g573(n1888 ,n1787 ,n1688);
    not g574(n2145 ,n2026);
    nand g575(n1225 ,n7[23] ,n847);
    nor g576(n1348 ,n2407 ,n1147);
    nand g577(n2233 ,n51[13] ,n1991);
    nand g578(n1185 ,n14[3] ,n295);
    nand g579(n1800 ,n1216 ,n1474);
    nand g580(n1647 ,n1095 ,n1413);
    nand g581(n632 ,n420 ,n504);
    nand g582(n698 ,n46[9] ,n529);
    nand g583(n1021 ,n13[5] ,n848);
    not g584(n337 ,n44[0]);
    nand g585(n2327 ,n2021 ,n2241);
    nand g586(n1930 ,n1569 ,n1758);
    not g587(n481 ,n480);
    nand g588(n1753 ,n1278 ,n1300);
    or g589(n345 ,n39[0] ,n39[1]);
    nand g590(n1173 ,n15[7] ,n299);
    nand g591(n1381 ,n1134 ,n1017);
    not g592(n1565 ,n1518);
    nand g593(n1596 ,n42[23] ,n289);
    nand g594(n288 ,n34[14] ,n287);
    nand g595(n1294 ,n993 ,n994);
    nand g596(n818 ,n31[5] ,n666);
    nand g597(n891 ,n726 ,n745);
    dff g598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2372), .Q(n52[8]));
    nand g599(n2292 ,n53[10] ,n2259);
    or g600(n2411 ,n65 ,n68);
    dff g601(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n900), .Q(n49[8]));
    dff g602(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2332), .Q(n50[15]));
    xnor g603(n490 ,n41[5] ,n51[5]);
    nand g604(n416 ,n53[14] ,n318);
    not g605(n1545 ,n1463);
    nand g606(n1307 ,n41[9] ,n292);
    dff g607(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2170), .Q(n42[12]));
    nor g608(n412 ,n43[1] ,n43[2]);
    not g609(n89 ,n50[4]);
    nand g610(n765 ,n522 ,n613);
    nand g611(n688 ,n2449 ,n528);
    nand g612(n1668 ,n1265 ,n1562);
    xnor g613(n2524 ,n34[8] ,n276);
    nand g614(n2379 ,n1943 ,n2300);
    dff g615(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n904), .Q(n46[7]));
    nand g616(n1515 ,n42[16] ,n292);
    nand g617(n679 ,n2523 ,n523);
    or g618(n370 ,n316 ,n53[4]);
    not g619(n690 ,n529);
    nand g620(n1923 ,n831 ,n1829);
    nand g621(n1278 ,n6[20] ,n295);
    not g622(n101 ,n100);
    dff g623(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1898), .Q(n40[31]));
    dff g624(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n31[6]));
    xnor g625(n2451 ,n46[5] ,n208);
    dff g626(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1859), .Q(n42[25]));
    nand g627(n2047 ,n26[5] ,n1695);
    nand g628(n1369 ,n829 ,n1011);
    not g629(n320 ,n41[15]);
    nand g630(n888 ,n706 ,n701);
    nand g631(n272 ,n34[5] ,n270);
    dff g632(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2325), .Q(n51[7]));
    nand g633(n1001 ,n5[7] ,n298);
    nand g634(n1482 ,n40[23] ,n1139);
    dff g635(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n890), .Q(n48[4]));
    nand g636(n1928 ,n1571 ,n1751);
    nand g637(n2231 ,n51[15] ,n1991);
    nand g638(n2247 ,n1966 ,n2086);
    nand g639(n1043 ,n4[1] ,n297);
    dff g640(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2283), .Q(n50[0]));
    nor g641(n671 ,n44[1] ,n533);
    not g642(n645 ,n587);
    nand g643(n1131 ,n6[29] ,n295);
    nand g644(n2109 ,n12[8] ,n1694);
    nand g645(n444 ,n50[4] ,n316);
    not g646(n1149 ,n1101);
    not g647(n2162 ,n2121);
    or g648(n1855 ,n1740 ,n1655);
    nand g649(n1047 ,n13[9] ,n848);
    nand g650(n972 ,n608 ,n304);
    nand g651(n1076 ,n5[13] ,n848);
    nand g652(n1787 ,n1172 ,n1308);
    nand g653(n1251 ,n6[3] ,n296);
    nand g654(n439 ,n53[4] ,n316);
    or g655(n1842 ,n1722 ,n1709);
    nand g656(n942 ,n11[19] ,n294);
    nand g657(n1253 ,n8[6] ,n300);
    nand g658(n1805 ,n1227 ,n1483);
    nand g659(n1977 ,n25[19] ,n1693);
    nand g660(n1339 ,n40[9] ,n292);
    nor g661(n562 ,n39[0] ,n473);
    nand g662(n1215 ,n9[27] ,n849);
    nand g663(n1784 ,n1166 ,n1305);
    nand g664(n2014 ,n1603 ,n1602);
    nand g665(n2182 ,n50[0] ,n1992);
    not g666(n152 ,n151);
    dff g667(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2379), .Q(n53[2]));
    nand g668(n417 ,n52[2] ,n325);
    nand g669(n728 ,n2446 ,n526);
    nand g670(n1393 ,n1282 ,n1283);
    nand g671(n694 ,n46[8] ,n529);
    nand g672(n941 ,n11[20] ,n293);
    nand g673(n1139 ,n531 ,n791);
    or g674(n601 ,n2409 ,n532);
    not g675(n323 ,n41[11]);
    nand g676(n2002 ,n26[26] ,n1695);
    nand g677(n1918 ,n1567 ,n1577);
    nor g678(n1228 ,n2407 ,n971);
    dff g679(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1894), .Q(n41[3]));
    dff g680(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n883), .Q(n48[9]));
    nand g681(n1168 ,n14[10] ,n295);
    xnor g682(n2515 ,n50[15] ,n116);
    dff g683(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2334), .Q(n50[13]));
    nand g684(n1764 ,n29[3] ,n1399);
    or g685(n1849 ,n1731 ,n1649);
    nand g686(n1799 ,n1214 ,n1471);
    nand g687(n2189 ,n2011 ,n2138);
    nand g688(n916 ,n16[2] ,n664);
    not g689(n1837 ,n1801);
    not g690(n2383 ,n2384);
    nand g691(n1721 ,n40[27] ,n1397);
    nand g692(n1036 ,n4[11] ,n297);
    dff g693(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2255), .Q(n25[23]));
    nand g694(n2086 ,n12[30] ,n1694);
    dff g695(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1907), .Q(n40[19]));
    nand g696(n188 ,n53[7] ,n187);
    not g697(n959 ,n913);
    nor g698(n380 ,n325 ,n50[2]);
    nand g699(n2332 ,n1949 ,n2212);
    nor g700(n2486 ,n122 ,n120);
    nor g701(n847 ,n591 ,n601);
    dff g702(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1364), .Q(n31[0]));
    nand g703(n1240 ,n7[16] ,n295);
    nand g704(n1458 ,n1180 ,n1051);
    nand g705(n2285 ,n52[0] ,n2260);
    nand g706(n2095 ,n12[22] ,n1694);
    nand g707(n2127 ,n25[0] ,n1693);
    or g708(n500 ,n403 ,n381);
    nand g709(n1810 ,n1493 ,n1072);
    nand g710(n661 ,n2526 ,n523);
    nor g711(n105 ,n90 ,n104);
    nand g712(n2019 ,n2489 ,n1701);
    nand g713(n1692 ,n42[10] ,n289);
    nand g714(n1178 ,n15[13] ,n299);
    dff g715(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2177), .Q(n40[17]));
    nand g716(n1005 ,n5[5] ,n297);
    or g717(n1871 ,n1771 ,n1671);
    nand g718(n2060 ,n2485 ,n1696);
    or g719(n2281 ,n2178 ,n1881);
    xnor g720(n2506 ,n50[6] ,n100);
    dff g721(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2192), .Q(n26[19]));
    nand g722(n2348 ,n1914 ,n2285);
    nand g723(n775 ,n514 ,n626);
    nand g724(n2098 ,n12[19] ,n1694);
    nand g725(n1347 ,n40[5] ,n292);
    nand g726(n2330 ,n2083 ,n2244);
    nand g727(n778 ,n639 ,n302);
    nand g728(n1517 ,n42[17] ,n1139);
    nand g729(n1102 ,n815 ,n783);
    or g730(n1876 ,n1774 ,n1672);
    dff g731(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2258), .Q(n26[1]));
    not g732(n173 ,n53[4]);
    not g733(n340 ,n46[0]);
    not g734(n64 ,n24[1]);
    xnor g735(n2474 ,n52[4] ,n153);
    nand g736(n1031 ,n4[16] ,n848);
    nand g737(n1431 ,n42[0] ,n292);
    nand g738(n424 ,n51[12] ,n326);
    nand g739(n622 ,n38[1] ,n532);
    nand g740(n2338 ,n1955 ,n2218);
    not g741(n1527 ,n1439);
    dff g742(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1124), .Q(n34[0]));
    nand g743(n936 ,n11[25] ,n294);
    nand g744(n1038 ,n13[15] ,n297);
    dff g745(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n869), .Q(n47[5]));
    nand g746(n1091 ,n9[7] ,n849);
    nand g747(n915 ,n16[3] ,n664);
    not g748(n1833 ,n1766);
    or g749(n1911 ,n1813 ,n1708);
    nor g750(n347 ,n38[0] ,n3[2]);
    nand g751(n1925 ,n872 ,n1830);
    nand g752(n939 ,n11[22] ,n664);
    nand g753(n1823 ,n1193 ,n1544);
    not g754(n303 ,n847);
    nand g755(n1118 ,n7[1] ,n847);
    nand g756(n1186 ,n15[2] ,n849);
    not g757(n280 ,n279);
    nand g758(n1622 ,n40[11] ,n1397);
    dff g759(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n972), .Q(n38[0]));
    nor g760(n2471 ,n150 ,n148);
    not g761(n309 ,n2533);
    nand g762(n1840 ,n308 ,n1697);
    dff g763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2360), .Q(n53[5]));
    nand g764(n1235 ,n9[18] ,n849);
    nand g765(n1673 ,n1259 ,n1524);
    dff g766(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n793), .Q(n48[0]));
    not g767(n1525 ,n1434);
    nand g768(n420 ,n51[14] ,n318);
    dff g769(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2368), .Q(n52[12]));
    dff g770(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1896), .Q(n41[1]));
    nor g771(n561 ,n39[1] ,n481);
    nand g772(n2309 ,n52[8] ,n2260);
    nand g773(n193 ,n53[10] ,n192);
    nand g774(n1037 ,n4[10] ,n297);
    nand g775(n1244 ,n7[15] ,n295);
    nand g776(n1593 ,n40[24] ,n1397);
    nand g777(n824 ,n11[2] ,n664);
    or g778(n1853 ,n1735 ,n1652);
    nand g779(n1615 ,n42[14] ,n289);
    nand g780(n1946 ,n2465 ,n1698);
    nor g781(n984 ,n512 ,n767);
    xor g782(n2420 ,n49[1] ,n49[0]);
    not g783(n1839 ,n1810);
    nand g784(n1135 ,n6[27] ,n296);
    dff g785(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2194), .Q(n26[17]));
    nand g786(n1961 ,n2504 ,n1700);
    nand g787(n1947 ,n1176 ,n1834);
    or g788(n1575 ,n992 ,n1295);
    buf g789(n33[2], 1'b0);
    dff g790(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2200), .Q(n26[11]));
    nand g791(n1669 ,n305 ,n1504);
    nand g792(n2359 ,n1939 ,n2296);
    nand g793(n716 ,n34[4] ,n524);
    xnor g794(n2500 ,n51[15] ,n144);
    nand g795(n1460 ,n916 ,n1053);
    not g796(n312 ,n43[0]);
    nand g797(n1239 ,n9[16] ,n299);
    nand g798(n1745 ,n1288 ,n1386);
    or g799(n2179 ,n1343 ,n1920);
    dff g800(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1928), .Q(n36[2]));
    dff g801(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2246), .Q(n25[31]));
    nand g802(n225 ,n47[5] ,n224);
    nand g803(n636 ,n2520 ,n523);
    nand g804(n1758 ,n36[0] ,n1400);
    nand g805(n995 ,n5[12] ,n848);
    nand g806(n1719 ,n1246 ,n1558);
    xor g807(n2447 ,n46[1] ,n46[0]);
    nand g808(n360 ,n53[0] ,n317);
    nand g809(n2125 ,n26[28] ,n1695);
    nand g810(n67 ,n24[0] ,n66);
    xnor g811(n2504 ,n50[4] ,n97);
    or g812(n585 ,n331 ,n347);
    nand g813(n2056 ,n26[1] ,n1695);
    nor g814(n600 ,n502 ,n543);
    dff g815(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2249), .Q(n25[28]));
    dff g816(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1847), .Q(n40[6]));
    nand g817(n1469 ,n42[10] ,n1139);
    not g818(n957 ,n864);
    nand g819(n1252 ,n8[9] ,n300);
    nand g820(n438 ,n53[2] ,n325);
    nand g821(n2122 ,n26[30] ,n1695);
    nor g822(n168 ,n147 ,n167);
    nand g823(n2000 ,n1721 ,n1720);
    nand g824(n793 ,n727 ,n606);
    or g825(n497 ,n380 ,n391);
    nor g826(n2422 ,n250 ,n252);
    nand g827(n1234 ,n7[19] ,n847);
    or g828(n401 ,n320 ,n52[15]);
    nand g829(n1074 ,n5[15] ,n297);
    nand g830(n1634 ,n40[6] ,n1397);
    not g831(n1828 ,n1736);
    nand g832(n692 ,n46[7] ,n529);
    nand g833(n1499 ,n948 ,n1002);
    nand g834(n1372 ,n42[31] ,n1139);
    nand g835(n1922 ,n828 ,n1828);
    nand g836(n772 ,n38[0] ,n667);
    or g837(n400 ,n316 ,n50[4]);
    nand g838(n1224 ,n9[23] ,n300);
    not g839(n2401 ,n2419);
    nand g840(n687 ,n2435 ,n530);
    nand g841(n2082 ,n2488 ,n1701);
    nand g842(n243 ,n48[7] ,n241);
    nand g843(n890 ,n749 ,n704);
    dff g844(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1192), .Q(n34[15]));
    dff g845(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n885), .Q(n48[8]));
    dff g846(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n878), .Q(n49[9]));
    nand g847(n1177 ,n15[5] ,n299);
    nand g848(n2083 ,n2487 ,n1701);
    nor g849(n211 ,n202 ,n210);
    nand g850(n768 ,n499 ,n596);
    dff g851(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n840), .Q(n49[2]));
    dff g852(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1842), .Q(n40[13]));
    nand g853(n938 ,n11[23] ,n293);
    nor g854(n2444 ,n227 ,n229);
    xor g855(n520 ,n41[11] ,n53[11]);
    nand g856(n896 ,n649 ,n730);
    dff g857(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1200), .Q(n34[9]));
    nor g858(n357 ,n311 ,n3[3]);
    nor g859(n1196 ,n2407 ,n964);
    nand g860(n1939 ,n2461 ,n1698);
    nand g861(n1203 ,n8[1] ,n299);
    nand g862(n2306 ,n52[11] ,n2260);
    nor g863(n87 ,n86 ,n84);
    nand g864(n1595 ,n799 ,n1405);
    nand g865(n2341 ,n1959 ,n2221);
    nand g866(n2030 ,n1617 ,n1618);
    nand g867(n2343 ,n1964 ,n2226);
    or g868(n1903 ,n1804 ,n1817);
    nand g869(n1385 ,n1138 ,n1019);
    nand g870(n1975 ,n25[21] ,n1693);
    nand g871(n821 ,n31[3] ,n666);
    nand g872(n2326 ,n2081 ,n2240);
    not g873(n174 ,n53[8]);
    or g874(n760 ,n372 ,n630);
    nand g875(n2403 ,n22[0] ,n2402);
    nand g876(n200 ,n53[14] ,n199);
    dff g877(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2251), .Q(n25[26]));
    not g878(n304 ,n848);
    or g879(n1886 ,n1785 ,n1686);
    nand g880(n1985 ,n25[11] ,n1693);
    nand g881(n1358 ,n40[3] ,n292);
    nand g882(n738 ,n46[0] ,n529);
    nor g883(n68 ,n2412 ,n67);
    nand g884(n1237 ,n9[17] ,n849);
    or g885(n589 ,n311 ,n414);
    nand g886(n2282 ,n1579 ,n2181);
    nand g887(n948 ,n11[14] ,n293);
    dff g888(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n895), .Q(n47[7]));
    nand g889(n480 ,n35[1] ,n2533);
    or g890(n1872 ,n1775 ,n1675);
    nand g891(n2018 ,n26[18] ,n1695);
    nand g892(n425 ,n51[11] ,n323);
    nand g893(n1303 ,n41[13] ,n292);
    dff g894(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1879), .Q(n41[15]));
    xor g895(n2438 ,n47[1] ,n47[0]);
    xnor g896(n2461 ,n53[6] ,n184);
    nand g897(n1190 ,n15[1] ,n299);
    dff g898(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2370), .Q(n52[9]));
    nand g899(n723 ,n48[9] ,n527);
    nand g900(n1018 ,n4[26] ,n298);
    nor g901(n1124 ,n2407 ,n779);
    nand g902(n943 ,n11[18] ,n664);
    nand g903(n2265 ,n2131 ,n2113);
    nand g904(n944 ,n11[17] ,n664);
    nand g905(n502 ,n362 ,n404);
    nand g906(n1477 ,n935 ,n1218);
    dff g907(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2269), .Q(n25[8]));
    dff g908(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2331), .Q(n51[1]));
    dff g909(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2210), .Q(n25[19]));
    nand g910(n1791 ,n1181 ,n1312);
    nand g911(n2370 ,n2066 ,n2308);
    nand g912(n1598 ,n40[22] ,n291);
    nor g913(n388 ,n324 ,n53[6]);
    nand g914(n1042 ,n4[8] ,n297);
    nand g915(n2187 ,n2007 ,n2136);
    not g916(n2141 ,n2016);
    nor g917(n176 ,n53[1] ,n53[0]);
    nand g918(n1776 ,n1184 ,n1440);
    nand g919(n905 ,n696 ,n691);
    nand g920(n907 ,n16[7] ,n294);
    nand g921(n754 ,n34[6] ,n524);
    nand g922(n486 ,n35[3] ,n308);
    nand g923(n1713 ,n42[30] ,n289);
    nand g924(n2080 ,n2492 ,n1701);
    nand g925(n1663 ,n843 ,n1404);
    xnor g926(n2448 ,n46[2] ,n203);
    nand g927(n631 ,n451 ,n491);
    nand g928(n2337 ,n1954 ,n2217);
    dff g929(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2351), .Q(n53[14]));
    nand g930(n2017 ,n26[19] ,n1695);
    buf g931(n32[5], 1'b0);
    nand g932(n634 ,n2518 ,n523);
    nor g933(n472 ,n329 ,n43[2]);
    nor g934(n1364 ,n2407 ,n1158);
    xor g935(n513 ,n41[3] ,n50[3]);
    not g936(n2158 ,n2053);
    nand g937(n828 ,n23[0] ,n293);
    or g938(n348 ,n37[0] ,n37[1]);
    dff g939(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n623), .Q(n39[0]));
    dff g940(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n901), .Q(n47[1]));
    nand g941(n1500 ,n909 ,n1050);
    nor g942(n852 ,n301 ,n620);
    or g943(n346 ,n37[2] ,n37[3]);
    nand g944(n1678 ,n1241 ,n1408);
    nand g945(n1257 ,n8[8] ,n849);
    nand g946(n928 ,n755 ,n648);
    not g947(n327 ,n41[7]);
    nand g948(n2335 ,n1953 ,n2216);
    nand g949(n1801 ,n1475 ,n1062);
    not g950(n117 ,n51[4]);
    nand g951(n1792 ,n1185 ,n1313);
    dff g952(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2267), .Q(n25[6]));
    nand g953(n1614 ,n42[15] ,n289);
    nand g954(n484 ,n44[0] ,n312);
    not g955(n1564 ,n1516);
    not g956(n958 ,n873);
    nand g957(n899 ,n652 ,n733);
    nand g958(n1438 ,n830 ,n1249);
    nand g959(n1220 ,n7[25] ,n296);
    nand g960(n1440 ,n42[4] ,n1139);
    nor g961(n196 ,n175 ,n195);
    nand g962(n1809 ,n1236 ,n1492);
    nand g963(n1452 ,n1165 ,n1023);
    nand g964(n2350 ,n2132 ,n2287);
    nand g965(n1586 ,n850 ,n1323);
    nand g966(n767 ,n510 ,n595);
    nand g967(n1766 ,n1507 ,n1035);
    nand g968(n2400 ,n2418 ,n2409);
    nand g969(n730 ,n2443 ,n526);
    nor g970(n488 ,n472 ,n353);
    nand g971(n1284 ,n8[23] ,n299);
    nand g972(n2111 ,n12[6] ,n1694);
    not g973(n1156 ,n1111);
    nand g974(n649 ,n47[6] ,n587);
    nand g975(n2386 ,n45[0] ,n2383);
    nand g976(n1631 ,n42[7] ,n289);
    nand g977(n1948 ,n912 ,n1835);
    not g978(n1552 ,n1485);
    nand g979(n1497 ,n1242 ,n1074);
    not g980(n91 ,n50[12]);
    nor g981(n1401 ,n574 ,n975);
    nand g982(n1964 ,n2501 ,n1700);
    not g983(n147 ,n52[12]);
    nand g984(n547 ,n442 ,n374);
    not g985(n122 ,n121);
    or g986(n1860 ,n1747 ,n1660);
    nand g987(n233 ,n48[1] ,n48[0]);
    xnor g988(n2465 ,n53[10] ,n191);
    dff g989(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2193), .Q(n26[18]));
    dff g990(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2326), .Q(n51[6]));
    dff g991(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2318), .Q(n51[14]));
    not g992(n341 ,n48[0]);
    not g993(n657 ,n588);
    nand g994(n680 ,n2522 ,n523);
    nand g995(n1379 ,n834 ,n1016);
    nand g996(n842 ,n10[20] ,n293);
    nand g997(n1782 ,n1162 ,n1303);
    dff g998(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2167), .Q(n42[23]));
    nand g999(n1126 ,n6[31] ,n295);
    nand g1000(n816 ,n31[7] ,n666);
    dff g1001(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2169), .Q(n42[14]));
    nand g1002(n1265 ,n8[13] ,n849);
    nand g1003(n2286 ,n1915 ,n2183);
    nand g1004(n1365 ,n40[2] ,n1139);
    nand g1005(n1944 ,n2464 ,n1698);
    or g1006(n1883 ,n1782 ,n1683);
    nor g1007(n776 ,n422 ,n628);
    nand g1008(n1346 ,n810 ,n1005);
    nand g1009(n437 ,n35[2] ,n308);
    nand g1010(n2253 ,n1974 ,n2095);
    nand g1011(n1661 ,n841 ,n1426);
    nor g1012(n277 ,n262 ,n276);
    not g1013(n1562 ,n1509);
    not g1014(n246 ,n49[2]);
    nand g1015(n2290 ,n53[12] ,n2259);
    nand g1016(n610 ,n354 ,n586);
    not g1017(n1547 ,n1470);
    dff g1018(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2171), .Q(n42[5]));
    nand g1019(n545 ,n436 ,n393);
    nand g1020(n1995 ,n930 ,n1836);
    nand g1021(n749 ,n48[4] ,n527);
    nand g1022(n744 ,n48[1] ,n527);
    nand g1023(n709 ,n2442 ,n526);
    nand g1024(n2273 ,n1984 ,n2105);
    not g1025(n2397 ,n2409);
    nand g1026(n137 ,n51[10] ,n136);
    nand g1027(n1300 ,n42[20] ,n1139);
    or g1028(n2417 ,n55 ,n58);
    nand g1029(n2128 ,n25[1] ,n1693);
    or g1030(n1885 ,n1784 ,n1685);
    nand g1031(n2190 ,n2013 ,n2139);
    nand g1032(n549 ,n445 ,n400);
    nor g1033(n2456 ,n178 ,n176);
    or g1034(n1298 ,n552 ,n986);
    nand g1035(n1114 ,n825 ,n790);
    or g1036(n2177 ,n1494 ,n1999);
    dff g1037(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n908), .Q(n46[3]));
    not g1038(n202 ,n46[6]);
    dff g1039(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1206), .Q(n34[3]));
    nor g1040(n2435 ,n242 ,n244);
    dff g1041(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2250), .Q(n25[27]));
    nand g1042(n2121 ,n1714 ,n1713);
    nand g1043(n1612 ,n40[15] ,n1397);
    nand g1044(n1774 ,n946 ,n1469);
    xnor g1045(n2507 ,n50[7] ,n102);
    nand g1046(n934 ,n752 ,n662);
    nand g1047(n1380 ,n42[28] ,n1139);
    nand g1048(n898 ,n683 ,n732);
    nand g1049(n1637 ,n42[4] ,n289);
    not g1050(n171 ,n170);
    dff g1051(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2394), .Q(n45[0]));
    nand g1052(n1054 ,n13[10] ,n298);
    nand g1053(n1941 ,n2459 ,n1698);
    dff g1054(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2196), .Q(n26[15]));
    xnor g1055(n2466 ,n53[11] ,n193);
    or g1056(n1893 ,n1791 ,n1691);
    xnor g1057(n2481 ,n52[11] ,n165);
    nor g1058(n560 ,n39[2] ,n475);
    or g1059(n603 ,n563 ,n547);
    nand g1060(n810 ,n11[5] ,n293);
    nand g1061(n1322 ,n37[1] ,n1140);
    nand g1062(n1657 ,n835 ,n1422);
    nand g1063(n455 ,n52[8] ,n319);
    nand g1064(n2064 ,n2481 ,n1696);
    nand g1065(n1328 ,n35[1] ,n1140);
    nand g1066(n925 ,n11[30] ,n293);
    nand g1067(n95 ,n50[2] ,n94);
    nand g1068(n1816 ,n1226 ,n1551);
    nand g1069(n656 ,n49[8] ,n588);
    not g1070(n268 ,n267);
    or g1071(n1992 ,n852 ,n1702);
    not g1072(n539 ,n538);
    nand g1073(n2239 ,n51[7] ,n1991);
    nand g1074(n1658 ,n836 ,n1423);
    nand g1075(n2007 ,n26[24] ,n1695);
    nand g1076(n88 ,n49[7] ,n87);
    nand g1077(n722 ,n2420 ,n525);
    nand g1078(n1779 ,n1441 ,n1059);
    nand g1079(n2238 ,n51[8] ,n1991);
    nand g1080(n1137 ,n6[26] ,n296);
    nand g1081(n902 ,n16[8] ,n294);
    nand g1082(n1057 ,n5[31] ,n297);
    not g1083(n131 ,n130);
    nand g1084(n1665 ,n845 ,n1565);
    nand g1085(n1262 ,n6[12] ,n295);
    nand g1086(n769 ,n503 ,n600);
    nor g1087(n2505 ,n99 ,n101);
    nor g1088(n1142 ,n2407 ,n851);
    or g1089(n1851 ,n1732 ,n1650);
    dff g1090(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2391), .Q(n45[2]));
    not g1091(n307 ,n1397);
    nand g1092(n1125 ,n7[0] ,n847);
    nand g1093(n1052 ,n13[3] ,n297);
    nand g1094(n80 ,n48[6] ,n48[5]);
    nand g1095(n696 ,n46[6] ,n529);
    not g1096(n961 ,n919);
    nand g1097(n814 ,n11[4] ,n293);
    nand g1098(n781 ,n37[2] ,n665);
    nand g1099(n2293 ,n53[9] ,n2259);
    xnor g1100(n2489 ,n51[4] ,n125);
    nand g1101(n551 ,n448 ,n376);
    xnor g1102(n2433 ,n48[5] ,n238);
    nand g1103(n1718 ,n40[28] ,n291);
    nand g1104(n2072 ,n2473 ,n1696);
    dff g1105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2189), .Q(n26[22]));
    or g1106(n674 ,n333 ,n544);
    nand g1107(n2248 ,n1967 ,n2087);
    nor g1108(n361 ,n317 ,n53[0]);
    xnor g1109(n2462 ,n53[7] ,n186);
    nor g1110(n625 ,n2407 ,n560);
    nand g1111(n1223 ,n15[14] ,n300);
    nand g1112(n1378 ,n42[29] ,n292);
    nand g1113(n2288 ,n53[14] ,n2259);
    nand g1114(n2355 ,n1946 ,n2292);
    not g1115(n231 ,n48[2]);
    nand g1116(n1441 ,n42[3] ,n1139);
    dff g1117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1584), .Q(n29[1]));
    nor g1118(n112 ,n91 ,n111);
    nand g1119(n2112 ,n12[5] ,n1694);
    or g1120(n1913 ,n495 ,n1574);
    not g1121(n2140 ,n2014);
    nor g1122(n450 ,n335 ,n41[1]);
    nand g1123(n1739 ,n1125 ,n1374);
    nand g1124(n2216 ,n50[11] ,n1992);
    nand g1125(n2123 ,n1715 ,n1716);
    not g1126(n96 ,n95);
    nand g1127(n742 ,n34[8] ,n524);
    not g1128(n1522 ,n1427);
    not g1129(n94 ,n93);
    dff g1130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n796), .Q(n46[0]));
    dff g1131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1876), .Q(n42[10]));
    nand g1132(n1041 ,n4[0] ,n297);
    not g1133(n1422 ,n1381);
    nand g1134(n1825 ,n1186 ,n1542);
    nand g1135(n755 ,n34[2] ,n524);
    dff g1136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2281), .Q(n27));
    nand g1137(n929 ,n678 ,n644);
    nand g1138(n1455 ,n902 ,n1048);
    not g1139(n2160 ,n2057);
    nand g1140(n736 ,n2450 ,n528);
    nand g1141(n2131 ,n25[4] ,n1693);
    nor g1142(n1397 ,n533 ,n1146);
    nand g1143(n2322 ,n2078 ,n2235);
    not g1144(n1566 ,n1520);
    not g1145(n963 ,n921);
    not g1146(n1697 ,n1698);
    not g1147(n344 ,n45[1]);
    nand g1148(n1034 ,n4[13] ,n297);
    nand g1149(n1730 ,n1098 ,n1347);
    nand g1150(n2264 ,n2130 ,n2114);
    nand g1151(n1690 ,n1123 ,n1559);
    nor g1152(n369 ,n324 ,n50[6]);
    nand g1153(n1283 ,n6[22] ,n295);
    nand g1154(n1217 ,n9[26] ,n299);
    xnor g1155(n2437 ,n48[9] ,n245);
    xnor g1156(n2485 ,n52[15] ,n172);
    nand g1157(n1274 ,n6[18] ,n295);
    not g1158(n1413 ,n1346);
    nand g1159(n2256 ,n1975 ,n2096);
    nor g1160(n2475 ,n155 ,n157);
    not g1161(n175 ,n53[12]);
    nand g1162(n2032 ,n1620 ,n1619);
    nand g1163(n1115 ,n7[2] ,n295);
    nand g1164(n799 ,n11[12] ,n294);
    nand g1165(n654 ,n47[1] ,n587);
    nor g1166(n522 ,n368 ,n369);
    not g1167(n1538 ,n1456);
    nand g1168(n1714 ,n40[30] ,n1397);
    nand g1169(n1165 ,n15[11] ,n849);
    or g1170(n366 ,n319 ,n52[8]);
    nand g1171(n430 ,n52[15] ,n320);
    xnor g1172(n2450 ,n46[4] ,n206);
    nand g1173(n114 ,n50[13] ,n112);
    nand g1174(n782 ,n37[1] ,n665);
    nand g1175(n1103 ,n7[4] ,n295);
    dff g1176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1857), .Q(n42[27]));
    nand g1177(n574 ,n308 ,n482);
    dff g1178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1208), .Q(n34[1]));
    nand g1179(n805 ,n11[8] ,n293);
    nand g1180(n2404 ,n22[1] ,n2402);
    or g1181(n1868 ,n1765 ,n1668);
    not g1182(n1560 ,n1501);
    dff g1183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2273), .Q(n25[12]));
    nand g1184(n441 ,n53[13] ,n315);
    not g1185(n1555 ,n1491);
    not g1186(n2149 ,n2034);
    dff g1187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2173), .Q(n42[3]));
    nand g1188(n274 ,n34[6] ,n273);
    nand g1189(n454 ,n51[3] ,n322);
    nand g1190(n1343 ,n808 ,n1092);
    dff g1191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n874), .Q(n49[7]));
    dff g1192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2286), .Q(n51[0]));
    nand g1193(n2048 ,n1638 ,n1637);
    nand g1194(n2085 ,n12[31] ,n1694);
    nand g1195(n670 ,n38[2] ,n536);
    nand g1196(n2367 ,n2062 ,n2304);
    nand g1197(n281 ,n34[10] ,n280);
    nand g1198(n1184 ,n8[4] ,n849);
    nand g1199(n789 ,n39[1] ,n665);
    nor g1200(n506 ,n394 ,n405);
    nand g1201(n922 ,n748 ,n642);
    nand g1202(n845 ,n10[17] ,n294);
    or g1203(n857 ,n477 ,n674);
    nand g1204(n1674 ,n305 ,n1430);
    nand g1205(n1078 ,n9[12] ,n849);
    nand g1206(n1351 ,n1096 ,n1006);
    nand g1207(n471 ,n53[9] ,n313);
    nand g1208(n2214 ,n50[13] ,n1992);
    nand g1209(n1516 ,n795 ,n1031);
    nand g1210(n873 ,n716 ,n682);
    dff g1211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2371), .Q(n52[10]));
    dff g1212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1853), .Q(n40[1]));
    nor g1213(n1201 ,n2407 ,n966);
    nor g1214(n1192 ,n2407 ,n961);
    nand g1215(n640 ,n49[1] ,n588);
    nor g1216(n848 ,n675 ,n602);
    dff g1217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1350), .Q(n32[1]));
    nand g1218(n1189 ,n14[1] ,n296);
    not g1219(n1406 ,n1333);
    nand g1220(n1682 ,n932 ,n1531);
    not g1221(n1412 ,n1344);
    nand g1222(n255 ,n49[5] ,n254);
    dff g1223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2256), .Q(n25[21]));
    nor g1224(n1354 ,n2407 ,n1151);
    nand g1225(n2365 ,n2060 ,n2302);
    dff g1226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1932), .Q(n30[3]));
    nor g1227(n849 ,n2410 ,n700);
    nand g1228(n2110 ,n12[7] ,n1694);
    dff g1229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2268), .Q(n25[7]));
    nand g1230(n583 ,n425 ,n424);
    nand g1231(n1304 ,n41[12] ,n292);
    or g1232(n1909 ,n1809 ,n1706);
    nand g1233(n1187 ,n14[2] ,n296);
    dff g1234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2324), .Q(n51[8]));
    dff g1235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1910), .Q(n40[16]));
    nand g1236(n741 ,n2424 ,n525);
    nand g1237(n1072 ,n5[17] ,n848);
    nand g1238(n1010 ,n17[1] ,n848);
    nand g1239(n1132 ,n8[28] ,n299);
    xnor g1240(n507 ,n41[14] ,n50[14]);
    nand g1241(n788 ,n39[3] ,n665);
    nand g1242(n2413 ,n2406 ,n2404);
    nand g1243(n1254 ,n6[0] ,n296);
    nand g1244(n2031 ,n26[13] ,n1695);
    nand g1245(n715 ,n2438 ,n526);
    nand g1246(n463 ,n51[9] ,n313);
    nand g1247(n1342 ,n40[7] ,n1139);
    not g1248(n970 ,n929);
    dff g1249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1864), .Q(n42[18]));
    nor g1250(n1698 ,n535 ,n1398);
    nand g1251(n2325 ,n2080 ,n2239);
    nand g1252(n1120 ,n21[0] ,n300);
    dff g1253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1903), .Q(n40[23]));
    or g1254(n611 ,n357 ,n585);
    nand g1255(n2094 ,n12[23] ,n1694);
    nand g1256(n1587 ,n850 ,n1325);
    nor g1257(n1296 ,n497 ,n982);
    not g1258(n239 ,n238);
    dff g1259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2263), .Q(n25[2]));
    nand g1260(n1191 ,n15[0] ,n300);
    nand g1261(n2023 ,n26[17] ,n1695);
    nor g1262(n988 ,n583 ,n758);
    nand g1263(n1447 ,n1257 ,n1042);
    nand g1264(n2199 ,n2033 ,n2148);
    dff g1265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1581), .Q(n35[0]));
    nand g1266(n927 ,n725 ,n655);
    or g1267(n2165 ,n1371 ,n1922);
    nand g1268(n1804 ,n1225 ,n1482);
    not g1269(n1693 ,n1694);
    nand g1270(n2194 ,n2023 ,n2143);
    nand g1271(n1820 ,n1213 ,n1547);
    xnor g1272(n516 ,n41[5] ,n53[5]);
    nand g1273(n2113 ,n12[4] ,n1694);
    buf g1274(n32[7], 1'b0);
    nand g1275(n1134 ,n8[27] ,n300);
    nor g1276(n505 ,n409 ,n378);
    nand g1277(n2300 ,n53[2] ,n2259);
    xnor g1278(n2454 ,n46[8] ,n213);
    dff g1279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1855), .Q(n42[29]));
    nand g1280(n2130 ,n25[3] ,n1693);
    nand g1281(n1993 ,n25[5] ,n1693);
    nand g1282(n2392 ,n2388 ,n2390);
    nand g1283(n1315 ,n41[1] ,n1139);
    nand g1284(n2027 ,n26[15] ,n1695);
    or g1285(n1906 ,n1806 ,n1815);
    nand g1286(n835 ,n10[27] ,n664);
    nand g1287(n2297 ,n53[5] ,n2259);
    nand g1288(n2021 ,n2490 ,n1701);
    nand g1289(n998 ,n5[9] ,n297);
    or g1290(n1856 ,n1741 ,n1656);
    nand g1291(n153 ,n52[3] ,n152);
    nand g1292(n2221 ,n50[6] ,n1992);
    nand g1293(n1915 ,n332 ,n1701);
    nand g1294(n1991 ,n855 ,n1703);
    or g1295(n1908 ,n582 ,n1578);
    nand g1296(n1762 ,n1512 ,n1033);
    nand g1297(n478 ,n2[3] ,n2411);
    nand g1298(n195 ,n53[11] ,n194);
    nand g1299(n1968 ,n25[28] ,n1693);
    nand g1300(n1506 ,n952 ,n1262);
    not g1301(n295 ,n303);
    dff g1302(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2252), .Q(n25[25]));
    nand g1303(n660 ,n2527 ,n523);
    nand g1304(n1083 ,n6[2] ,n295);
    xnor g1305(n2492 ,n51[7] ,n130);
    nand g1306(n1473 ,n1215 ,n1061);
    nand g1307(n2037 ,n1626 ,n1692);
    dff g1308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1863), .Q(n42[19]));
    dff g1309(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2270), .Q(n25[18]));
    nand g1310(n1578 ,n501 ,n1318);
    nand g1311(n2010 ,n1598 ,n1597);
    nor g1312(n358 ,n317 ,n52[0]);
    nand g1313(n2369 ,n2064 ,n2306);
    nand g1314(n2405 ,n2415 ,n2410);
    nand g1315(n1390 ,n42[23] ,n292);
    nand g1316(n1491 ,n943 ,n1071);
    nand g1317(n910 ,n684 ,n728);
    nor g1318(n619 ,n2407 ,n519);
    dff g1319(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2172), .Q(n44[1]));
    nand g1320(n286 ,n34[13] ,n284);
    nand g1321(n1965 ,n25[31] ,n1693);
    nand g1322(n733 ,n2439 ,n526);
    not g1323(n1152 ,n1105);
    dff g1324(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2197), .Q(n26[14]));
    not g1325(n531 ,n532);
    nand g1326(n2295 ,n53[7] ,n2259);
    nand g1327(n1055 ,n13[1] ,n297);
    nand g1328(n2115 ,n12[2] ,n1694);
    nand g1329(n606 ,n341 ,n530);
    dff g1330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1887), .Q(n41[9]));
    nand g1331(n642 ,n2521 ,n523);
    dff g1332(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1198), .Q(n34[10]));
    nand g1333(n2016 ,n1605 ,n1604);
    nand g1334(n2388 ,n45[1] ,n2383);
    dff g1335(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2188), .Q(n26[23]));
    nand g1336(n806 ,n694 ,n734);
    nand g1337(n1653 ,n1122 ,n1418);
    nand g1338(n1707 ,n945 ,n1556);
    nand g1339(n2087 ,n12[29] ,n1694);
    nor g1340(n1701 ,n543 ,n1398);
    nand g1341(n711 ,n48[2] ,n527);
    nor g1342(n189 ,n174 ,n188);
    not g1343(n244 ,n243);
    nor g1344(n1143 ,n477 ,n772);
    nand g1345(n1667 ,n1269 ,n1563);
    or g1346(n1875 ,n1778 ,n1679);
    nand g1347(n2078 ,n2496 ,n1701);
    nor g1348(n2501 ,n94 ,n92);
    dff g1349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2320), .Q(n51[12]));
    nand g1350(n719 ,n2425 ,n525);
    nand g1351(n1649 ,n814 ,n1414);
    not g1352(n143 ,n142);
    or g1353(n1845 ,n1726 ,n1623);
    nor g1354(n2494 ,n134 ,n136);
    nand g1355(n913 ,n754 ,n661);
    nand g1356(n1489 ,n40[19] ,n292);
    nand g1357(n605 ,n340 ,n528);
    dff g1358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n31[2]));
    or g1359(n375 ,n328 ,n50[1]);
    nand g1360(n564 ,n312 ,n485);
    nand g1361(n2416 ,n2401 ,n2399);
    nand g1362(n1607 ,n40[18] ,n291);
    nand g1363(n2271 ,n1986 ,n2107);
    nand g1364(n2034 ,n1622 ,n1621);
    nand g1365(n1813 ,n1244 ,n1498);
    nand g1366(n1002 ,n5[14] ,n297);
    or g1367(n602 ,n2408 ,n532);
    nand g1368(n841 ,n10[21] ,n294);
    nor g1369(n1400 ,n572 ,n978);
    not g1370(n247 ,n49[6]);
    dff g1371(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2247), .Q(n25[30]));
    nand g1372(n1789 ,n1175 ,n1310);
    nand g1373(n2267 ,n1990 ,n2111);
    nand g1374(n1434 ,n868 ,n1041);
    nand g1375(n695 ,n2453 ,n528);
    dff g1376(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n899), .Q(n47[2]));
    nand g1377(n2043 ,n26[7] ,n1695);
    xnor g1378(n2518 ,n34[14] ,n286);
    nand g1379(n1589 ,n40[26] ,n291);
    dff g1380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1848), .Q(n40[5]));
    nor g1381(n1402 ,n570 ,n976);
    nand g1382(n1232 ,n7[20] ,n847);
    nor g1383(n493 ,n385 ,n397);
    nand g1384(n855 ,n308 ,n615);
    or g1385(n1857 ,n1742 ,n1657);
    nand g1386(n2408 ,n2[0] ,n2516);
    nand g1387(n236 ,n48[3] ,n234);
    not g1388(n331 ,n38[1]);
    nand g1389(n725 ,n34[3] ,n524);
    nand g1390(n198 ,n53[13] ,n196);
    nand g1391(n2192 ,n2017 ,n2141);
    nand g1392(n604 ,n338 ,n525);
    or g1393(n1905 ,n1807 ,n1814);
    nand g1394(n2051 ,n26[3] ,n1695);
    nand g1395(n2106 ,n12[11] ,n1694);
    nand g1396(n795 ,n10[16] ,n664);
    nand g1397(n2126 ,n1718 ,n1717);
    nand g1398(n1613 ,n801 ,n1407);
    nand g1399(n684 ,n47[9] ,n587);
    nand g1400(n434 ,n51[7] ,n327);
    nor g1401(n597 ,n358 ,n566);
    nand g1402(n1508 ,n42[13] ,n292);
    nor g1403(n133 ,n118 ,n132);
    nand g1404(n2224 ,n50[3] ,n1992);
    dff g1405(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2202), .Q(n26[9]));
    xnor g1406(n2520 ,n34[12] ,n283);
    nand g1407(n1924 ,n1144 ,n1744);
    xnor g1408(n2441 ,n47[4] ,n221);
    nand g1409(n1204 ,n7[30] ,n295);
    not g1410(n316 ,n41[4]);
    nand g1411(n991 ,n622 ,n303);
    dff g1412(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n875), .Q(n47[4]));
    not g1413(n1418 ,n1369);
    nand g1414(n1605 ,n40[19] ,n291);
    nand g1415(n1004 ,n4[7] ,n297);
    or g1416(n1846 ,n1727 ,n1624);
    not g1417(n1827 ,n1734);
    nor g1418(n372 ,n324 ,n52[6]);
    nand g1419(n1751 ,n36[2] ,n1402);
    dff g1420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2262), .Q(n25[1]));
    dff g1421(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1085), .Q(n34[13]));
    nor g1422(n1359 ,n2407 ,n1154);
    nand g1423(n577 ,n439 ,n435);
    nand g1424(n2412 ,n2405 ,n2403);
    xnor g1425(n2493 ,n51[8] ,n132);
    nand g1426(n2186 ,n2005 ,n2135);
    not g1427(n315 ,n41[13]);
    nand g1428(n581 ,n458 ,n446);
    not g1429(n293 ,n302);
    dff g1430(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1746), .Q(n37[2]));
    or g1431(n1865 ,n1757 ,n1665);
    dff g1432(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2230), .Q(n26[28]));
    nand g1433(n57 ,n20[0] ,n56);
    nand g1434(n2050 ,n1639 ,n1641);
    dff g1435(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1911), .Q(n40[15]));
    dff g1436(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2373), .Q(n52[7]));
    nand g1437(n1729 ,n1094 ,n1345);
    nor g1438(n60 ,n59 ,n2416);
    nand g1439(n1310 ,n41[6] ,n292);
    nand g1440(n1484 ,n939 ,n1067);
    not g1441(n2153 ,n2042);
    nor g1442(n594 ,n576 ,n549);
    nand g1443(n2242 ,n51[4] ,n1991);
    nand g1444(n2313 ,n1963 ,n2225);
    nand g1445(n1630 ,n40[8] ,n1397);
    nor g1446(n618 ,n2407 ,n521);
    nand g1447(n1956 ,n2508 ,n1700);
    dff g1448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1846), .Q(n40[8]));
    nand g1449(n1510 ,n30[2] ,n1141);
    nand g1450(n1056 ,n13[0] ,n297);
    dff g1451(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2353), .Q(n53[12]));
    nand g1452(n2377 ,n2072 ,n2314);
    nand g1453(n823 ,n31[1] ,n666);
    dff g1454(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n905), .Q(n46[6]));
    not g1455(n329 ,n43[1]);
    or g1456(n1841 ,n1723 ,n1595);
    nand g1457(n384 ,n41[3] ,n336);
    nand g1458(n170 ,n52[13] ,n168);
    nand g1459(n546 ,n438 ,n384);
    nand g1460(n2129 ,n25[2] ,n1693);
    or g1461(n374 ,n327 ,n50[7]);
    nand g1462(n1735 ,n1118 ,n1368);
    or g1463(n514 ,n312 ,n412);
    or g1464(n758 ,n382 ,n632);
    nor g1465(n1702 ,n669 ,n1293);
    nand g1466(n470 ,n35[0] ,n308);
    nand g1467(n2236 ,n51[10] ,n1991);
    nand g1468(n158 ,n52[6] ,n157);
    not g1469(n328 ,n41[1]);
    nand g1470(n731 ,n2441 ,n526);
    nand g1471(n1266 ,n6[14] ,n847);
    xnor g1472(n2430 ,n48[2] ,n233);
    or g1473(n376 ,n325 ,n52[2]);
    not g1474(n1542 ,n1460);
    not g1475(n2156 ,n2048);
    dff g1476(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1934), .Q(n29[3]));
    nor g1477(n664 ,n478 ,n532);
    nand g1478(n662 ,n2525 ,n523);
    dff g1479(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2339), .Q(n50[8]));
    nor g1480(n354 ,n43[1] ,n2[1]);
    or g1481(n2166 ,n1373 ,n1923);
    nand g1482(n1439 ,n807 ,n1040);
    nand g1483(n1309 ,n41[7] ,n1139);
    nand g1484(n56 ,n2419 ,n54);
    nand g1485(n2255 ,n1973 ,n2094);
    not g1486(n2138 ,n2010);
    nor g1487(n183 ,n53[5] ,n182);
    nand g1488(n1167 ,n15[10] ,n849);
    nand g1489(n997 ,n5[10] ,n298);
    dff g1490(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1904), .Q(n40[22]));
    nor g1491(n58 ,n2418 ,n57);
    dff g1492(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1860), .Q(n42[24]));
    nand g1493(n1513 ,n42[15] ,n1139);
    nand g1494(n1311 ,n41[5] ,n292);
    nand g1495(n1493 ,n40[17] ,n292);
    nand g1496(n1584 ,n303 ,n1326);
    nand g1497(n135 ,n51[9] ,n133);
    not g1498(n326 ,n41[12]);
    nand g1499(n221 ,n47[3] ,n219);
    or g1500(n669 ,n2407 ,n538);
    not g1501(n262 ,n34[8]);
    nand g1502(n410 ,n43[0] ,n308);
    nand g1503(n1812 ,n1247 ,n1502);
    nand g1504(n1210 ,n9[29] ,n299);
    nor g1505(n1579 ,n989 ,n1299);
    nand g1506(n1798 ,n1467 ,n1044);
    not g1507(n296 ,n303);
    nand g1508(n887 ,n702 ,n703);
    dff g1509(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1924), .Q(n37[3]));
    nand g1510(n1621 ,n42[11] ,n289);
    nand g1511(n1978 ,n25[18] ,n1693);
    nand g1512(n544 ,n330 ,n472);
    nor g1513(n978 ,n541 ,n856);
    nand g1514(n908 ,n697 ,n688);
    nand g1515(n1302 ,n41[14] ,n292);
    nand g1516(n1979 ,n25[17] ,n1693);
    dff g1517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1844), .Q(n40[10]));
    nor g1518(n2523 ,n278 ,n280);
    nand g1519(n1060 ,n5[28] ,n297);
    nand g1520(n2211 ,n2058 ,n2160);
    nor g1521(n256 ,n247 ,n255);
    not g1522(n1832 ,n1762);
    xnor g1523(n2503 ,n50[3] ,n95);
    xnor g1524(n2427 ,n49[8] ,n258);
    nor g1525(n529 ,n2407 ,n474);
    nand g1526(n1603 ,n40[20] ,n291);
    nand g1527(n1478 ,n40[25] ,n292);
    nand g1528(n453 ,n51[2] ,n325);
    nand g1529(n1495 ,n1239 ,n1073);
    nand g1530(n2305 ,n52[12] ,n2260);
    nand g1531(n1065 ,n5[24] ,n848);
    nand g1532(n2001 ,n26[27] ,n1695);
    not g1533(n1529 ,n1447);
    nand g1534(n482 ,n35[3] ,n2535);
    nand g1535(n1287 ,n8[24] ,n849);
    not g1536(n2139 ,n2012);
    nand g1537(n1738 ,n1129 ,n1376);
    nand g1538(n1949 ,n2515 ,n1700);
    dff g1539(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1669), .Q(n29[2]));
    nand g1540(n1033 ,n4[14] ,n298);
    nand g1541(n448 ,n52[11] ,n323);
    nor g1542(n1195 ,n2407 ,n957);
    nand g1543(n830 ,n10[5] ,n293);
    nand g1544(n1456 ,n1173 ,n1049);
    nor g1545(n977 ,n593 ,n856);
    nand g1546(n1022 ,n4[23] ,n298);
    nand g1547(n973 ,n757 ,n771);
    nand g1548(n2357 ,n1944 ,n2293);
    nand g1549(n864 ,n751 ,n636);
    nand g1550(n1628 ,n42[9] ,n289);
    nand g1551(n1648 ,n40[0] ,n291);
    nand g1552(n1109 ,n9[3] ,n299);
    nand g1553(n2315 ,n52[2] ,n2260);
    nand g1554(n1030 ,n4[17] ,n848);
    not g1555(n259 ,n258);
    nand g1556(n573 ,n461 ,n428);
    not g1557(n1417 ,n1366);
    dff g1558(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1909), .Q(n40[18]));
    nand g1559(n567 ,n482 ,n476);
    dff g1560(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2168), .Q(n42[22]));
    nand g1561(n436 ,n53[6] ,n324);
    nand g1562(n548 ,n471 ,n370);
    nand g1563(n875 ,n650 ,n731);
    not g1564(n1703 ,n1702);
    nand g1565(n784 ,n36[3] ,n665);
    nand g1566(n1290 ,n485 ,n858);
    nand g1567(n1984 ,n25[12] ,n1693);
    nand g1568(n1957 ,n2507 ,n1700);
    nand g1569(n1754 ,n36[1] ,n1403);
    or g1570(n1907 ,n1808 ,n1705);
    dff g1571(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2187), .Q(n26[24]));
    nor g1572(n587 ,n309 ,n487);
    nor g1573(n2527 ,n271 ,n273);
    nand g1574(n865 ,n11[31] ,n664);
    nor g1575(n396 ,n319 ,n53[8]);
    nor g1576(n2426 ,n257 ,n259);
    or g1577(n1894 ,n1792 ,n1625);
    nand g1578(n1645 ,n42[1] ,n289);
    not g1579(n2164 ,n2126);
    nand g1580(n1748 ,n1390 ,n1022);
    nor g1581(n148 ,n52[1] ,n52[0]);
    not g1582(n1409 ,n1338);
    not g1583(n110 ,n109);
    not g1584(n1533 ,n1451);
    nand g1585(n1606 ,n42[18] ,n289);
    nand g1586(n2013 ,n26[21] ,n1695);
    dff g1587(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1849), .Q(n40[4]));
    not g1588(n201 ,n46[2]);
    or g1589(n2169 ,n1511 ,n1931);
    nand g1590(n1475 ,n40[26] ,n292);
    dff g1591(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2165), .Q(n44[0]));
    nand g1592(n945 ,n11[16] ,n293);
    not g1593(n54 ,n20[1]);
    nand g1594(n1104 ,n816 ,n784);
    nand g1595(n1659 ,n837 ,n1424);
    nand g1596(n1620 ,n40[12] ,n1397);
    nand g1597(n885 ,n713 ,n699);
    or g1598(n770 ,n555 ,n598);
    nand g1599(n1760 ,n1268 ,n1513);
    not g1600(n1407 ,n1335);
    nand g1601(n1480 ,n40[24] ,n292);
    dff g1602(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2204), .Q(n26[7]));
    nand g1603(n427 ,n53[8] ,n319);
    nand g1604(n2274 ,n1983 ,n2104);
    nand g1605(n552 ,n464 ,n371);
    or g1606(n1882 ,n50[0] ,n1699);
    nor g1607(n1318 ,n553 ,n987);
    not g1608(n706 ,n527);
    nand g1609(n1073 ,n5[16] ,n297);
    nand g1610(n2092 ,n12[25] ,n1694);
    nand g1611(n2320 ,n2077 ,n2234);
    not g1612(n2161 ,n2119);
    nand g1613(n156 ,n52[5] ,n154);
    nand g1614(n1623 ,n804 ,n1409);
    nor g1615(n92 ,n50[1] ,n50[0]);
    nand g1616(n172 ,n52[14] ,n171);
    nand g1617(n2020 ,n1607 ,n1606);
    nand g1618(n1270 ,n6[16] ,n295);
    nand g1619(n1936 ,n2467 ,n1698);
    nand g1620(n1130 ,n8[29] ,n300);
    dff g1621(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1568), .Q(n28));
    dff g1622(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2313), .Q(n50[2]));
    nor g1623(n521 ,n345 ,n349);
    nor g1624(n503 ,n407 ,n387);
    dff g1625(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2166), .Q(n42[31]));
    not g1626(n2157 ,n2050);
    nand g1627(n1618 ,n42[13] ,n289);
    nand g1628(n1518 ,n1273 ,n1030);
    nand g1629(n1773 ,n1436 ,n1045);
    nand g1630(n456 ,n51[8] ,n319);
    nand g1631(n832 ,n10[30] ,n294);
    or g1632(n543 ,n477 ,n415);
    nand g1633(n1313 ,n41[3] ,n1139);
    nand g1634(n1193 ,n14[0] ,n295);
    not g1635(n159 ,n158);
    nand g1636(n1040 ,n4[4] ,n848);
    nand g1637(n860 ,n627 ,n672);
    nand g1638(n1008 ,n5[2] ,n297);
    nand g1639(n2212 ,n50[15] ,n1992);
    not g1640(n1539 ,n1457);
    nand g1641(n1652 ,n826 ,n1417);
    nand g1642(n1035 ,n4[12] ,n298);
    xnor g1643(n2488 ,n51[3] ,n123);
    nand g1644(n2277 ,n1980 ,n2101);
    nand g1645(n1067 ,n5[22] ,n297);
    nand g1646(n1488 ,n40[20] ,n1139);
    nand g1647(n1229 ,n9[21] ,n849);
    or g1648(n393 ,n321 ,n53[10]);
    nand g1649(n2289 ,n53[13] ,n2259);
    dff g1650(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1856), .Q(n42[28]));
    not g1651(n164 ,n163);
    dff g1652(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2335), .Q(n50[11]));
    nand g1653(n1027 ,n4[20] ,n297);
    or g1654(n2414 ,n60 ,n63);
    nand g1655(n2349 ,n2282 ,n1918);
    nor g1656(n1917 ,n1576 ,n1575);
    nand g1657(n1486 ,n40[21] ,n1139);
    nand g1658(n1710 ,n42[31] ,n289);
    nand g1659(n894 ,n744 ,n743);
    nand g1660(n2262 ,n2128 ,n2116);
    nand g1661(n2044 ,n1634 ,n1633);
    not g1662(n473 ,n474);
    nand g1663(n787 ,n36[0] ,n665);
    nand g1664(n260 ,n49[8] ,n259);
    nand g1665(n1174 ,n14[7] ,n295);
    nand g1666(n2193 ,n2018 ,n2142);
    nand g1667(n2415 ,n2400 ,n2398);
    nand g1668(n248 ,n49[1] ,n49[0]);
    nand g1669(n826 ,n11[1] ,n293);
    nand g1670(n663 ,n47[8] ,n587);
    nand g1671(n2045 ,n26[6] ,n1695);
    nand g1672(n1326 ,n29[1] ,n1140);
    dff g1673(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n887), .Q(n48[6]));
    nand g1674(n1362 ,n824 ,n1008);
    nand g1675(n909 ,n16[6] ,n664);
    nand g1676(n165 ,n52[10] ,n164);
    nand g1677(n1170 ,n14[9] ,n296);
    nand g1678(n2235 ,n51[11] ,n1991);
    nand g1679(n582 ,n453 ,n452);
    nand g1680(n238 ,n48[4] ,n237);
    nand g1681(n432 ,n51[6] ,n324);
    nand g1682(n550 ,n417 ,n401);
    dff g1683(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1891), .Q(n41[6]));
    nor g1684(n773 ,n467 ,n599);
    nand g1685(n924 ,n742 ,n681);
    nand g1686(n1166 ,n14[11] ,n295);
    or g1687(n2170 ,n1506 ,n1933);
    nand g1688(n980 ,n508 ,n776);
    or g1689(n1884 ,n1783 ,n1684);
    nand g1690(n1811 ,n1240 ,n1496);
    not g1691(n1416 ,n1362);
    nand g1692(n1466 ,n40[30] ,n292);
    or g1693(n1859 ,n1745 ,n1659);
    dff g1694(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n898), .Q(n47[3]));
    nor g1695(n390 ,n326 ,n51[12]);
    dff g1696(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1354), .Q(n31[7]));
    nand g1697(n1394 ,n1281 ,n1026);
    nand g1698(n892 ,n711 ,n747);
    dff g1699(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1851), .Q(n40[3]));
    nor g1700(n559 ,n39[3] ,n483);
    nand g1701(n568 ,n444 ,n465);
    nand g1702(n1502 ,n40[14] ,n292);
    nand g1703(n1111 ,n822 ,n794);
    not g1704(n192 ,n191);
    or g1705(n1895 ,n1793 ,n1825);
    not g1706(n1414 ,n1351);
    or g1707(n1570 ,n301 ,n1403);
    dff g1708(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2377), .Q(n52[3]));
    nand g1709(n1737 ,n1372 ,n1013);
    not g1710(n1535 ,n1453);
    dff g1711(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2348), .Q(n52[0]));
    or g1712(n1863 ,n1755 ,n1663);
    dff g1713(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1867), .Q(n42[15]));
    nor g1714(n588 ,n310 ,n486);
    nand g1715(n1020 ,n4[24] ,n848);
    nand g1716(n2009 ,n26[23] ,n1695);
    dff g1717(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2327), .Q(n51[5]));
    nand g1718(n2040 ,n1630 ,n1629);
    nand g1719(n1740 ,n1131 ,n1378);
    nor g1720(n537 ,n38[0] ,n477);
    xnor g1721(n2432 ,n48[4] ,n236);
    nor g1722(n536 ,n38[0] ,n414);
    nand g1723(n1744 ,n37[3] ,n1399);
    nand g1724(n1633 ,n42[6] ,n289);
    nand g1725(n569 ,n454 ,n431);
    nand g1726(n1958 ,n2458 ,n1698);
    dff g1727(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n617), .Q(n33[5]));
    dff g1728(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1912), .Q(n40[14]));
    or g1729(n1877 ,n1772 ,n1680);
    dff g1730(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1854), .Q(n42[30]));
    nand g1731(n2077 ,n2497 ,n1701);
    dff g1732(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1890), .Q(n41[5]));
    dff g1733(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1872), .Q(n42[7]));
    nor g1734(n154 ,n145 ,n153);
    nand g1735(n1341 ,n1279 ,n1027);
    or g1736(n1569 ,n2407 ,n1400);
    not g1737(n2133 ,n2000);
    nand g1738(n666 ,n43[1] ,n542);
    nand g1739(n2195 ,n2025 ,n2144);
    nor g1740(n140 ,n119 ,n139);
    xnor g1741(n2470 ,n53[15] ,n200);
    nand g1742(n2011 ,n26[22] ,n1695);
    not g1743(n1838 ,n1802);
    dff g1744(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2344), .Q(n50[4]));
    nand g1745(n2362 ,n1958 ,n2299);
    nand g1746(n1687 ,n897 ,n1536);
    nand g1747(n1970 ,n25[26] ,n1693);
    xnor g1748(n2445 ,n47[8] ,n228);
    dff g1749(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1160), .Q(n34[4]));
    nand g1750(n2257 ,n1976 ,n2097);
    nand g1751(n1396 ,n40[8] ,n292);
    nand g1752(n163 ,n52[9] ,n161);
    dff g1753(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1889), .Q(n41[7]));
    nor g1754(n387 ,n323 ,n51[11]);
    xnor g1755(n2530 ,n34[2] ,n265);
    nand g1756(n641 ,n49[2] ,n588);
    nor g1757(n979 ,n500 ,n759);
    nor g1758(n182 ,n173 ,n181);
    not g1759(n592 ,n591);
    nand g1760(n1221 ,n9[24] ,n299);
    nand g1761(n2024 ,n1611 ,n1610);
    nand g1762(n868 ,n10[0] ,n293);
    xnor g1763(n2495 ,n51[10] ,n135);
    nand g1764(n591 ,n2410 ,n478);
    nor g1765(n190 ,n53[9] ,n189);
    nand g1766(n1026 ,n4[21] ,n297);
    nand g1767(n1086 ,n7[10] ,n847);
    nand g1768(n2091 ,n12[26] ,n1694);
    not g1769(n136 ,n135);
    nand g1770(n949 ,n16[5] ,n293);
    nand g1771(n831 ,n10[31] ,n294);
    nand g1772(n2269 ,n1988 ,n2109);
    nand g1773(n1824 ,n1189 ,n1543);
    or g1774(n404 ,n316 ,n51[4]);
    not g1775(n291 ,n307);
    dff g1776(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2209), .Q(n26[2]));
    nand g1777(n1113 ,n9[2] ,n299);
    nand g1778(n125 ,n51[3] ,n124);
    nand g1779(n2038 ,n1627 ,n1628);
    not g1780(n301 ,n308);
    nand g1781(n1980 ,n25[16] ,n1693);
    dff g1782(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2345), .Q(n50[3]));
    nand g1783(n2409 ,n2[1] ,n2417);
    dff g1784(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n651), .Q(n39[3]));
    nand g1785(n1786 ,n1170 ,n1307);
    nand g1786(n681 ,n2524 ,n523);
    nand g1787(n476 ,n35[2] ,n2534);
    nor g1788(n409 ,n322 ,n51[3]);
    nor g1789(n162 ,n52[9] ,n161);
    nand g1790(n809 ,n11[6] ,n293);
    nand g1791(n1487 ,n941 ,n1069);
    not g1792(n1419 ,n1375);
    nand g1793(n1763 ,n861 ,n1510);
    nand g1794(n798 ,n685 ,n736);
    nand g1795(n746 ,n34[10] ,n524);
    not g1796(n2163 ,n2123);
    or g1797(n489 ,n364 ,n386);
    nand g1798(n107 ,n50[9] ,n105);
    nor g1799(n1205 ,n2407 ,n967);
    not g1800(n2147 ,n2030);
    nand g1801(n1000 ,n5[8] ,n848);
    nand g1802(n1684 ,n1164 ,n1533);
    nand g1803(n2093 ,n12[24] ,n1694);
    nor g1804(n2431 ,n235 ,n237);
    not g1805(n411 ,n410);
    nand g1806(n1781 ,n1084 ,n1302);
    nand g1807(n1609 ,n42[17] ,n289);
    not g1808(n103 ,n102);
    nand g1809(n819 ,n11[3] ,n294);
    dff g1810(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1901), .Q(n40[27]));
    nand g1811(n558 ,n365 ,n430);
    nand g1812(n946 ,n10[10] ,n664);
    nand g1813(n1752 ,n1280 ,n1395);
    nand g1814(n1588 ,n42[26] ,n289);
    nor g1815(n270 ,n261 ,n269);
    nand g1816(n1327 ,n35[0] ,n1142);
    nand g1817(n883 ,n723 ,n705);
    nor g1818(n617 ,n2407 ,n518);
    nand g1819(n1929 ,n1570 ,n1754);
    nand g1820(n870 ,n10[8] ,n294);
    nand g1821(n1062 ,n5[26] ,n298);
    nand g1822(n1795 ,n797 ,n1316);
    nand g1823(n717 ,n2428 ,n525);
    nand g1824(n1175 ,n14[6] ,n295);
    dff g1825(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n910), .Q(n47[9]));
    nand g1826(n144 ,n51[14] ,n143);
    nand g1827(n1725 ,n1086 ,n1336);
    nand g1828(n1680 ,n1250 ,n1525);
    dff g1829(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n616), .Q(n33[6]));
    nand g1830(n2243 ,n51[3] ,n1991);
    nand g1831(n1601 ,n800 ,n1406);
    nor g1832(n398 ,n325 ,n53[2]);
    nand g1833(n1443 ,n42[2] ,n1139);
    nor g1834(n672 ,n567 ,n584);
    nand g1835(n914 ,n16[4] ,n294);
    dff g1836(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n886), .Q(n48[7]));
    nand g1837(n1982 ,n25[14] ,n1693);
    nor g1838(n1200 ,n2407 ,n965);
    nand g1839(n584 ,n480 ,n474);
    nand g1840(n1197 ,n9[31] ,n299);
    nand g1841(n2356 ,n1938 ,n2295);
    dff g1842(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1583), .Q(n30[1]));
    or g1843(n399 ,n318 ,n53[14]);
    nand g1844(n2308 ,n52[9] ,n2260);
    dff g1845(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2341), .Q(n50[6]));
    nand g1846(n1676 ,n1255 ,n1526);
    or g1847(n859 ,n589 ,n668);
    nand g1848(n1952 ,n2512 ,n1700);
    nand g1849(n1090 ,n7[8] ,n295);
    not g1850(n1532 ,n1450);
    nand g1851(n206 ,n46[3] ,n204);
    nand g1852(n2294 ,n53[8] ,n2259);
    nor g1853(n1317 ,n2407 ,n1245);
    nand g1854(n1617 ,n40[13] ,n1397);
    nand g1855(n1392 ,n42[22] ,n1139);
    nand g1856(n836 ,n10[26] ,n664);
    not g1857(n1557 ,n1497);
    nand g1858(n66 ,n2413 ,n64);
    nand g1859(n638 ,n49[0] ,n588);
    nand g1860(n726 ,n48[3] ,n527);
    dff g1861(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n624), .Q(n39[1]));
    nand g1862(n2334 ,n1951 ,n2214);
    nand g1863(n2303 ,n52[14] ,n2260);
    nand g1864(n1227 ,n7[22] ,n847);
    nand g1865(n627 ,n472 ,n564);
    not g1866(n966 ,n924);
    nand g1867(n839 ,n10[22] ,n293);
    nand g1868(n1683 ,n881 ,n1532);
    nand g1869(n2226 ,n50[1] ,n1992);
    nand g1870(n1238 ,n7[17] ,n295);
    nand g1871(n1496 ,n40[16] ,n292);
    not g1872(n224 ,n223);
    nor g1873(n235 ,n48[3] ,n234);
    nand g1874(n750 ,n34[14] ,n524);
    not g1875(n1148 ,n1100);
    nand g1876(n2097 ,n12[20] ,n1694);
    xnor g1877(n2480 ,n52[10] ,n163);
    not g1878(n232 ,n48[6]);
    or g1879(n1898 ,n1796 ,n1822);
    nand g1880(n1576 ,n983 ,n1296);
    xnor g1881(n2467 ,n53[12] ,n195);
    nand g1882(n1061 ,n5[27] ,n848);
    nand g1883(n1483 ,n40[22] ,n1139);
    xnor g1884(n2439 ,n47[2] ,n218);
    nand g1885(n2310 ,n52[7] ,n2260);
    nand g1886(n1382 ,n42[27] ,n292);
    nand g1887(n1519 ,n42[18] ,n292);
    nand g1888(n2075 ,n2499 ,n1701);
    nand g1889(n1715 ,n40[29] ,n291);
    nand g1890(n1051 ,n13[4] ,n848);
    nand g1891(n659 ,n49[7] ,n588);
    nor g1892(n2531 ,n266 ,n264);
    nand g1893(n1081 ,n7[11] ,n296);
    nand g1894(n445 ,n50[2] ,n325);
    nand g1895(n1248 ,n9[13] ,n299);
    nand g1896(n442 ,n50[6] ,n324);
    xnor g1897(n2434 ,n48[6] ,n240);
    nand g1898(n844 ,n10[18] ,n293);
    nand g1899(n878 ,n756 ,n717);
    dff g1900(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2340), .Q(n50[7]));
    not g1901(n335 ,n51[1]);
    nand g1902(n987 ,n490 ,n777);
    nand g1903(n1123 ,n15[6] ,n299);
    nor g1904(n2532 ,n70 ,n73);
    nand g1905(n2185 ,n2002 ,n2134);
    nor g1906(n2181 ,n769 ,n1908);
    nand g1907(n1472 ,n860 ,n1145);
    nand g1908(n1261 ,n8[11] ,n299);
    nand g1909(n866 ,n10[6] ,n293);
    nand g1910(n1796 ,n1199 ,n1464);
    nand g1911(n1727 ,n1090 ,n1396);
    nor g1912(n2519 ,n285 ,n287);
    xnor g1913(n2511 ,n50[11] ,n109);
    nand g1914(n1783 ,n884 ,n1304);
    nand g1915(n882 ,n640 ,n722);
    nand g1916(n1433 ,n867 ,n1075);
    nand g1917(n1954 ,n2510 ,n1700);
    dff g1918(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2261), .Q(n25[0]));
    not g1919(n118 ,n51[8]);
    dff g1920(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2356), .Q(n53[7]));
    nand g1921(n1272 ,n6[17] ,n847);
    nand g1922(n1765 ,n1264 ,n1508);
    nand g1923(n487 ,n35[1] ,n308);
    nor g1924(n79 ,n48[4] ,n48[3]);
    not g1925(n157 ,n156);
    nand g1926(n1374 ,n40[0] ,n1139);
    xnor g1927(n2525 ,n34[7] ,n274);
    nor g1928(n983 ,n513 ,n766);
    dff g1929(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2186), .Q(n26[25]));
    xnor g1930(n2478 ,n52[8] ,n160);
    nand g1931(n807 ,n10[4] ,n293);
    not g1932(n1553 ,n1487);
    or g1933(n2171 ,n1438 ,n1947);
    dff g1934(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n951), .Q(n46[2]));
    nand g1935(n895 ,n646 ,n712);
    xnor g1936(n491 ,n41[13] ,n51[13]);
    nand g1937(n822 ,n31[2] ,n666);
    dff g1938(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1877), .Q(n42[0]));
    nand g1939(n1428 ,n42[6] ,n292);
    or g1940(n2168 ,n1393 ,n1926);
    nand g1941(n1468 ,n1210 ,n1209);
    not g1942(n166 ,n165);
    nand g1943(n1006 ,n5[4] ,n297);
    nand g1944(n2342 ,n1960 ,n2222);
    nand g1945(n1260 ,n6[11] ,n296);
    nand g1946(n1246 ,n9[14] ,n299);
    dff g1947(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1869), .Q(n42[11]));
    nand g1948(n576 ,n429 ,n418);
    nand g1949(n1749 ,n36[3] ,n1401);
    nand g1950(n707 ,n46[2] ,n529);
    not g1951(n207 ,n206);
    nand g1952(n2116 ,n12[1] ,n1694);
    nand g1953(n1258 ,n15[15] ,n300);
    nand g1954(n1127 ,n8[31] ,n849);
    nand g1955(n1015 ,n4[29] ,n297);
    nor g1956(n761 ,n590 ,n670);
    nand g1957(n73 ,n46[7] ,n72);
    nand g1958(n825 ,n31[0] ,n666);
    nand g1959(n452 ,n51[4] ,n316);
    dff g1960(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1893), .Q(n41[4]));
    nand g1961(n1333 ,n1080 ,n996);
    nand g1962(n1453 ,n893 ,n1054);
    nand g1963(n2204 ,n2043 ,n2153);
    nand g1964(n2229 ,n2124 ,n2163);
    nand g1965(n1951 ,n2513 ,n1700);
    or g1966(n1571 ,n301 ,n1402);
    nor g1967(n596 ,n551 ,n550);
    nand g1968(n646 ,n47[7] ,n587);
    nand g1969(n2219 ,n50[8] ,n1992);
    nand g1970(n1383 ,n1136 ,n1018);
    nand g1971(n644 ,n2531 ,n523);
    nand g1972(n739 ,n34[5] ,n524);
    dff g1973(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2277), .Q(n25[16]));
    nand g1974(n428 ,n3[0] ,n311);
    nand g1975(n900 ,n656 ,n693);
    dff g1976(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n863), .Q(n49[4]));
    nand g1977(n621 ,n38[2] ,n532);
    nand g1978(n208 ,n46[4] ,n207);
    or g1979(n2176 ,n1476 ,n1997);
    not g1980(n318 ,n41[14]);
    dff g1981(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1885), .Q(n41[11]));
    nand g1982(n2206 ,n2047 ,n2155);
    nor g1983(n1085 ,n2407 ,n963);
    not g1984(n1408 ,n1337);
    nand g1985(n1263 ,n8[12] ,n300);
    or g1986(n1850 ,n1733 ,n1651);
    nor g1987(n2180 ,n1913 ,n1916);
    nand g1988(n1209 ,n7[29] ,n295);
    nand g1989(n1521 ,n42[19] ,n292);
    nor g1990(n614 ,n545 ,n520);
    dff g1991(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1862), .Q(n42[20]));
    nand g1992(n937 ,n11[24] ,n294);
    or g1993(n2280 ,n1917 ,n2180);
    nand g1994(n686 ,n34[13] ,n524);
    nand g1995(n2361 ,n1941 ,n2298);
    dff g1996(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1289), .Q(n34[6]));
    dff g1997(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n31[5]));
    nand g1998(n1095 ,n9[5] ,n299);
    nand g1999(n1182 ,n6[7] ,n847);
    nand g2000(n1761 ,n30[3] ,n1399);
    nand g2001(n1011 ,n5[0] ,n297);
    nand g2002(n1164 ,n14[12] ,n296);
    nand g2003(n1724 ,n1081 ,n1334);
    nand g2004(n1039 ,n4[6] ,n297);
    nand g2005(n1368 ,n40[1] ,n292);
    nand g2006(n2312 ,n52[5] ,n2260);
    nand g2007(n1096 ,n9[4] ,n299);
    nand g2008(n629 ,n427 ,n534);
    or g2009(n352 ,n36[2] ,n36[3]);
    nand g2010(n1679 ,n1203 ,n1528);
    nand g2011(n1146 ,n337 ,n858);
    or g2012(n590 ,n312 ,n479);
    nand g2013(n1214 ,n7[28] ,n295);
    nand g2014(n1082 ,n9[10] ,n300);
    nand g2015(n1141 ,n669 ,n855);
    nor g2016(n2382 ,n306 ,n2381);
    nand g2017(n2410 ,n2[2] ,n2414);
    nand g2018(n451 ,n51[15] ,n320);
    nand g2019(n1642 ,n42[2] ,n289);
    dff g2020(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2369), .Q(n52[11]));
    nand g2021(n215 ,n46[8] ,n214);
    dff g2022(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1930), .Q(n36[0]));
    xnor g2023(n2457 ,n53[2] ,n177);
    nand g2024(n2344 ,n1961 ,n2223);
    nand g2025(n1627 ,n40[9] ,n291);
    or g2026(n764 ,n565 ,n603);
    dff g2027(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2323), .Q(n51[10]));
    nand g2028(n2374 ,n2069 ,n2311);
    nand g2029(n1108 ,n821 ,n788);
    nor g2030(n204 ,n201 ,n203);
    not g2031(n138 ,n137);
    nor g2032(n2385 ,n488 ,n2383);
    nand g2033(n1277 ,n8[19] ,n299);
    dff g2034(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1875), .Q(n42[1]));
    xnor g2035(n2436 ,n48[8] ,n243);
    nor g2036(n504 ,n408 ,n383);
    nand g2037(n797 ,n16[0] ,n294);
    nand g2038(n1230 ,n7[21] ,n296);
    nand g2039(n2218 ,n50[9] ,n1992);
    nand g2040(n1336 ,n40[10] ,n292);
    nand g2041(n1507 ,n42[12] ,n1139);
    nand g2042(n1994 ,n2469 ,n1698);
    nand g2043(n1444 ,n871 ,n1043);
    not g2044(n1537 ,n1455);
    nor g2045(n469 ,n344 ,n301);
    nand g2046(n901 ,n654 ,n715);
    nand g2047(n1591 ,n42[25] ,n289);
    nor g2048(n985 ,n498 ,n768);
    not g2049(n287 ,n286);
    nand g2050(n1802 ,n1478 ,n1063);
    nand g2051(n1501 ,n1248 ,n1076);
    nand g2052(n2036 ,n26[10] ,n1695);
    not g2053(n535 ,n534);
    nand g2054(n1159 ,n6[1] ,n847);
    dff g2055(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1582), .Q(n37[1]));
    nand g2056(n1335 ,n1082 ,n997);
    dff g2057(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1674), .Q(n35[2]));
    dff g2058(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1880), .Q(n41[14]));
    dff g2059(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n32[2]));
    not g2060(n1415 ,n1356);
    nand g2061(n1717 ,n42[28] ,n289);
    nand g2062(n2258 ,n2056 ,n2159);
    nand g2063(n633 ,n2519 ,n523);
    nand g2064(n2389 ,n860 ,n2384);
    not g2065(n333 ,n44[1]);
    nand g2066(n1306 ,n41[10] ,n1139);
    nor g2067(n2449 ,n205 ,n207);
    nand g2068(n1331 ,n1078 ,n995);
    nand g2069(n1914 ,n334 ,n1696);
    not g2070(n965 ,n923);
    dff g2071(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n31[1]));
    not g2072(n1549 ,n1479);
    not g2073(n334 ,n52[0]);
    or g2074(n355 ,n35[0] ,n35[3]);
    nor g2075(n383 ,n325 ,n51[2]);
    nand g2076(n83 ,n48[7] ,n82);
    nand g2077(n1750 ,n1392 ,n1025);
    not g2078(n2144 ,n2024);
    buf g2079(n32[4], 1'b0);
    nor g2080(n220 ,n47[3] ,n219);
    nand g2081(n877 ,n663 ,n729);
    nand g2082(n801 ,n11[10] ,n293);
    not g2083(n322 ,n41[3]);
    nand g2084(n1019 ,n4[25] ,n848);
    nand g2085(n718 ,n2426 ,n525);
    nand g2086(n2107 ,n12[10] ,n1694);
    nand g2087(n85 ,n49[6] ,n49[5]);
    nand g2088(n2373 ,n2068 ,n2310);
    not g2089(n1153 ,n1106);
    nand g2090(n2213 ,n50[14] ,n1992);
    nand g2091(n2100 ,n12[17] ,n1694);
    or g2092(n541 ,n38[0] ,n484);
    xnor g2093(n511 ,n41[12] ,n52[12]);
    nand g2094(n2354 ,n1937 ,n2291);
    nand g2095(n2254 ,n1972 ,n2093);
    nand g2096(n2376 ,n2071 ,n2346);
    nand g2097(n1708 ,n947 ,n1557);
    nand g2098(n2250 ,n1969 ,n2090);
    xnor g2099(n2497 ,n51[12] ,n139);
    nand g2100(n1514 ,n955 ,n1032);
    nor g2101(n993 ,n578 ,n763);
    nand g2102(n635 ,n2517 ,n523);
    nand g2103(n2324 ,n2054 ,n2238);
    nand g2104(n1340 ,n1089 ,n1000);
    not g2105(n2142 ,n2020);
    nand g2106(n2364 ,n1945 ,n2301);
    nand g2107(n2230 ,n2125 ,n2164);
    dff g2108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2275), .Q(n25[14]));
    nand g2109(n840 ,n641 ,n721);
    nand g2110(n2084 ,n2486 ,n1701);
    nand g2111(n415 ,n311 ,n330);
    nor g2112(n976 ,n541 ,n857);
    nand g2113(n926 ,n739 ,n660);
    nand g2114(n130 ,n51[6] ,n129);
    nand g2115(n423 ,n53[7] ,n327);
    not g2116(n1561 ,n1505);
    nand g2117(n1933 ,n1263 ,n1833);
    nand g2118(n1574 ,n494 ,n1320);
    nand g2119(n1163 ,n15[12] ,n849);
    nor g2120(n249 ,n246 ,n248);
    nand g2121(n570 ,n308 ,n476);
    or g2122(n986 ,n558 ,n760);
    nand g2123(n2244 ,n51[2] ,n1991);
    nand g2124(n1731 ,n1103 ,n1353);
    not g2125(n1556 ,n1495);
    nand g2126(n1459 ,n1183 ,n1052);
    nand g2127(n2090 ,n12[27] ,n1694);
    or g2128(n392 ,n327 ,n51[7]);
    or g2129(n1852 ,n1739 ,n1653);
    nand g2130(n699 ,n2436 ,n530);
    dff g2131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n991), .Q(n38[1]));
    nor g2132(n205 ,n46[3] ,n204);
    nand g2133(n1180 ,n15[4] ,n299);
    nand g2134(n1927 ,n1572 ,n1749);
    nand g2135(n2245 ,n51[1] ,n1991);
    nand g2136(n2004 ,n1590 ,n1591);
    nand g2137(n1308 ,n41[8] ,n292);
    dff g2138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2359), .Q(n53[6]));
    or g2139(n2167 ,n1391 ,n1925);
    nor g2140(n542 ,n43[0] ,n472);
    xnor g2141(n509 ,n41[10] ,n50[10]);
    nand g2142(n100 ,n50[5] ,n98);
    not g2143(n1543 ,n1461);
    nor g2144(n1355 ,n2407 ,n1152);
    nand g2145(n827 ,n23[1] ,n664);
    nand g2146(n2104 ,n12[13] ,n1694);
    nand g2147(n1377 ,n1130 ,n1015);
    nand g2148(n1016 ,n4[28] ,n298);
    nand g2149(n1059 ,n4[3] ,n298);
    nand g2150(n1107 ,n820 ,n787);
    nand g2151(n1675 ,n1182 ,n1523);
    nand g2152(n2076 ,n2498 ,n1701);
    nand g2153(n75 ,n47[6] ,n47[5]);
    nand g2154(n930 ,n11[29] ,n293);
    nand g2155(n1503 ,n42[11] ,n1139);
    or g2156(n367 ,n313 ,n50[9]);
    dff g2157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1888), .Q(n41[8]));
    nand g2158(n1371 ,n1121 ,n1012);
    nand g2159(n1314 ,n41[2] ,n292);
    nand g2160(n2319 ,n2076 ,n2233);
    nand g2161(n1093 ,n7[6] ,n295);
    xnor g2162(n2514 ,n50[14] ,n114);
    not g2163(n1424 ,n1385);
    nand g2164(n1688 ,n1171 ,n1537);
    nand g2165(n932 ,n16[14] ,n293);
    not g2166(n310 ,n2535);
    nand g2167(n167 ,n52[11] ,n166);
    nand g2168(n1461 ,n918 ,n1055);
    dff g2169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2378), .Q(n52[1]));
    not g2170(n1420 ,n1377);
    nand g2171(n1044 ,n5[29] ,n298);
    dff g2172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2175), .Q(n40[26]));
    not g2173(n1530 ,n1448);
    dff g2174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2254), .Q(n25[24]));
    nand g2175(n1759 ,n1270 ,n1515);
    nand g2176(n1963 ,n2502 ,n1700);
    or g2177(n1919 ,n301 ,n1696);
    nand g2178(n1819 ,n933 ,n1548);
    nand g2179(n850 ,n536 ,n667);
    nand g2180(n1009 ,n5[1] ,n298);
    nor g2181(n106 ,n50[9] ,n105);
    nand g2182(n1222 ,n7[24] ,n296);
    dff g2183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1228), .Q(n34[7]));
    nand g2184(n2203 ,n2041 ,n2152);
    nand g2185(n599 ,n379 ,n515);
    not g2186(n2407 ,n1);
    or g2187(n1864 ,n1756 ,n1664);
    or g2188(n981 ,n568 ,n764);
    nand g2189(n1815 ,n940 ,n1552);
    nand g2190(n1619 ,n42[12] ,n289);
    nand g2191(n532 ,n411 ,n412);
    dff g2192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1360), .Q(n31[3]));
    nand g2193(n2252 ,n1971 ,n2092);
    nand g2194(n2232 ,n51[14] ,n1991);
    nand g2195(n1395 ,n42[21] ,n1139);
    nand g2196(n1972 ,n25[24] ,n1693);
    nand g2197(n783 ,n37[0] ,n665);
    nand g2198(n1983 ,n25[13] ,n1693);
    nand g2199(n1373 ,n1127 ,n1126);
    nand g2200(n2207 ,n2049 ,n2156);
    nand g2201(n524 ,n43[0] ,n472);
    nand g2202(n213 ,n46[7] ,n211);
    xnor g2203(n2469 ,n53[14] ,n198);
    nand g2204(n2210 ,n1977 ,n2098);
    not g2205(n962 ,n920);
    xor g2206(n512 ,n41[13] ,n52[13]);
    nand g2207(n1770 ,n1252 ,n1429);
    not g2208(n2136 ,n2006);
    nor g2209(n250 ,n49[3] ,n249);
    not g2210(n317 ,n41[0]);
    nand g2211(n1183 ,n15[3] ,n300);
    nand g2212(n1242 ,n9[15] ,n300);
    or g2213(n1910 ,n1811 ,n1707);
    nand g2214(n1807 ,n1232 ,n1488);
    nand g2215(n571 ,n308 ,n480);
    nor g2216(n99 ,n50[5] ,n98);
    nand g2217(n1273 ,n8[17] ,n299);
    nand g2218(n1981 ,n25[15] ,n1693);
    nand g2219(n735 ,n2451 ,n528);
    nand g2220(n2301 ,n53[1] ,n2259);
    nand g2221(n1969 ,n25[27] ,n1693);
    nand g2222(n1048 ,n13[8] ,n298);
    nand g2223(n267 ,n34[2] ,n266);
    nand g2224(n1088 ,n7[9] ,n296);
    dff g2225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1580), .Q(n29[0]));
    not g2226(n263 ,n34[12]);
    nand g2227(n1959 ,n2506 ,n1700);
    not g2228(n1826 ,n1728);
    nand g2229(n2033 ,n26[12] ,n1695);
    dff g2230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n903), .Q(n46[9]));
    xnor g2231(n2508 ,n50[8] ,n104);
    nand g2232(n1580 ,n304 ,n1329);
    or g2233(n414 ,n38[1] ,n38[3]);
    nand g2234(n2270 ,n1978 ,n2099);
    nand g2235(n2008 ,n1594 ,n1596);
    nand g2236(n817 ,n31[6] ,n666);
    not g2237(n313 ,n41[9]);
    or g2238(n1887 ,n1786 ,n1687);
    nor g2239(n2468 ,n197 ,n199);
    not g2240(n967 ,n926);
    nor g2241(n530 ,n2534 ,n437);
    nand g2242(n580 ,n419 ,n426);
    nand g2243(n2183 ,n51[0] ,n1991);
    nand g2244(n1592 ,n42[24] ,n289);
    not g2245(n275 ,n274);
    nand g2246(n2371 ,n2065 ,n2307);
    nand g2247(n1024 ,n13[12] ,n297);
    nand g2248(n1133 ,n6[28] ,n296);
    nand g2249(n1430 ,n35[2] ,n1141);
    or g2250(n2174 ,n1468 ,n1995);
    not g2251(n1425 ,n1387);
    nand g2252(n879 ,n653 ,n719);
    xnor g2253(n499 ,n41[9] ,n52[9]);
    nand g2254(n2200 ,n2035 ,n2149);
    not g2255(n180 ,n179);
    dff g2256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1843), .Q(n40[11]));
    nand g2257(n2246 ,n1965 ,n2085);
    nor g2258(n459 ,n343 ,n2407);
    nor g2259(n528 ,n2532 ,n470);
    nand g2260(n1976 ,n25[20] ,n1693);
    dff g2261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2184), .Q(n26[27]));
    nand g2262(n708 ,n46[1] ,n529);
    not g2263(n59 ,n22[1]);
    nand g2264(n2237 ,n51[9] ,n1991);
    or g2265(n2516 ,n18[1] ,n18[0]);
    nand g2266(n1049 ,n13[7] ,n848);
    dff g2267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1897), .Q(n41[0]));
    xnor g2268(n2491 ,n51[6] ,n128);
    nand g2269(n2028 ,n1616 ,n1615);
    not g2270(n475 ,n476);
    xnor g2271(n2442 ,n47[5] ,n223);
    nand g2272(n732 ,n2440 ,n526);
    or g2273(n1854 ,n1738 ,n1654);
    or g2274(n1870 ,n1770 ,n1673);
    nand g2275(n2375 ,n2070 ,n2312);
    nor g2276(n2260 ,n761 ,n1919);
    not g2277(n483 ,n482);
    nand g2278(n1255 ,n6[6] ,n295);
    nand g2279(n811 ,n32[3] ,n666);
    not g2280(n129 ,n128);
    nand g2281(n1756 ,n1274 ,n1519);
    nand g2282(n1058 ,n5[30] ,n298);
    nand g2283(n1032 ,n4[15] ,n297);
    nor g2284(n74 ,n47[4] ,n47[3]);
    not g2285(n217 ,n47[6]);
    dff g2286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2364), .Q(n53[1]));
    nand g2287(n109 ,n50[10] ,n108);
    nand g2288(n1324 ,n30[1] ,n1140);
    nand g2289(n2272 ,n1985 ,n2106);
    nand g2290(n800 ,n11[11] ,n293);
    dff g2291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1902), .Q(n40[24]));
    not g2292(n1836 ,n1798);
    or g2293(n477 ,n331 ,n38[3]);
    nand g2294(n838 ,n10[24] ,n293);
    nand g2295(n533 ,n411 ,n472);
    nand g2296(n903 ,n698 ,n740);
    or g2297(n1398 ,n533 ,n1290);
    nor g2298(n2419 ,n2395 ,n2408);
    nand g2299(n1520 ,n1275 ,n1029);
    xnor g2300(n2482 ,n52[12] ,n167);
    nand g2301(n2390 ,n1145 ,n2384);
    not g2302(n222 ,n221);
    dff g2303(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1886), .Q(n41[10]));
    or g2304(n373 ,n319 ,n51[8]);
    not g2305(n668 ,n667);
    nand g2306(n128 ,n51[5] ,n126);
    nand g2307(n1775 ,n1256 ,n1437);
    nand g2308(n1685 ,n889 ,n1534);
    nand g2309(n802 ,n10[7] ,n664);
    not g2310(n90 ,n50[8]);
    nand g2311(n1066 ,n5[23] ,n848);
    nand g2312(n812 ,n32[1] ,n666);
    nand g2313(n2003 ,n1589 ,n1588);
    nand g2314(n1319 ,n511 ,n979);
    not g2315(n237 ,n236);
    nand g2316(n886 ,n724 ,n687);
    nand g2317(n2353 ,n1936 ,n2290);
    nand g2318(n1594 ,n40[23] ,n1397);
    not g2319(n308 ,n2407);
    nor g2320(n113 ,n50[13] ,n112);
    nand g2321(n2261 ,n2127 ,n2117);
    nand g2322(n554 ,n434 ,n363);
    nand g2323(n1625 ,n915 ,n1541);
    xnor g2324(n2463 ,n53[8] ,n188);
    nor g2325(n1293 ,n544 ,n1290);
    nand g2326(n2015 ,n26[20] ,n1695);
    nand g2327(n2070 ,n2475 ,n1696);
    dff g2328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2176), .Q(n40[25]));
    nand g2329(n1644 ,n40[1] ,n291);
    dff g2330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n778), .Q(n38[3]));
    nand g2331(n1640 ,n1093 ,n1412);
    not g2332(n343 ,n45[2]);
    dff g2333(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2376), .Q(n52[4]));
    nand g2334(n2022 ,n1608 ,n1609);
    nand g2335(n889 ,n16[11] ,n293);
    nor g2336(n82 ,n81 ,n79);
    nand g2337(n745 ,n2431 ,n530);
    nand g2338(n1641 ,n42[3] ,n289);
    nor g2339(n385 ,n313 ,n53[9]);
    nor g2340(n169 ,n52[13] ,n168);
    nand g2341(n1662 ,n842 ,n1411);
    nand g2342(n2304 ,n52[13] ,n2260);
    nand g2343(n565 ,n443 ,n367);
    nand g2344(n1583 ,n859 ,n1324);
    not g2345(n413 ,n412);
    not g2346(n851 ,n850);
    nand g2347(n790 ,n39[0] ,n665);
    not g2348(n2396 ,n18[0]);
    nand g2349(n1288 ,n6[25] ,n847);
    or g2350(n1879 ,n1780 ,n1681);
    not g2351(n1154 ,n1107);
    nand g2352(n1366 ,n1116 ,n1009);
    or g2353(n2175 ,n1477 ,n1998);
    dff g2354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2374), .Q(n52[6]));
    nor g2355(n2483 ,n169 ,n171);
    nand g2356(n1077 ,n7[13] ,n847);
    nor g2357(n1881 ,n524 ,n1704);
    nand g2358(n683 ,n47[3] ,n587);
    nor g2359(n2509 ,n106 ,n108);
    nand g2360(n1793 ,n1187 ,n1314);
    nand g2361(n1386 ,n42[25] ,n1139);
    nand g2362(n1389 ,n42[24] ,n1139);
    or g2363(n1862 ,n1753 ,n1662);
    not g2364(n1536 ,n1454);
    not g2365(n1404 ,n1292);
    nor g2366(n2440 ,n220 ,n222);
    nand g2367(n1780 ,n1161 ,n1301);
    xnor g2368(n2459 ,n53[4] ,n181);
    nand g2369(n2201 ,n2036 ,n2150);
    not g2370(n292 ,n306);
    nand g2371(n61 ,n2416 ,n59);
    nor g2372(n1399 ,n301 ,n1143);
    nand g2373(n1470 ,n931 ,n1060);
    nand g2374(n1250 ,n8[0] ,n299);
    nand g2375(n2068 ,n2477 ,n1696);
    nand g2376(n447 ,n52[4] ,n316);
    dff g2377(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n618), .Q(n33[4]));
    nand g2378(n2222 ,n50[5] ,n1992);
    nand g2379(n1014 ,n4[30] ,n298);
    nor g2380(n534 ,n440 ,n415);
    nand g2381(n2302 ,n52[15] ,n2260);
    nand g2382(n1188 ,n6[4] ,n295);
    dff g2383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2357), .Q(n53[9]));
    nand g2384(n2284 ,n53[0] ,n2259);
    or g2385(n1843 ,n1724 ,n1601);
    nand g2386(n1677 ,n1188 ,n1527);
    nor g2387(n467 ,n319 ,n50[8]);
    nor g2388(n226 ,n217 ,n225);
    dff g2389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2274), .Q(n25[13]));
    nand g2390(n1202 ,n9[30] ,n300);
    xnor g2391(n2452 ,n46[6] ,n210);
    nand g2392(n418 ,n50[15] ,n320);
    nand g2393(n1064 ,n13[14] ,n298);
    not g2394(n108 ,n107);
    nand g2395(n474 ,n35[0] ,n2532);
    nor g2396(n1704 ,n540 ,n291);
    nand g2397(n919 ,n689 ,n635);
    nor g2398(n219 ,n216 ,n218);
    dff g2399(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2375), .Q(n52[5]));
    nand g2400(n276 ,n34[7] ,n275);
    nand g2401(n1098 ,n7[5] ,n295);
    nand g2402(n97 ,n50[3] ,n96);
    nand g2403(n1624 ,n805 ,n1410);
    nand g2404(n359 ,n50[0] ,n317);
    nand g2405(n1590 ,n40[25] ,n291);
    not g2406(n305 ,n849);
    dff g2407(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n882), .Q(n49[1]));
    nor g2408(n974 ,n524 ,n854);
    nand g2409(n1454 ,n1169 ,n1047);
    nand g2410(n2314 ,n52[3] ,n2260);
    nand g2411(n1312 ,n41[4] ,n292);
    not g2412(n1544 ,n1462);
    nand g2413(n685 ,n46[4] ,n529);
    nand g2414(n1723 ,n1079 ,n1332);
    nand g2415(n1023 ,n13[11] ,n297);
    nand g2416(n1733 ,n1115 ,n1365);
    nand g2417(n658 ,n49[4] ,n588);
    dff g2418(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1205), .Q(n34[5]));
    nand g2419(n703 ,n2434 ,n530);
    nand g2420(n1464 ,n40[31] ,n292);
    not g2421(n1528 ,n1444);
    nand g2422(n1955 ,n2509 ,n1700);
    nand g2423(n1384 ,n42[26] ,n1139);
    nand g2424(n2209 ,n2052 ,n2158);
    nor g2425(n1567 ,n670 ,n1319);
    nand g2426(n1267 ,n8[14] ,n849);
    nand g2427(n2391 ,n2387 ,n2389);
    nor g2428(n72 ,n71 ,n69);
    not g2429(n145 ,n52[4]);
    nor g2430(n2490 ,n127 ,n129);
    nand g2431(n1450 ,n1178 ,n1046);
    nand g2432(n1337 ,n803 ,n999);
    nand g2433(n2196 ,n2027 ,n2145);
    nand g2434(n2331 ,n2084 ,n2245);
    nand g2435(n1651 ,n1113 ,n1416);
    or g2436(n1897 ,n1795 ,n1823);
    nand g2437(n1161 ,n14[15] ,n847);
    nor g2438(n2534 ,n80 ,n83);
    nand g2439(n2291 ,n53[11] ,n2259);
    nand g2440(n253 ,n49[4] ,n252);
    nand g2441(n1937 ,n2466 ,n1698);
    nand g2442(n956 ,n708 ,n710);
    nand g2443(n727 ,n48[0] ,n527);
    nor g2444(n407 ,n321 ,n51[10]);
    nand g2445(n729 ,n2445 ,n526);
    or g2446(n1873 ,n1769 ,n1676);
    nor g2447(n2513 ,n113 ,n115);
    nand g2448(n1953 ,n2511 ,n1700);
    nor g2449(n994 ,n548 ,n762);
    dff g2450(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2264), .Q(n25[3]));
    dff g2451(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1845), .Q(n40[9]));
    nand g2452(n1646 ,n42[0] ,n289);
    nand g2453(n682 ,n2528 ,n523);
    nand g2454(n1171 ,n15[8] ,n299);
    dff g2455(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n798), .Q(n46[4]));
    nor g2456(n234 ,n231 ,n233);
    nand g2457(n116 ,n50[14] ,n115);
    dff g2458(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n956), .Q(n46[1]));
    nand g2459(n139 ,n51[11] ,n138);
    nand g2460(n1935 ,n302 ,n1768);
    nand g2461(n2266 ,n1993 ,n2112);
    not g2462(n2143 ,n2022);
    nor g2463(n397 ,n315 ,n53[13]);
    nand g2464(n846 ,n647 ,n607);
    nand g2465(n921 ,n686 ,n633);
    nor g2466(n1206 ,n2407 ,n968);
    not g2467(n187 ,n186);
    dff g2468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2322), .Q(n51[11]));
    nand g2469(n1582 ,n859 ,n1322);
    nor g2470(n63 ,n2415 ,n62);
    nand g2471(n704 ,n2432 ,n530);
    nand g2472(n2311 ,n52[6] ,n2260);
    nand g2473(n1321 ,n44[1] ,n1139);
    nand g2474(n689 ,n34[15] ,n524);
    dff g2475(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1858), .Q(n42[26]));
    nand g2476(n762 ,n506 ,n614);
    nand g2477(n2317 ,n2074 ,n2231);
    not g2478(n214 ,n213);
    nand g2479(n2227 ,n2120 ,n2161);
    nand g2480(n1028 ,n4[19] ,n297);
    nand g2481(n697 ,n46[3] ,n529);
    dff g2482(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n990), .Q(n38[2]));
    nand g2483(n933 ,n11[27] ,n293);
    nand g2484(n1080 ,n9[11] ,n300);
    nand g2485(n1608 ,n40[17] ,n291);
    nand g2486(n1286 ,n6[24] ,n295);
    dff g2487(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1852), .Q(n40[0]));
    nand g2488(n177 ,n53[1] ,n53[0]);
    nand g2489(n1046 ,n13[13] ,n848);
    nand g2490(n876 ,n16[15] ,n293);
    nand g2491(n2368 ,n2063 ,n2305);
    nand g2492(n1375 ,n832 ,n1014);
    nand g2493(n1741 ,n1133 ,n1380);
    or g2494(n856 ,n414 ,n674);
    dff g2495(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1927), .Q(n36[3]));
    nor g2496(n2178 ,n2407 ,n2118);
    dff g2497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1348), .Q(n32[3]));
    nand g2498(n1276 ,n6[19] ,n295);
    nand g2499(n2062 ,n2483 ,n1696);
    nand g2500(n1689 ,n907 ,n1538);
    dff g2501(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1895), .Q(n41[2]));
    nor g2502(n540 ,n43[0] ,n413);
    nand g2503(n861 ,n537 ,n667);
    nand g2504(n2316 ,n52[1] ,n2260);
    nand g2505(n820 ,n31[4] ,n666);
    nand g2506(n421 ,n52[7] ,n327);
    nor g2507(n1700 ,n677 ,n1398);
    nor g2508(n612 ,n590 ,n535);
    nand g2509(n2079 ,n2494 ,n1701);
    dff g2510(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2278), .Q(n25[17]));
    nand g2511(n756 ,n49[9] ,n588);
    nand g2512(n1068 ,n5[21] ,n848);
    nor g2513(n777 ,n450 ,n631);
    nand g2514(n935 ,n11[26] ,n293);
    nand g2515(n1344 ,n809 ,n1003);
    nand g2516(n2228 ,n2122 ,n2162);
    nand g2517(n1785 ,n1168 ,n1306);
    nand g2518(n1602 ,n42[20] ,n289);
    nand g2519(n2119 ,n1711 ,n1710);
    not g2520(n300 ,n305);
    not g2521(n297 ,n304);
    nand g2522(n996 ,n5[11] ,n298);
    nor g2523(n460 ,n342 ,n2407);
    nand g2524(n2069 ,n2476 ,n1696);
    nand g2525(n2042 ,n1632 ,n1631);
    nand g2526(n955 ,n10[15] ,n664);
    nor g2527(n1403 ,n571 ,n977);
    nand g2528(n2101 ,n12[16] ,n1694);
    nand g2529(n1329 ,n29[0] ,n1142);
    nand g2530(n1998 ,n1217 ,n1837);
    nor g2531(n2479 ,n162 ,n164);
    nand g2532(n647 ,n47[0] ,n587);
    nand g2533(n458 ,n52[1] ,n328);
    nand g2534(n142 ,n51[13] ,n140);
    nand g2535(n2263 ,n2129 ,n2115);
    nand g2536(n479 ,n43[2] ,n329);
    nand g2537(n1987 ,n25[9] ,n1693);
    nor g2538(n65 ,n64 ,n2413);
    nand g2539(n1504 ,n29[2] ,n1141);
    nand g2540(n1101 ,n812 ,n782);
    nand g2541(n920 ,n750 ,n634);
    nand g2542(n419 ,n50[1] ,n328);
    dff g2543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1841), .Q(n40[12]));
    nand g2544(n815 ,n32[0] ,n666);
    nand g2545(n1122 ,n9[0] ,n849);
    nand g2546(n449 ,n52[5] ,n314);
    nand g2547(n1457 ,n1177 ,n1021);
    dff g2548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2337), .Q(n50[10]));
    nand g2549(n990 ,n621 ,n305);
    nand g2550(n796 ,n738 ,n605);
    nand g2551(n721 ,n2421 ,n525);
    nand g2552(n1462 ,n1191 ,n1056);
    not g2553(n2137 ,n2008);
    nand g2554(n1788 ,n1174 ,n1309);
    xnor g2555(n2423 ,n49[4] ,n251);
    nand g2556(n1971 ,n25[25] ,n1693);
    nand g2557(n1921 ,n1117 ,n1827);
    nand g2558(n2096 ,n12[21] ,n1694);
    nand g2559(n999 ,n4[2] ,n297);
    nand g2560(n2240 ,n51[6] ,n1991);
    not g2561(n2148 ,n2032);
    nand g2562(n737 ,n2448 ,n528);
    nand g2563(n251 ,n49[3] ,n249);
    nand g2564(n759 ,n366 ,n597);
    nand g2565(n794 ,n39[2] ,n665);
    nand g2566(n2336 ,n1952 ,n2215);
    dff g2567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n879), .Q(n49[6]));
    not g2568(n1546 ,n1465);
    xnor g2569(n2476 ,n52[6] ,n156);
    nor g2570(n651 ,n2407 ,n559);
    dff g2571(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1352), .Q(n32[0]));
    not g2572(n1158 ,n1114);
    nand g2573(n1050 ,n13[6] ,n848);
    not g2574(n254 ,n253);
    nor g2575(n406 ,n318 ,n51[14]);
    not g2576(n1426 ,n1394);
    nand g2577(n1069 ,n5[20] ,n297);
    nand g2578(n1117 ,n19[1] ,n296);
    nand g2579(n556 ,n456 ,n468);
    nand g2580(n1926 ,n839 ,n1831);
    nand g2581(n1950 ,n2514 ,n1700);
    nand g2582(n1471 ,n40[28] ,n1139);
    not g2583(n1523 ,n1432);
    nand g2584(n1463 ,n865 ,n1057);
    nand g2585(n953 ,n10[13] ,n293);
    nand g2586(n1172 ,n14[8] ,n295);
    nor g2587(n69 ,n46[4] ,n46[3]);
    nand g2588(n743 ,n2429 ,n530);
    dff g2589(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2257), .Q(n25[20]));
    nand g2590(n1581 ,n304 ,n1327);
    nand g2591(n2012 ,n1599 ,n1600);
    not g2592(n853 ,n852);
    nand g2593(n1670 ,n1260 ,n1561);
    nand g2594(n1084 ,n14[14] ,n295);
    dff g2595(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1900), .Q(n40[28]));
    dff g2596(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2266), .Q(n25[5]));
    xnor g2597(n2512 ,n50[12] ,n111);
    not g2598(n289 ,n290);
    nand g2599(n2251 ,n1970 ,n2091);
    nand g2600(n1025 ,n4[22] ,n298);
    or g2601(n350 ,n36[0] ,n36[1]);
    or g2602(n1912 ,n1812 ,n1719);
    nand g2603(n1966 ,n25[30] ,n1693);
    not g2604(n1551 ,n1484);
    nand g2605(n893 ,n16[10] ,n293);
    nand g2606(n2065 ,n2480 ,n1696);
    nand g2607(n1325 ,n30[0] ,n1142);
    nor g2608(n141 ,n51[13] ,n140);
    nand g2609(n1017 ,n4[27] ,n298);
    nand g2610(n76 ,n47[9] ,n47[8]);
    nand g2611(n1794 ,n1190 ,n1315);
    not g2612(n1831 ,n1750);
    nand g2613(n2191 ,n2015 ,n2140);
    not g2614(n2402 ,n2410);
    not g2615(n298 ,n304);
    nand g2616(n1778 ,n1159 ,n1445);
    not g2617(n336 ,n53[3]);
    nor g2618(n623 ,n2407 ,n562);
    nand g2619(n1435 ,n1253 ,n1039);
    xnor g2620(n2425 ,n49[6] ,n255);
    nand g2621(n1767 ,n862 ,n1503);
    not g2622(n332 ,n51[0]);
    or g2623(n1858 ,n1743 ,n1658);
    nand g2624(n947 ,n11[15] ,n293);
    nand g2625(n1932 ,n1144 ,n1761);
    xnor g2626(n515 ,n41[13] ,n50[13]);
    nand g2627(n2220 ,n50[7] ,n1992);
    nand g2628(n1712 ,n949 ,n1539);
    nand g2629(n748 ,n34[11] ,n524);
    nand g2630(n1736 ,n1120 ,n1370);
    nand g2631(n123 ,n51[2] ,n122);
    nor g2632(n2460 ,n183 ,n185);
    not g2633(n523 ,n524);
    nor g2634(n1694 ,n44[1] ,n307);
    not g2635(n273 ,n272);
    not g2636(n1830 ,n1748);
    nand g2637(n1007 ,n5[3] ,n297);
    nand g2638(n578 ,n457 ,n433);
    dff g2639(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2201), .Q(n26[10]));
    not g2640(n2406 ,n2416);
    nand g2641(n184 ,n53[5] ,n182);
    or g2642(n1878 ,n1777 ,n1678);
    dff g2643(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n894), .Q(n48[1]));
    nor g2644(n1573 ,n774 ,n1294);
    nand g2645(n1626 ,n40[10] ,n291);
    nand g2646(n1616 ,n40[14] ,n1397);
    or g2647(n1889 ,n1788 ,n1689);
    nor g2648(n264 ,n34[1] ,n34[0]);
    dff g2649(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1905), .Q(n40[20]));
    nand g2650(n1162 ,n14[13] ,n847);
    nand g2651(n435 ,n53[10] ,n321);
    nand g2652(n1818 ,n1222 ,n1549);
    nand g2653(n1353 ,n40[4] ,n1139);
    nand g2654(n833 ,n10[29] ,n294);
    or g2655(n598 ,n569 ,n554);
    nand g2656(n1960 ,n2505 ,n1700);
    nand g2657(n691 ,n2452 ,n528);
    nand g2658(n808 ,n11[7] ,n293);
    nand g2659(n1757 ,n1272 ,n1517);
    or g2660(n1572 ,n301 ,n1401);
    nand g2661(n1635 ,n42[5] ,n289);
    nand g2662(n734 ,n2454 ,n528);
    nand g2663(n1474 ,n40[27] ,n1139);
    or g2664(n1295 ,n677 ,n981);
    dff g2665(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1201), .Q(n34[8]));
    nor g2666(n1357 ,n2407 ,n1153);
    not g2667(n2151 ,n2038);
    nand g2668(n1771 ,n870 ,n1446);
    dff g2669(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1865), .Q(n42[17]));
    or g2670(n677 ,n38[2] ,n589);
    nor g2671(n975 ,n593 ,n857);
    nor g2672(n2498 ,n141 ,n143);
    nand g2673(n1268 ,n6[15] ,n847);
    nand g2674(n446 ,n52[14] ,n318);
    nand g2675(n179 ,n53[2] ,n178);
    nand g2676(n563 ,n466 ,n375);
    nand g2677(n1747 ,n1286 ,n1389);
    xnor g2678(n2487 ,n51[2] ,n121);
    nand g2679(n269 ,n34[3] ,n268);
    nor g2680(n2535 ,n85 ,n88);
    dff g2681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1207), .Q(n34[2]));
    nor g2682(n771 ,n43[2] ,n673);
    nand g2683(n2329 ,n2082 ,n2243);
    nand g2684(n858 ,n637 ,n611);
    dff g2685(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2185), .Q(n26[26]));
    nand g2686(n2363 ,n2073 ,n2315);
    nand g2687(n700 ,n478 ,n531);
    nand g2688(n2081 ,n2491 ,n1701);
    nand g2689(n2208 ,n2051 ,n2157);
    nand g2690(n279 ,n34[9] ,n277);
    nor g2691(n1349 ,n2407 ,n1148);
    nand g2692(n1945 ,n2456 ,n1698);
    nor g2693(n2380 ,n2349 ,n2280);
    nand g2694(n917 ,n746 ,n680);
    not g2695(n330 ,n38[2]);
    nand g2696(n863 ,n658 ,n714);
    nand g2697(n766 ,n509 ,n594);
    nand g2698(n575 ,n447 ,n421);
    nand g2699(n2059 ,n2471 ,n1696);
    nand g2700(n1245 ,n28 ,n854);
    dff g2701(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n877), .Q(n47[8]));
    not g2702(n216 ,n47[2]);
    nand g2703(n86 ,n49[9] ,n49[8]);
    nand g2704(n829 ,n11[0] ,n294);
    not g2705(n1563 ,n1514);
    not g2706(n1534 ,n1452);
    nand g2707(n1638 ,n40[4] ,n1397);
    nor g2708(n620 ,n312 ,n589);
    xnor g2709(n2521 ,n34[11] ,n281);
    or g2710(n349 ,n39[2] ,n39[3]);
    nand g2711(n1769 ,n866 ,n1428);
    nor g2712(n368 ,n314 ,n50[5]);
    xnor g2713(n2502 ,n50[2] ,n93);
    nand g2714(n2046 ,n1636 ,n1635);
    nand g2715(n1654 ,n1128 ,n1419);
    or g2716(n371 ,n327 ,n52[7]);
    nand g2717(n2225 ,n50[2] ,n1992);
    nand g2718(n2249 ,n1968 ,n2089);
    nand g2719(n867 ,n10[9] ,n294);
    nand g2720(n2279 ,n1987 ,n2108);
    dff g2721(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1884), .Q(n41[12]));
    dff g2722(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1196), .Q(n34[11]));
    nand g2723(n1045 ,n4[5] ,n298);
    nand g2724(n431 ,n51[10] ,n321);
    nand g2725(n572 ,n308 ,n474);
    nand g2726(n2089 ,n12[28] ,n1694);
    dff g2727(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2350), .Q(n53[15]));
    nand g2728(n2071 ,n2474 ,n1696);
    nand g2729(n2026 ,n1612 ,n1614);
    dff g2730(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n911), .Q(n49[3]));
    dff g2731(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2333), .Q(n50[14]));
    nand g2732(n1071 ,n5[18] ,n297);
    not g2733(n1835 ,n1779);
    nand g2734(n2276 ,n1981 ,n2102);
    nor g2735(n492 ,n388 ,n395);
    or g2736(n356 ,n2[3] ,n2[2]);
    nand g2737(n557 ,n359 ,n462);
    not g2738(n1554 ,n1490);
    nand g2739(n258 ,n49[7] ,n256);
    nand g2740(n2346 ,n52[4] ,n2260);
    not g2741(n2135 ,n2004);
    nand g2742(n2117 ,n12[0] ,n1694);
    nand g2743(n2347 ,n1874 ,n2284);
    nand g2744(n1790 ,n1179 ,n1311);
    nand g2745(n2057 ,n1648 ,n1646);
    or g2746(n1880 ,n1781 ,n1682);
    or g2747(n498 ,n389 ,n377);
    nand g2748(n1305 ,n41[11] ,n292);
    dff g2749(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2392), .Q(n45[1]));
    nand g2750(n2108 ,n12[9] ,n1694);
    dff g2751(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1873), .Q(n42[6]));
    nor g2752(n155 ,n52[5] ,n154);
    nand g2753(n1247 ,n7[14] ,n295);
    nor g2754(n1289 ,n2407 ,n959);
    nand g2755(n1116 ,n9[1] ,n299);
    nand g2756(n1746 ,n861 ,n1388);
    nand g2757(n2039 ,n26[9] ,n1695);
    dff g2758(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2365), .Q(n52[15]));
    nand g2759(n433 ,n53[15] ,n320);
    or g2760(n1847 ,n1729 ,n1640);
    not g2761(n302 ,n664);
    nand g2762(n1722 ,n1077 ,n1330);
    nand g2763(n713 ,n48[8] ,n527);
    not g2764(n229 ,n228);
    dff g2765(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2195), .Q(n26[16]));
    nand g2766(n1199 ,n7[31] ,n295);
    buf g2767(n32[6], 1'b0);
    not g2768(n1559 ,n1500);
    nand g2769(n869 ,n645 ,n709);
    or g2770(n1874 ,n53[0] ,n1697);
    nand g2771(n1967 ,n25[29] ,n1693);
    nand g2772(n884 ,n16[12] ,n664);
    not g2773(n1531 ,n1449);
    nand g2774(n714 ,n2423 ,n525);
    nand g2775(n813 ,n32[2] ,n666);
    dff g2776(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2279), .Q(n25[9]));
    dff g2777(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n460), .Q(n43[0]));
    nand g2778(n951 ,n707 ,n737);
    dff g2779(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2207), .Q(n26[4]));
    nand g2780(n160 ,n52[7] ,n159);
    nand g2781(n2394 ,n2386 ,n2393);
    nand g2782(n1211 ,n8[10] ,n299);
    dff g2783(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2330), .Q(n51[2]));
    nand g2784(n1275 ,n8[18] ,n299);
    nand g2785(n1356 ,n819 ,n1007);
    nand g2786(n1181 ,n14[4] ,n847);
    nand g2787(n2029 ,n26[14] ,n1695);
    nand g2788(n1119 ,n21[1] ,n299);
    nand g2789(n720 ,n2422 ,n525);
    nand g2790(n1075 ,n4[9] ,n297);
    nand g2791(n786 ,n36[1] ,n665);
    not g2792(n673 ,n672);
    nand g2793(n1249 ,n6[5] ,n295);
    nand g2794(n1999 ,n1237 ,n1839);
    nand g2795(n1934 ,n302 ,n1764);
    nand g2796(n1916 ,n516 ,n1573);
    dff g2797(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1906), .Q(n40[21]));
    nand g2798(n1940 ,n2460 ,n1698);
    nand g2799(n1666 ,n1271 ,n1564);
    dff g2800(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1195), .Q(n34[12]));
    nand g2801(n2041 ,n26[8] ,n1695);
    nand g2802(n2358 ,n1942 ,n2294);
    nand g2803(n1943 ,n2457 ,n1698);
    nand g2804(n1974 ,n25[22] ,n1693);
    nor g2805(n278 ,n34[9] ,n277);
    nand g2806(n1986 ,n25[10] ,n1693);
    dff g2807(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2367), .Q(n52[13]));
endmodule
