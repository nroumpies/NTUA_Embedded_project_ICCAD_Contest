module top (n0, n1, n2, n3, n4, n5, n6, n7);
    input n0, n1, n2, n3;
    input [15:0] n4;
    output [15:0] n5;
    output n6, n7;
    wire n0, n1, n2, n3;
    wire [15:0] n4;
    wire [15:0] n5;
    wire n6, n7;
    wire [15:0] n8;
    wire [15:0] n9;
    wire [15:0] n10;
    wire [15:0] n11;
    wire [15:0] n12;
    wire [15:0] n13;
    wire [15:0] n14;
    wire [15:0] n15;
    wire [15:0] n16;
    wire [15:0] n17;
    wire [15:0] n18;
    wire [15:0] n19;
    wire [15:0] n20;
    wire [15:0] n21;
    wire [15:0] n22;
    wire [15:0] n23;
    wire [15:0] n24;
    wire [15:0] n25;
    wire [15:0] n26;
    wire [15:0] n27;
    wire [15:0] n28;
    wire [15:0] n29;
    wire [15:0] n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
    wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
    wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
    wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
    wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
    wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
    wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
    wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
    wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
    wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
    wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
    wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
    wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
    wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
    wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
    wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
    wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
    wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
    wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
    wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
    wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
    wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
    wire n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742;
    wire n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750;
    wire n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758;
    wire n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766;
    wire n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774;
    wire n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782;
    wire n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790;
    wire n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798;
    wire n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806;
    wire n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814;
    wire n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822;
    wire n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
    wire n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838;
    wire n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846;
    wire n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854;
    wire n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
    wire n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870;
    wire n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878;
    wire n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886;
    wire n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894;
    wire n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902;
    wire n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910;
    wire n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918;
    wire n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
    wire n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934;
    wire n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
    wire n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950;
    wire n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958;
    wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
    wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974;
    wire n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982;
    wire n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990;
    wire n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998;
    wire n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
    wire n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014;
    wire n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022;
    wire n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;
    wire n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038;
    wire n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046;
    wire n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054;
    wire n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062;
    wire n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070;
    wire n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078;
    wire n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086;
    wire n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094;
    wire n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102;
    wire n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110;
    wire n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118;
    wire n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126;
    wire n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134;
    wire n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142;
    wire n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150;
    wire n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158;
    wire n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166;
    wire n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174;
    wire n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182;
    wire n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190;
    wire n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198;
    wire n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206;
    wire n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214;
    wire n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222;
    wire n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230;
    wire n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238;
    wire n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246;
    wire n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254;
    wire n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262;
    wire n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270;
    wire n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278;
    wire n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286;
    wire n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294;
    wire n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302;
    wire n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310;
    wire n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318;
    wire n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326;
    wire n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334;
    wire n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342;
    wire n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350;
    wire n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358;
    wire n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366;
    wire n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374;
    wire n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382;
    wire n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390;
    wire n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398;
    wire n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406;
    wire n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414;
    wire n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422;
    wire n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430;
    wire n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438;
    wire n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446;
    wire n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454;
    wire n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462;
    wire n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470;
    wire n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478;
    wire n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486;
    wire n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494;
    wire n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502;
    wire n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510;
    wire n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518;
    wire n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526;
    wire n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534;
    wire n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542;
    wire n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550;
    wire n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558;
    wire n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566;
    wire n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574;
    wire n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582;
    wire n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590;
    wire n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598;
    wire n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606;
    wire n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614;
    wire n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622;
    wire n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630;
    wire n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638;
    wire n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646;
    wire n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654;
    wire n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662;
    wire n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670;
    wire n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678;
    wire n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686;
    wire n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694;
    wire n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702;
    wire n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710;
    wire n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718;
    wire n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726;
    wire n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734;
    wire n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742;
    wire n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750;
    wire n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758;
    wire n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766;
    wire n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774;
    wire n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782;
    wire n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790;
    wire n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798;
    wire n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806;
    wire n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814;
    wire n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822;
    wire n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830;
    wire n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838;
    wire n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846;
    wire n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854;
    wire n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862;
    wire n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870;
    wire n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878;
    wire n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886;
    wire n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894;
    wire n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902;
    wire n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910;
    wire n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918;
    wire n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926;
    wire n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934;
    wire n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942;
    wire n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950;
    wire n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958;
    wire n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966;
    wire n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974;
    wire n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982;
    wire n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990;
    wire n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998;
    wire n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006;
    wire n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014;
    wire n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022;
    wire n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030;
    wire n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038;
    wire n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046;
    wire n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054;
    wire n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062;
    wire n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070;
    wire n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078;
    wire n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086;
    wire n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094;
    wire n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102;
    wire n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110;
    wire n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118;
    wire n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126;
    wire n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134;
    wire n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142;
    wire n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150;
    wire n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158;
    wire n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166;
    wire n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174;
    wire n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182;
    wire n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190;
    wire n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198;
    wire n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206;
    wire n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214;
    wire n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222;
    wire n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230;
    wire n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238;
    wire n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246;
    wire n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254;
    wire n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262;
    wire n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270;
    wire n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278;
    wire n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286;
    wire n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294;
    wire n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302;
    wire n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310;
    wire n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318;
    wire n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326;
    wire n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334;
    wire n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342;
    wire n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350;
    wire n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358;
    wire n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366;
    wire n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374;
    wire n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382;
    wire n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390;
    wire n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398;
    wire n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406;
    wire n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414;
    wire n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422;
    wire n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430;
    wire n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438;
    wire n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446;
    wire n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454;
    wire n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462;
    wire n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470;
    wire n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478;
    wire n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486;
    wire n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494;
    wire n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502;
    wire n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510;
    wire n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518;
    wire n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526;
    wire n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534;
    wire n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542;
    wire n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550;
    wire n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558;
    wire n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566;
    wire n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574;
    wire n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582;
    wire n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590;
    wire n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598;
    wire n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606;
    wire n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614;
    wire n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622;
    wire n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630;
    wire n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638;
    wire n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646;
    wire n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654;
    wire n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662;
    wire n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670;
    wire n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678;
    wire n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686;
    wire n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694;
    wire n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702;
    wire n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710;
    wire n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718;
    wire n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726;
    wire n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734;
    wire n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742;
    wire n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750;
    wire n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758;
    wire n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766;
    wire n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774;
    wire n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782;
    wire n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790;
    wire n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798;
    wire n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806;
    wire n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814;
    wire n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822;
    wire n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830;
    wire n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838;
    wire n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846;
    wire n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854;
    wire n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862;
    wire n3863, n3864, n3865, n3866, n3867, n3868, n3869;
    nand g0(n634 ,n180 ,n445);
    xnor g1(n2104 ,n1945 ,n2039);
    dff g2(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1426), .Q(n12[13]));
    nand g3(n1048 ,n22[15] ,n463);
    nand g4(n1167 ,n22[6] ,n451);
    not g5(n2066 ,n2067);
    dff g6(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1398), .Q(n12[12]));
    nand g7(n3280 ,n3184 ,n3247);
    nand g8(n2032 ,n3850 ,n1986);
    nand g9(n3523 ,n3461 ,n3498);
    nor g10(n2529 ,n2463 ,n2497);
    nand g11(n1722 ,n1680 ,n1679);
    xor g12(n2985 ,n2761 ,n2715);
    nand g13(n990 ,n19[13] ,n482);
    nor g14(n471 ,n213 ,n412);
    nand g15(n1102 ,n15[14] ,n443);
    nand g16(n2193 ,n2070 ,n2129);
    xnor g17(n3328 ,n3224 ,n3157);
    nand g18(n1223 ,n14[12] ,n466);
    dff g19(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1468), .Q(n10[11]));
    nand g20(n2023 ,n3852 ,n1987);
    nand g21(n3096 ,n2888 ,n3025);
    nor g22(n1315 ,n788 ,n771);
    nand g23(n1119 ,n15[4] ,n443);
    nor g24(n493 ,n211 ,n406);
    nor g25(n2166 ,n2105 ,n2148);
    not g26(n77 ,n76);
    xnor g27(n3231 ,n3156 ,n3152);
    xnor g28(n2643 ,n2609 ,n2567);
    nand g29(n1928 ,n3853 ,n1922);
    nand g30(n1585 ,n871 ,n1053);
    nand g31(n549 ,n183 ,n449);
    nand g32(n338 ,n26[7] ,n247);
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1555), .Q(n18[11]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n229), .Q(n27[3]));
    nand g35(n3403 ,n3331 ,n3365);
    nand g36(n3141 ,n3054 ,n3055);
    nand g37(n3386 ,n3249 ,n3343);
    nor g38(n1285 ,n779 ,n798);
    nand g39(n1165 ,n13[10] ,n501);
    nand g40(n426 ,n315 ,n381);
    nand g41(n2033 ,n3856 ,n1985);
    nor g42(n2401 ,n2356 ,n2400);
    nand g43(n567 ,n204 ,n485);
    nand g44(n1877 ,n41 ,n40);
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1364), .Q(n21[8]));
    nand g46(n1160 ,n22[9] ,n451);
    nand g47(n590 ,n187 ,n453);
    xnor g48(n3527 ,n3481 ,n3493);
    nor g49(n347 ,n322 ,n318);
    not g50(n108 ,n27[6]);
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1533), .Q(n22[4]));
    nand g52(n1144 ,n8[3] ,n489);
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1520), .Q(n14[1]));
    nand g54(n3402 ,n3296 ,n3369);
    nand g55(n304 ,n132 ,n241);
    nand g56(n758 ,n182 ,n488);
    nand g57(n39 ,n26[5] ,n36);
    nor g58(n3615 ,n3843 ,n3827);
    nand g59(n3770 ,n3687 ,n3702);
    nand g60(n1163 ,n9[11] ,n459);
    nand g61(n922 ,n13[8] ,n448);
    nor g62(n2432 ,n2407 ,n2421);
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1462), .Q(n10[13]));
    nand g64(n1183 ,n9[6] ,n459);
    xor g65(n3811 ,n28[1] ,n27[1]);
    nor g66(n3818 ,n2953 ,n2900);
    or g67(n3469 ,n3410 ,n3445);
    nand g68(n1376 ,n939 ,n568);
    xnor g69(n2578 ,n2531 ,n2447);
    xnor g70(n1910 ,n27[6] ,n27[5]);
    or g71(n1789 ,n359 ,n1771);
    xnor g72(n3369 ,n3265 ,n3271);
    nand g73(n1339 ,n1274 ,n524);
    nand g74(n1207 ,n13[13] ,n501);
    nor g75(n2566 ,n2506 ,n2516);
    nand g76(n1093 ,n16[3] ,n444);
    nand g77(n2771 ,n27[6] ,n4[1]);
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1415), .Q(n19[5]));
    nand g79(n2003 ,n3855 ,n1963);
    not g80(n2595 ,n2594);
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1476), .Q(n15[9]));
    or g82(n1859 ,n1798 ,n1854);
    xnor g83(n2261 ,n2204 ,n1896);
    nand g84(n2025 ,n3851 ,n1986);
    nand g85(n1196 ,n22[12] ,n463);
    nand g86(n374 ,n276 ,n307);
    nor g87(n764 ,n10[3] ,n503);
    nor g88(n1884 ,n92 ,n90);
    nand g89(n3021 ,n2851 ,n2909);
    xnor g90(n2124 ,n2064 ,n1955);
    nand g91(n2745 ,n27[6] ,n4[5]);
    xnor g92(n2254 ,n2202 ,n2122);
    nand g93(n1003 ,n20[2] ,n452);
    nand g94(n1328 ,n865 ,n510);
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n382), .Q(n24[2]));
    nand g96(n1392 ,n959 ,n587);
    nand g97(n1076 ,n16[9] ,n444);
    nand g98(n942 ,n20[15] ,n452);
    xnor g99(n2126 ,n2058 ,n1957);
    nand g100(n1435 ,n1039 ,n668);
    nand g101(n636 ,n182 ,n457);
    xnor g102(n2323 ,n2252 ,n2285);
    xnor g103(n3224 ,n3106 ,n3108);
    nand g104(n419 ,n5[2] ,n359);
    nand g105(n716 ,n181 ,n488);
    not g106(n2406 ,n5[3]);
    xnor g107(n3242 ,n3133 ,n3094);
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1380), .Q(n20[13]));
    not g109(n2770 ,n2769);
    or g110(n1814 ,n29[2] ,n1784);
    nand g111(n1120 ,n15[3] ,n443);
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n430), .Q(n26[13]));
    nand g113(n672 ,n186 ,n440);
    nand g114(n1577 ,n1032 ,n1218);
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1384), .Q(n20[11]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1407), .Q(n19[10]));
    xor g117(n3436 ,n3399 ,n3414);
    nand g118(n2188 ,n2126 ,n2124);
    nand g119(n2022 ,n3850 ,n1985);
    nor g120(n789 ,n10[8] ,n503);
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n225), .Q(n28[7]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1561), .Q(n18[6]));
    nand g123(n3007 ,n2725 ,n2904);
    nand g124(n2755 ,n28[5] ,n26[0]);
    nand g125(n3286 ,n3175 ,n3253);
    nor g126(n3646 ,n3637 ,n3645);
    nand g127(n1932 ,n3855 ,n1922);
    nand g128(n1656 ,n1267 ,n1018);
    nand g129(n3059 ,n2885 ,n3014);
    xnor g130(n2287 ,n2142 ,n2247);
    nand g131(n1106 ,n15[11] ,n443);
    nand g132(n855 ,n17[10] ,n484);
    nand g133(n1213 ,n9[0] ,n459);
    nand g134(n159 ,n24[6] ,n94);
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1510), .Q(n14[4]));
    nand g136(n2712 ,n27[7] ,n4[0]);
    nand g137(n877 ,n11[0] ,n478);
    nand g138(n638 ,n188 ,n445);
    nand g139(n882 ,n9[0] ,n496);
    nor g140(n834 ,n14[8] ,n467);
    xnor g141(n2211 ,n2137 ,n2101);
    or g142(n2637 ,n2552 ,n2613);
    xnor g143(n2202 ,n2135 ,n2155);
    nand g144(n1648 ,n1254 ,n1016);
    nand g145(n959 ,n20[5] ,n452);
    not g146(n106 ,n6);
    nor g147(n2271 ,n2177 ,n2244);
    nand g148(n1562 ,n1252 ,n675);
    xnor g149(n3330 ,n3223 ,n3242);
    nand g150(n330 ,n26[3] ,n247);
    xnor g151(n230 ,n152 ,n29[1]);
    nand g152(n2930 ,n2719 ,n2819);
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1565), .Q(n10[10]));
    nor g154(n2646 ,n2598 ,n2627);
    nand g155(n1381 ,n945 ,n571);
    nand g156(n2828 ,n28[7] ,n26[7]);
    nor g157(n1291 ,n805 ,n804);
    or g158(n3448 ,n3408 ,n3422);
    nand g159(n3767 ,n3716 ,n3747);
    or g160(n1314 ,n782 ,n813);
    nor g161(n1816 ,n29[8] ,n1794);
    nand g162(n1624 ,n1217 ,n1216);
    xnor g163(n1875 ,n26[15] ,n85);
    nand g164(n3555 ,n3535 ,n2705);
    xnor g165(n3543 ,n3518 ,n3492);
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1559), .Q(n18[8]));
    or g167(n3196 ,n3074 ,n3103);
    xnor g168(n2980 ,n2742 ,n2804);
    nand g169(n1346 ,n900 ,n530);
    xnor g170(n2959 ,n2832 ,n2800);
    nand g171(n2728 ,n28[3] ,n26[6]);
    nand g172(n1121 ,n10[5] ,n481);
    not g173(n245 ,n246);
    or g174(n34 ,n26[3] ,n32);
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n386), .Q(n26[0]));
    or g176(n2187 ,n2125 ,n2130);
    nand g177(n1458 ,n1090 ,n627);
    nor g178(n2192 ,n2072 ,n2153);
    nand g179(n3562 ,n3545 ,n3561);
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1362), .Q(n21[9]));
    nand g181(n630 ,n186 ,n445);
    nand g182(n352 ,n275 ,n340);
    nand g183(n2834 ,n28[1] ,n26[7]);
    nand g184(n750 ,n187 ,n490);
    nand g185(n2847 ,n27[3] ,n4[2]);
    nand g186(n885 ,n19[14] ,n482);
    nand g187(n1405 ,n854 ,n599);
    nor g188(n2159 ,n2106 ,n2118);
    nand g189(n1927 ,n3854 ,n1922);
    nand g190(n3079 ,n2870 ,n3035);
    nor g191(n132 ,n26[13] ,n26[14]);
    nor g192(n1808 ,n29[15] ,n1765);
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1441), .Q(n8[9]));
    nand g194(n1708 ,n1310 ,n1309);
    xnor g195(n2154 ,n1956 ,n2093);
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1552), .Q(n18[13]));
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1564), .Q(n18[4]));
    nand g198(n1475 ,n1109 ,n681);
    nand g199(n2663 ,n2635 ,n2648);
    nor g200(n1671 ,n1595 ,n1594);
    xnor g201(n2656 ,n2624 ,n2611);
    xnor g202(n189 ,n98 ,n4[6]);
    not g203(n2702 ,n2703);
    xnor g204(n3099 ,n3003 ,n2724);
    nand g205(n1988 ,n3850 ,n1960);
    nand g206(n1268 ,n21[6] ,n471);
    nand g207(n2031 ,n3851 ,n1985);
    nand g208(n2418 ,n3814 ,n4[4]);
    nand g209(n3582 ,n26[2] ,n4[2]);
    nand g210(n3181 ,n3091 ,n3136);
    nand g211(n1416 ,n989 ,n606);
    nand g212(n2019 ,n3853 ,n1986);
    not g213(n2784 ,n2783);
    nand g214(n1464 ,n1096 ,n631);
    xnor g215(n2606 ,n2580 ,n2528);
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n328), .Q(n25[6]));
    nand g217(n1587 ,n893 ,n1055);
    xor g218(n181 ,n4[12] ,n29[12]);
    not g219(n58 ,n26[4]);
    not g220(n55 ,n54);
    nand g221(n3763 ,n3743 ,n3742);
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n214), .Q(n27[5]));
    or g223(n2268 ,n2228 ,n2233);
    nand g224(n2820 ,n27[6] ,n4[6]);
    nand g225(n3061 ,n2871 ,n3013);
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n397), .Q(n26[15]));
    or g227(n3544 ,n3527 ,n3534);
    not g228(n480 ,n481);
    xnor g229(n2577 ,n2530 ,n2533);
    or g230(n3048 ,n2830 ,n2999);
    nand g231(n517 ,n191 ,n487);
    nor g232(n2906 ,n2840 ,n2754);
    nand g233(n732 ,n187 ,n480);
    nand g234(n1142 ,n9[15] ,n459);
    nor g235(n2305 ,n2253 ,n2285);
    nand g236(n401 ,n5[0] ,n359);
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1859), .Q(n5[2]));
    xor g238(n1895 ,n2118 ,n2106);
    nand g239(n2912 ,n2818 ,n2827);
    nand g240(n2269 ,n2116 ,n2250);
    nor g241(n1825 ,n29[5] ,n1781);
    xnor g242(n216 ,n151 ,n29[14]);
    nand g243(n3383 ,n3217 ,n3330);
    nand g244(n3779 ,n3727 ,n3723);
    nand g245(n2040 ,n1929 ,n1995);
    xnor g246(n3491 ,n3437 ,n3425);
    nand g247(n522 ,n182 ,n446);
    nand g248(n3695 ,n3861 ,n30[10]);
    or g249(n2885 ,n2736 ,n2808);
    nand g250(n1505 ,n1139 ,n744);
    nand g251(n3784 ,n3692 ,n3707);
    nand g252(n62 ,n26[1] ,n26[0]);
    nor g253(n2882 ,n2802 ,n2801);
    not g254(n3670 ,n2);
    nor g255(n1688 ,n1641 ,n1640);
    not g256(n2321 ,n2317);
    nand g257(n1247 ,n18[10] ,n456);
    nor g258(n57 ,n26[14] ,n55);
    nand g259(n1360 ,n920 ,n549);
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1408), .Q(n12[9]));
    nand g261(n1544 ,n1185 ,n707);
    nand g262(n2700 ,n2675 ,n2699);
    nand g263(n1138 ,n12[1] ,n476);
    nand g264(n357 ,n269 ,n312);
    nand g265(n861 ,n9[4] ,n496);
    nor g266(n1754 ,n1627 ,n1728);
    dff g267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1463), .Q(n16[2]));
    nand g268(n1506 ,n1141 ,n726);
    nand g269(n76 ,n26[9] ,n74);
    nand g270(n150 ,n25[3] ,n94);
    nand g271(n3452 ,n3408 ,n3422);
    nor g272(n821 ,n13[9] ,n500);
    xnor g273(n3397 ,n3310 ,n3188);
    or g274(n3453 ,n3350 ,n3420);
    dff g275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1354), .Q(n13[11]));
    nand g276(n1529 ,n1162 ,n746);
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1498), .Q(n8[4]));
    nand g278(n730 ,n192 ,n480);
    nand g279(n2010 ,n3857 ,n1964);
    nand g280(n1027 ,n11[10] ,n441);
    not g281(n105 ,n28[2]);
    xnor g282(n3623 ,n3849 ,n3833);
    xnor g283(n2127 ,n2060 ,n1955);
    nor g284(n247 ,n172 ,n202);
    nand g285(n3088 ,n2895 ,n3037);
    nor g286(n1290 ,n803 ,n790);
    nor g287(n774 ,n17[9] ,n469);
    nand g288(n3058 ,n2881 ,n3030);
    nor g289(n124 ,n26[2] ,n26[3]);
    nand g290(n1545 ,n1186 ,n708);
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1514), .Q(n22[15]));
    nand g292(n1173 ,n22[1] ,n451);
    not g293(n2570 ,n2562);
    nor g294(n2627 ,n2596 ,n2612);
    nand g295(n2648 ,n2640 ,n2638);
    or g296(n2898 ,n2727 ,n2740);
    nand g297(n1097 ,n10[12] ,n481);
    nand g298(n945 ,n13[2] ,n448);
    nand g299(n738 ,n181 ,n490);
    nand g300(n2645 ,n2621 ,n2629);
    nand g301(n1591 ,n1064 ,n1063);
    nor g302(n1675 ,n1632 ,n1605);
    xnor g303(n3314 ,n3239 ,n3262);
    nor g304(n1790 ,n359 ,n1772);
    xnor g305(n226 ,n150 ,n29[11]);
    nand g306(n1725 ,n1689 ,n1688);
    xnor g307(n3130 ,n2984 ,n2756);
    nand g308(n147 ,n1879 ,n94);
    not g309(n2245 ,n2244);
    nand g310(n1151 ,n22[14] ,n451);
    not g311(n3222 ,n3209);
    not g312(n488 ,n489);
    nand g313(n1480 ,n1114 ,n684);
    nand g314(n1991 ,n3858 ,n1964);
    not g315(n140 ,n141);
    nor g316(n2447 ,n2406 ,n2423);
    xnor g317(n3311 ,n3258 ,n3191);
    not g318(n367 ,n351);
    nand g319(n3600 ,n3581 ,n3599);
    not g320(n2350 ,n2349);
    nor g321(n3654 ,n3625 ,n3653);
    dff g322(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1445), .Q(n11[2]));
    xnor g323(n3861 ,n3624 ,n3655);
    or g324(n29[10] ,n3767 ,n3795);
    not g325(n100 ,n29[2]);
    nor g326(n2616 ,n2593 ,n2594);
    xnor g327(n3626 ,n3843 ,n3827);
    nand g328(n1317 ,n970 ,n607);
    nand g329(n1517 ,n1152 ,n751);
    not g330(n1960 ,n1961);
    nand g331(n1453 ,n1079 ,n674);
    nand g332(n883 ,n19[0] ,n472);
    nand g333(n397 ,n331 ,n367);
    not g334(n359 ,n360);
    nand g335(n415 ,n27[3] ,n365);
    nand g336(n2653 ,n2583 ,n2636);
    nand g337(n1573 ,n1021 ,n1219);
    nand g338(n1947 ,n1914 ,n1940);
    nand g339(n3750 ,n3845 ,n3685);
    nand g340(n1495 ,n1128 ,n735);
    nand g341(n3754 ,n3846 ,n3685);
    dff g342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1511), .Q(n9[14]));
    nand g343(n1861 ,n47 ,n46);
    nor g344(n1869 ,n75 ,n77);
    nand g345(n2506 ,n5[0] ,n2445);
    nand g346(n2000 ,n3854 ,n1964);
    xnor g347(n3844 ,n2381 ,n2390);
    nand g348(n3796 ,n3752 ,n3774);
    not g349(n2734 ,n2733);
    not g350(n2407 ,n5[0]);
    nand g351(n2695 ,n2679 ,n2694);
    not g352(n2760 ,n2759);
    nand g353(n3019 ,n2860 ,n2911);
    nand g354(n3687 ,n3869 ,n30[2]);
    xnor g355(n2969 ,n2718 ,n2821);
    nand g356(n2786 ,n28[6] ,n26[3]);
    nor g357(n2863 ,n2706 ,n2707);
    or g358(n2907 ,n2742 ,n2804);
    nand g359(n3752 ,n3835 ,n3685);
    nand g360(n719 ,n180 ,n480);
    nand g361(n1511 ,n1147 ,n695);
    nand g362(n2922 ,n2800 ,n2832);
    nand g363(n2061 ,n1981 ,n2019);
    nand g364(n613 ,n186 ,n485);
    xnor g365(n2380 ,n2365 ,n2350);
    dff g366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1736), .Q(n7));
    or g367(n1855 ,n1804 ,n1850);
    nand g368(n696 ,n180 ,n458);
    xnor g369(n3108 ,n2959 ,n2841);
    nand g370(n154 ,n1877 ,n94);
    nor g371(n2169 ,n2100 ,n2149);
    xnor g372(n2381 ,n2364 ,n2339);
    nor g373(n2234 ,n2170 ,n2218);
    nand g374(n1031 ,n22[4] ,n463);
    or g375(n3348 ,n3238 ,n3272);
    xnor g376(n30[10] ,n2676 ,n2698);
    not g377(n2441 ,n2442);
    nand g378(n3571 ,n3547 ,n3570);
    nand g379(n1444 ,n1050 ,n700);
    nand g380(n1041 ,n8[11] ,n489);
    not g381(n249 ,n248);
    nand g382(n3718 ,n3818 ,n3684);
    nand g383(n3026 ,n2760 ,n2937);
    nand g384(n920 ,n13[9] ,n448);
    nand g385(n3186 ,n3049 ,n3145);
    nor g386(n449 ,n138 ,n416);
    nand g387(n3198 ,n3069 ,n3138);
    xnor g388(n2579 ,n2535 ,n2465);
    not g389(n3299 ,n3298);
    nand g390(n173 ,n2 ,n110);
    nand g391(n1645 ,n1239 ,n1176);
    not g392(n3269 ,n3268);
    xnor g393(n3464 ,n3397 ,n3421);
    xnor g394(n3400 ,n3312 ,n3272);
    nor g395(n2289 ,n2114 ,n2272);
    nand g396(n316 ,n1890 ,n245);
    nand g397(n918 ,n21[12] ,n454);
    nor g398(n770 ,n11[5] ,n479);
    xnor g399(n3134 ,n2997 ,n2901);
    dff g400(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1857), .Q(n5[12]));
    or g401(n1848 ,n1812 ,n1828);
    dff g402(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1485), .Q(n10[6]));
    nand g403(n1941 ,n1908 ,n1921);
    dff g404(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n231), .Q(n27[0]));
    nand g405(n3775 ,n3717 ,n3746);
    dff g406(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n375), .Q(n24[3]));
    nand g407(n655 ,n186 ,n450);
    xnor g408(n2209 ,n2130 ,n2125);
    xor g409(n1959 ,n1943 ,n1949);
    nand g410(n2013 ,n3857 ,n1958);
    dff g411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1524), .Q(n22[9]));
    nor g412(n812 ,n16[5] ,n498);
    nand g413(n1319 ,n850 ,n593);
    nand g414(n676 ,n179 ,n442);
    nor g415(n485 ,n137 ,n411);
    nand g416(n531 ,n204 ,n446);
    nor g417(n3674 ,n3862 ,n30[9]);
    nand g418(n1131 ,n14[13] ,n491);
    nand g419(n3618 ,n3848 ,n3832);
    nand g420(n2242 ,n2191 ,n2225);
    nand g421(n3091 ,n2886 ,n3015);
    nand g422(n2047 ,n3858 ,n1985);
    nand g423(n899 ,n23[3] ,n447);
    nand g424(n1600 ,n1187 ,n973);
    xnor g425(n3443 ,n3388 ,n3412);
    nand g426(n2923 ,n2823 ,n2745);
    nor g427(n3655 ,n3608 ,n3654);
    not g428(n63 ,n62);
    nand g429(n3790 ,n3725 ,n3724);
    nand g430(n3798 ,n3757 ,n3784);
    xnor g431(n2367 ,n2319 ,n2326);
    or g432(n2899 ,n2794 ,n2743);
    nand g433(n3755 ,n3836 ,n3685);
    nand g434(n1375 ,n937 ,n564);
    xnor g435(n3838 ,n2304 ,n2299);
    xnor g436(n3241 ,n3097 ,n2905);
    nand g437(n579 ,n185 ,n453);
    xnor g438(n2130 ,n1955 ,n2061);
    nand g439(n78 ,n26[10] ,n77);
    not g440(n474 ,n475);
    nand g441(n1029 ,n11[9] ,n441);
    nor g442(n3577 ,n26[7] ,n4[7]);
    dff g443(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n376), .Q(n25[1]));
    nor g444(n772 ,n11[8] ,n479);
    nand g445(n915 ,n21[14] ,n454);
    nand g446(n1349 ,n907 ,n537);
    nand g447(n1352 ,n911 ,n541);
    nor g448(n3060 ,n2896 ,n3041);
    nand g449(n1456 ,n1088 ,n626);
    nand g450(n3204 ,n3117 ,n3116);
    dff g451(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n438), .Q(n26[5]));
    nor g452(n290 ,n201 ,n215);
    xnor g453(n2131 ,n2086 ,n1955);
    nand g454(n3451 ,n3370 ,n3425);
    nor g455(n763 ,n10[5] ,n503);
    nand g456(n1909 ,n28[0] ,n27[0]);
    nand g457(n2306 ,n2248 ,n2283);
    not g458(n2214 ,n2213);
    nand g459(n3234 ,n3088 ,n3195);
    nor g460(n1668 ,n1587 ,n1586);
    nand g461(n3258 ,n3144 ,n3212);
    nand g462(n1925 ,n3850 ,n1922);
    nand g463(n167 ,n29[7] ,n1885);
    xnor g464(n3517 ,n3443 ,n3489);
    nor g465(n3804 ,n2565 ,n2553);
    nand g466(n2005 ,n3854 ,n1963);
    nand g467(n1822 ,n29[11] ,n1791);
    nand g468(n631 ,n204 ,n445);
    nor g469(n291 ,n1889 ,n246);
    nand g470(n2076 ,n1967 ,n2052);
    dff g471(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1512), .Q(n8[3]));
    nand g472(n2938 ,n2826 ,n2730);
    not g473(n2467 ,n2466);
    nor g474(n2434 ,n2408 ,n2421);
    nand g475(n3414 ,n3341 ,n3361);
    nand g476(n2822 ,n28[7] ,n26[5]);
    nand g477(n2751 ,n27[3] ,n4[3]);
    xnor g478(n1868 ,n26[8] ,n73);
    nand g479(n1135 ,n10[1] ,n481);
    xor g480(n2957 ,n2785 ,n2737);
    nand g481(n3259 ,n3140 ,n3198);
    xnor g482(n3232 ,n3124 ,n3075);
    nand g483(n271 ,n1862 ,n206);
    xnor g484(n2667 ,n2641 ,n2621);
    xnor g485(n2999 ,n2849 ,n2837);
    nand g486(n2520 ,n2472 ,n2485);
    not g487(n3459 ,n3458);
    nand g488(n912 ,n19[15] ,n472);
    nand g489(n866 ,n17[3] ,n484);
    nand g490(n714 ,n184 ,n488);
    nand g491(n3620 ,n3836 ,n3820);
    nand g492(n1880 ,n35 ,n34);
    nand g493(n1043 ,n11[6] ,n441);
    xnor g494(n2372 ,n2327 ,n2351);
    nand g495(n2740 ,n27[7] ,n4[1]);
    nand g496(n1327 ,n876 ,n534);
    xnor g497(n2676 ,n2632 ,n2664);
    nor g498(n3504 ,n3443 ,n3489);
    or g499(n1782 ,n359 ,n1763);
    nor g500(n2599 ,n2543 ,n2582);
    xnor g501(n3441 ,n3311 ,n3413);
    nor g502(n1693 ,n1655 ,n1654);
    not g503(n3240 ,n3239);
    nor g504(n800 ,n22[3] ,n462);
    dff g505(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1529), .Q(n8[2]));
    nand g506(n87 ,n28[1] ,n28[0]);
    nand g507(n2173 ,n2097 ,n2151);
    xnor g508(n3239 ,n3099 ,n2904);
    nand g509(n2681 ,n2661 ,n2668);
    nand g510(n1343 ,n897 ,n527);
    xnor g511(n2989 ,n2721 ,n2790);
    not g512(n2954 ,n2939);
    not g513(n446 ,n447);
    nand g514(n1834 ,n395 ,n1800);
    nand g515(n1331 ,n867 ,n567);
    nor g516(n2244 ,n2184 ,n2221);
    nand g517(n305 ,n26[4] ,n247);
    nor g518(n1752 ,n1604 ,n1733);
    xnor g519(n3635 ,n3847 ,n3831);
    xnor g520(n234 ,n163 ,n29[9]);
    xnor g521(n2110 ,n1945 ,n2045);
    nand g522(n1187 ,n14[15] ,n466);
    not g523(n2949 ,n2948);
    not g524(n490 ,n491);
    nand g525(n416 ,n28[2] ,n362);
    nand g526(n709 ,n186 ,n458);
    nand g527(n2062 ,n1968 ,n2020);
    or g528(n3373 ,n3217 ,n3330);
    nand g529(n2559 ,n2509 ,n2527);
    nor g530(n1278 ,n794 ,n795);
    nand g531(n1465 ,n1097 ,n720);
    nor g532(n54 ,n26[13] ,n52);
    nor g533(n817 ,n18[9] ,n475);
    xnor g534(n3370 ,n3266 ,n3218);
    nand g535(n3376 ,n3219 ,n3346);
    nand g536(n1234 ,n18[10] ,n474);
    nand g537(n266 ,n24[3] ,n201);
    nand g538(n2805 ,n27[7] ,n4[2]);
    nand g539(n276 ,n1866 ,n206);
    dff g540(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1526), .Q(n22[8]));
    or g541(n3151 ,n3058 ,n3078);
    nand g542(n3233 ,n3111 ,n3188);
    nand g543(n1073 ,n16[10] ,n444);
    nand g544(n1415 ,n988 ,n591);
    nand g545(n3728 ,n3820 ,n3684);
    nand g546(n3035 ,n2842 ,n2922);
    not g547(n414 ,n415);
    nand g548(n1353 ,n913 ,n544);
    xnor g549(n1882 ,n27[3] ,n93);
    nand g550(n1830 ,n418 ,n1805);
    xnor g551(n1942 ,n1901 ,n1915);
    nand g552(n1238 ,n18[15] ,n456);
    nand g553(n1208 ,n21[13] ,n471);
    nand g554(n1132 ,n8[4] ,n489);
    nand g555(n1514 ,n1149 ,n639);
    nor g556(n2333 ,n2243 ,n2310);
    nand g557(n328 ,n254 ,n258);
    nand g558(n1549 ,n1213 ,n697);
    nor g559(n445 ,n135 ,n411);
    nand g560(n1629 ,n1222 ,n958);
    nand g561(n911 ,n13[12] ,n448);
    or g562(n2412 ,n3810 ,n4[0]);
    nand g563(n984 ,n19[7] ,n482);
    nand g564(n1318 ,n848 ,n892);
    nand g565(n1386 ,n952 ,n580);
    nand g566(n2858 ,n28[7] ,n26[1]);
    xnor g567(n30[4] ,n2665 ,n2663);
    nand g568(n3044 ,n2772 ,n2944);
    xnor g569(n2997 ,n2846 ,n2858);
    nand g570(n2626 ,n2586 ,n2610);
    nand g571(n2120 ,n1955 ,n2075);
    nand g572(n2053 ,n3856 ,n2015);
    nand g573(n2090 ,n2007 ,n2031);
    nand g574(n355 ,n271 ,n310);
    nand g575(n1046 ,n8[13] ,n489);
    nand g576(n3599 ,n3594 ,n3598);
    not g577(n2753 ,n2752);
    nand g578(n3381 ,n3351 ,n3327);
    nand g579(n2926 ,n2834 ,n2825);
    nand g580(n1569 ,n1265 ,n713);
    nor g581(n2524 ,n2466 ,n2503);
    dff g582(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1431), .Q(n8[12]));
    or g583(n2890 ,n2723 ,n2816);
    nand g584(n3006 ,n2798 ,n2948);
    nand g585(n2011 ,n3857 ,n1963);
    nand g586(n3731 ,n3839 ,n3685);
    nand g587(n3565 ,n3564 ,n3555);
    nor g588(n1470 ,n1 ,n842);
    dff g589(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1394), .Q(n20[4]));
    nor g590(n3708 ,n3698 ,n3680);
    nand g591(n3537 ,n3497 ,n3525);
    dff g592(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1484), .Q(n15[5]));
    nand g593(n1374 ,n938 ,n565);
    nand g594(n746 ,n186 ,n488);
    nor g595(n2633 ,n2615 ,n2616);
    nor g596(n3647 ,n3610 ,n3646);
    nor g597(n818 ,n20[9] ,n460);
    xnor g598(n2575 ,n2515 ,n2510);
    nor g599(n815 ,n20[8] ,n460);
    xnor g600(n3843 ,n2360 ,n2388);
    nand g601(n1259 ,n18[4] ,n456);
    nand g602(n1074 ,n23[0] ,n465);
    nand g603(n467 ,n210 ,n404);
    nand g604(n648 ,n184 ,n450);
    not g605(n1989 ,n1988);
    nand g606(n2561 ,n2510 ,n2515);
    nand g607(n879 ,n8[0] ,n494);
    nand g608(n1254 ,n18[7] ,n474);
    nand g609(n2787 ,n27[4] ,n4[6]);
    nor g610(n782 ,n19[8] ,n473);
    nand g611(n1101 ,n8[7] ,n489);
    nand g612(n2225 ,n1896 ,n2168);
    not g613(n2994 ,n2993);
    nand g614(n3034 ,n2770 ,n2933);
    nand g615(n3794 ,n3749 ,n3769);
    xnor g616(n1917 ,n28[6] ,n27[6]);
    xnor g617(n3227 ,n3155 ,n3153);
    nand g618(n1461 ,n1093 ,n629);
    nand g619(n3777 ,n3735 ,n3754);
    or g620(n3183 ,n3077 ,n3121);
    dff g621(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1562), .Q(n11[15]));
    nand g622(n375 ,n266 ,n296);
    nor g623(n2477 ,n2408 ,n2446);
    dff g624(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1842), .Q(n5[7]));
    nand g625(n2171 ,n1956 ,n2131);
    nor g626(n2555 ,n2525 ,n2519);
    nand g627(n2012 ,n3858 ,n1963);
    or g628(n42 ,n26[7] ,n40);
    nand g629(n3261 ,n3005 ,n3210);
    nand g630(n3289 ,n3218 ,n3235);
    dff g631(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1500), .Q(n10[1]));
    nand g632(n1126 ,n14[15] ,n491);
    nand g633(n2804 ,n28[4] ,n26[3]);
    nand g634(n725 ,n178 ,n488);
    or g635(n2892 ,n2828 ,n2793);
    nand g636(n1130 ,n10[2] ,n481);
    nand g637(n1273 ,n11[12] ,n441);
    nand g638(n3139 ,n2940 ,n3095);
    nor g639(n2517 ,n2455 ,n2478);
    nand g640(n1593 ,n878 ,n1072);
    nand g641(n1553 ,n1182 ,n757);
    xnor g642(n2142 ,n2067 ,n1946);
    nand g643(n3160 ,n3007 ,n3071);
    nand g644(n1248 ,n20[14] ,n461);
    nand g645(n2348 ,n2320 ,n2326);
    nand g646(n1606 ,n847 ,n968);
    nand g647(n2397 ,n2369 ,n2396);
    nand g648(n986 ,n10[12] ,n502);
    nand g649(n1908 ,n28[4] ,n28[3]);
    nand g650(n3711 ,n30[5] ,n3699);
    nand g651(n1022 ,n8[12] ,n489);
    xnor g652(n3119 ,n2975 ,n2749);
    not g653(n1926 ,n27[0]);
    nand g654(n1023 ,n14[6] ,n466);
    nand g655(n558 ,n178 ,n455);
    nand g656(n619 ,n182 ,n450);
    nand g657(n403 ,n5[5] ,n359);
    nand g658(n1982 ,n3851 ,n1960);
    nand g659(n735 ,n188 ,n490);
    not g660(n2708 ,n27[4]);
    nand g661(n659 ,n186 ,n457);
    nand g662(n3771 ,n3721 ,n3750);
    nor g663(n3174 ,n3117 ,n3116);
    not g664(n1898 ,n3854);
    nor g665(n68 ,n26[5] ,n67);
    xnor g666(n3823 ,n3479 ,n3494);
    not g667(n2591 ,n2590);
    nand g668(n948 ,n20[12] ,n452);
    nor g669(n1694 ,n1657 ,n1656);
    xnor g670(n2128 ,n2084 ,n1955);
    nand g671(n1341 ,n895 ,n525);
    nand g672(n867 ,n17[1] ,n484);
    not g673(n3085 ,n3084);
    or g674(n2875 ,n2799 ,n2731);
    nor g675(n2449 ,n2406 ,n2419);
    nand g676(n1385 ,n951 ,n579);
    or g677(n2876 ,n2722 ,n2820);
    nand g678(n3064 ,n2873 ,n3022);
    nand g679(n329 ,n255 ,n282);
    nand g680(n1603 ,n1190 ,n1012);
    xnor g681(n3170 ,n3061 ,n2903);
    not g682(n372 ,n357);
    nand g683(n2504 ,n5[0] ,n2441);
    not g684(n454 ,n455);
    not g685(n2359 ,n2358);
    not g686(n3001 ,n3000);
    or g687(n2666 ,n2653 ,n2655);
    nand g688(n589 ,n180 ,n487);
    dff g689(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1549), .Q(n9[0]));
    nand g690(n3158 ,n3008 ,n3070);
    xnor g691(n3117 ,n2971 ,n2783);
    nor g692(n3245 ,n3130 ,n3216);
    xnor g693(n3392 ,n3320 ,n3288);
    nand g694(n3030 ,n2845 ,n2924);
    dff g695(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1843), .Q(n5[6]));
    nor g696(n2325 ,n2275 ,n2308);
    nand g697(n1136 ,n14[10] ,n491);
    xnor g698(n3550 ,n3537 ,n3520);
    xnor g699(n3846 ,n2382 ,n2394);
    xnor g700(n3434 ,n3322 ,n3416);
    dff g701(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1410), .Q(n12[8]));
    dff g702(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1660), .Q(n15[13]));
    xnor g703(n3837 ,n2251 ,n2246);
    xnor g704(n2607 ,n2572 ,n2587);
    nand g705(n324 ,n252 ,n259);
    nor g706(n2452 ,n2407 ,n2424);
    not g707(n500 ,n501);
    not g708(n2748 ,n2747);
    not g709(n2105 ,n2104);
    nand g710(n893 ,n19[1] ,n472);
    nand g711(n1325 ,n863 ,n594);
    nand g712(n3084 ,n2866 ,n3021);
    nor g713(n2511 ,n2453 ,n2481);
    nor g714(n2537 ,n2464 ,n2473);
    nand g715(n1472 ,n1105 ,n679);
    xor g716(n3169 ,n3074 ,n3088);
    or g717(n2893 ,n2814 ,n2807);
    nand g718(n3781 ,n3760 ,n3729);
    nand g719(n149 ,n24[2] ,n94);
    not g720(n320 ,n319);
    nand g721(n3664 ,n3628 ,n3663);
    nand g722(n3036 ,n2857 ,n2916);
    nand g723(n526 ,n189 ,n446);
    nand g724(n1482 ,n1129 ,n725);
    nand g725(n1061 ,n23[15] ,n465);
    nand g726(n1995 ,n3855 ,n1964);
    or g727(n1795 ,n359 ,n1761);
    nand g728(n382 ,n270 ,n297);
    nand g729(n175 ,n27[1] ,n108);
    or g730(n3384 ,n3335 ,n3332);
    or g731(n3439 ,n3398 ,n3421);
    nand g732(n1556 ,n1247 ,n641);
    dff g733(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1333), .Q(n23[15]));
    nor g734(n2273 ,n2246 ,n2231);
    nand g735(n2924 ,n2835 ,n2803);
    xnor g736(n3359 ,n3268 ,n3280);
    xnor g737(n3106 ,n2983 ,n2847);
    nand g738(n1827 ,n29[12] ,n1790);
    nand g739(n2502 ,n5[0] ,n2436);
    xnor g740(n2966 ,n2740 ,n2727);
    xnor g741(n1962 ,n1946 ,n1925);
    xnor g742(n3839 ,n2303 ,n2343);
    dff g743(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n378), .Q(n25[3]));
    nand g744(n1179 ,n9[7] ,n459);
    not g745(n3628 ,n3627);
    nand g746(n2660 ,n2620 ,n2647);
    xor g747(n179 ,n4[15] ,n29[15]);
    xnor g748(n3639 ,n3844 ,n3828);
    nor g749(n3652 ,n3641 ,n3651);
    nand g750(n1454 ,n1084 ,n625);
    xnor g751(n3521 ,n3462 ,n3482);
    nand g752(n1936 ,n1917 ,n1910);
    dff g753(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1422), .Q(n19[1]));
    nand g754(n2762 ,n27[0] ,n4[4]);
    xnor g755(n2210 ,n2147 ,n2105);
    nand g756(n759 ,n183 ,n488);
    xnor g757(n3278 ,n3171 ,n3069);
    xnor g758(n3185 ,n2961 ,n3096);
    dff g759(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1569), .Q(n11[13]));
    nand g760(n606 ,n189 ,n487);
    nand g761(n255 ,n29[15] ,n202);
    not g762(n65 ,n64);
    nor g763(n1817 ,n95 ,n1785);
    nand g764(n3447 ,n3292 ,n3426);
    xnor g765(n190 ,n96 ,n4[7]);
    nor g766(n2371 ,n2291 ,n2346);
    nand g767(n968 ,n8[14] ,n494);
    or g768(n3644 ,n3634 ,n3643);
    nand g769(n3090 ,n2887 ,n3032);
    or g770(n1785 ,n359 ,n1767);
    xnor g771(n2644 ,n2586 ,n2610);
    nand g772(n3144 ,n2796 ,n3084);
    dff g773(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1488), .Q(n10[5]));
    dff g774(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1525), .Q(n14[0]));
    nand g775(n3757 ,n3843 ,n3685);
    nand g776(n1597 ,n1082 ,n1081);
    nand g777(n884 ,n10[14] ,n502);
    nand g778(n515 ,n184 ,n446);
    nor g779(n3214 ,n3080 ,n3122);
    nor g780(n806 ,n18[2] ,n475);
    xnor g781(n2121 ,n2069 ,n2071);
    xnor g782(n235 ,n162 ,n29[10]);
    nand g783(n169 ,n29[5] ,n1887);
    or g784(n3552 ,n3532 ,n3543);
    not g785(n2201 ,n2188);
    xnor g786(n3520 ,n3480 ,n3483);
    nand g787(n3065 ,n2898 ,n3028);
    nand g788(n3494 ,n3453 ,n3473);
    nand g789(n1793 ,n360 ,n1776);
    nor g790(n2351 ,n2307 ,n2336);
    not g791(n3221 ,n3206);
    nand g792(n2767 ,n28[6] ,n26[1]);
    nand g793(n917 ,n21[13] ,n454);
    nand g794(n1232 ,n13[11] ,n501);
    not g795(n136 ,n137);
    nand g796(n341 ,n26[11] ,n247);
    or g797(n1792 ,n359 ,n1775);
    xnor g798(n3819 ,n2900 ,n3225);
    nand g799(n705 ,n189 ,n458);
    nand g800(n155 ,n25[4] ,n94);
    nand g801(n2037 ,n1933 ,n1994);
    dff g802(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n21[10]));
    nand g803(n1344 ,n898 ,n528);
    or g804(n1780 ,n359 ,n1774);
    nand g805(n3187 ,n3051 ,n3135);
    nand g806(n293 ,n202 ,n235);
    nand g807(n1616 ,n1206 ,n976);
    nand g808(n1800 ,n95 ,n1767);
    nand g809(n308 ,n1872 ,n245);
    xnor g810(n30[3] ,n2643 ,n2640);
    dff g811(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1548), .Q(n9[1]));
    dff g812(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1517), .Q(n14[2]));
    nand g813(n653 ,n192 ,n457);
    xor g814(n2987 ,n2702 ,n2818);
    nand g815(n3005 ,n2734 ,n2900);
    nor g816(n3704 ,n3698 ,n3678);
    nand g817(n1189 ,n20[15] ,n461);
    or g818(n3295 ,n3118 ,n2704);
    nand g819(n682 ,n183 ,n442);
    xor g820(n1922 ,n27[0] ,n28[0]);
    nor g821(n2220 ,n2135 ,n2199);
    dff g822(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1453), .Q(n11[0]));
    xnor g823(n3116 ,n2970 ,n2751);
    not g824(n3630 ,n3629);
    nand g825(n2094 ,n2011 ,n2033);
    nand g826(n3380 ,n3160 ,n3337);
    nor g827(n829 ,n12[5] ,n477);
    nand g828(n1740 ,n1288 ,n1713);
    nand g829(n1369 ,n929 ,n557);
    xnor g830(n222 ,n98 ,n154);
    nand g831(n2548 ,n2465 ,n2536);
    nand g832(n3405 ,n3353 ,n3362);
    nor g833(n2389 ,n2352 ,n2388);
    or g834(n2868 ,n2720 ,n2789);
    nand g835(n2290 ,n2249 ,n2268);
    nand g836(n1389 ,n955 ,n583);
    nor g837(n3660 ,n3639 ,n3659);
    nand g838(n2027 ,n3852 ,n1985);
    or g839(n2638 ,n2567 ,n2609);
    nand g840(n1258 ,n15[13] ,n493);
    nand g841(n3773 ,n3720 ,n3719);
    nand g842(n2071 ,n1969 ,n2050);
    nand g843(n1799 ,n97 ,n1763);
    nand g844(n3513 ,n3441 ,n3490);
    nand g845(n1005 ,n8[6] ,n494);
    nand g846(n681 ,n185 ,n442);
    nand g847(n3712 ,n3823 ,n3684);
    nor g848(n3094 ,n2865 ,n3042);
    nor g849(n407 ,n105 ,n383);
    nand g850(n560 ,n181 ,n487);
    xnor g851(n2123 ,n2081 ,n1955);
    nand g852(n1626 ,n985 ,n1220);
    nand g853(n975 ,n10[13] ,n502);
    nand g854(n543 ,n191 ,n483);
    not g855(n2387 ,n2386);
    dff g856(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1560), .Q(n18[7]));
    nor g857(n1295 ,n807 ,n827);
    nand g858(n1019 ,n12[7] ,n486);
    nand g859(n1267 ,n22[6] ,n463);
    nor g860(n1787 ,n359 ,n1764);
    dff g861(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1523), .Q(n22[10]));
    dff g862(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1347), .Q(n23[1]));
    nand g863(n399 ,n337 ,n370);
    nor g864(n1287 ,n800 ,n765);
    nor g865(n3197 ,n3107 ,n3100);
    nand g866(n1087 ,n14[0] ,n466);
    dff g867(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1409), .Q(n19[9]));
    nand g868(n1345 ,n899 ,n529);
    xor g869(n3810 ,n28[0] ,n27[0]);
    dff g870(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1329), .Q(n17[3]));
    nor g871(n2296 ,n2197 ,n2257);
    xnor g872(n3437 ,n3370 ,n3415);
    nand g873(n314 ,n1869 ,n245);
    xnor g874(n3862 ,n3625 ,n3653);
    xnor g875(n3857 ,n3587 ,n3606);
    xnor g876(n3390 ,n3299 ,n3328);
    nand g877(n3598 ,n3582 ,n3597);
    nor g878(n2246 ,n2176 ,n2227);
    dff g879(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1327), .Q(n17[5]));
    nand g880(n979 ,n9[14] ,n496);
    nand g881(n1362 ,n923 ,n602);
    nor g882(n2070 ,n1973 ,n2051);
    nor g883(n2270 ,n2113 ,n2239);
    nor g884(n1682 ,n1623 ,n1622);
    nand g885(n1574 ,n1023 ,n1005);
    nor g886(n803 ,n20[3] ,n460);
    nand g887(n2733 ,n28[0] ,n26[1]);
    nand g888(n3318 ,n3240 ,n3270);
    nor g889(n1681 ,n1621 ,n1620);
    nand g890(n1395 ,n965 ,n590);
    xnor g891(n3854 ,n3600 ,n3584);
    not g892(n2853 ,n2852);
    nand g893(n3726 ,n3833 ,n3684);
    xnor g894(n3190 ,n3046 ,n3062);
    xnor g895(n3807 ,n3635 ,n3665);
    nand g896(n3291 ,n3118 ,n2704);
    nor g897(n1677 ,n1609 ,n1608);
    xor g898(n3812 ,n28[2] ,n27[2]);
    nand g899(n3062 ,n2868 ,n3023);
    nor g900(n1751 ,n1597 ,n1732);
    nand g901(n2790 ,n28[7] ,n26[6]);
    nand g902(n1257 ,n12[7] ,n476);
    nand g903(n3461 ,n3404 ,n3427);
    nand g904(n1222 ,n15[12] ,n493);
    nor g905(n3606 ,n3578 ,n3605);
    nand g906(n978 ,n17[13] ,n468);
    nor g907(n1664 ,n1577 ,n1576);
    nand g908(n3525 ,n3431 ,n3496);
    nand g909(n588 ,n192 ,n453);
    xor g910(n3226 ,n3115 ,n3161);
    not g911(n3329 ,n3328);
    nand g912(n3557 ,n3530 ,n3548);
    nand g913(n516 ,n180 ,n483);
    xor g914(n3852 ,n3592 ,n3596);
    nand g915(n1275 ,n23[10] ,n447);
    dff g916(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1849), .Q(n5[13]));
    not g917(n411 ,n410);
    nand g918(n1550 ,n1238 ,n646);
    dff g919(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1448), .Q(n16[11]));
    nand g920(n3015 ,n2764 ,n2938);
    nor g921(n86 ,n28[1] ,n28[0]);
    nand g922(n2045 ,n1932 ,n2000);
    dff g923(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1458), .Q(n16[5]));
    nand g924(n1063 ,n14[1] ,n466);
    nand g925(n1111 ,n10[8] ,n481);
    not g926(n3672 ,n3807);
    or g927(n1777 ,n1710 ,n1758);
    nand g928(n3143 ,n2903 ,n3059);
    nand g929(n3316 ,n3280 ,n3269);
    nor g930(n3661 ,n3614 ,n3660);
    xnor g931(n2206 ,n2127 ,n2145);
    xnor g932(n2157 ,n1956 ,n2089);
    nand g933(n1972 ,n3852 ,n1958);
    xor g934(n1896 ,n2120 ,n2110);
    or g935(n3449 ,n3370 ,n3425);
    nand g936(n544 ,n179 ,n455);
    nand g937(n1581 ,n1037 ,n1036);
    xnor g938(n3629 ,n3848 ,n3832);
    nand g939(n250 ,n29[7] ,n200);
    nand g940(n69 ,n26[5] ,n67);
    nor g941(n2900 ,n2864 ,n2788);
    nand g942(n3192 ,n2892 ,n3139);
    nand g943(n165 ,n25[1] ,n94);
    nand g944(n1660 ,n1104 ,n678);
    dff g945(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1396), .Q(n20[2]));
    xnor g946(n2961 ,n2823 ,n2745);
    nand g947(n1210 ,n18[13] ,n474);
    nor g948(n1284 ,n816 ,n764);
    nand g949(n1492 ,n1125 ,n693);
    nand g950(n640 ,n188 ,n450);
    nand g951(n1194 ,n8[0] ,n489);
    nor g952(n2309 ,n2288 ,n2254);
    nand g953(n1704 ,n1299 ,n1298);
    nand g954(n1152 ,n14[2] ,n491);
    nand g955(n565 ,n204 ,n455);
    nand g956(n1448 ,n1069 ,n621);
    nor g957(n1292 ,n767 ,n784);
    nand g958(n3534 ,n3510 ,n3522);
    nand g959(n545 ,n188 ,n455);
    or g960(n2877 ,n2824 ,n2712);
    dff g961(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1841), .Q(n5[8]));
    nand g962(n2621 ,n2550 ,n2603);
    nand g963(n868 ,n17[7] ,n468);
    nand g964(n1149 ,n22[15] ,n451);
    not g965(n3189 ,n3188);
    not g966(n2438 ,n2439);
    nor g967(n3360 ,n3299 ,n3329);
    nor g968(n3663 ,n3612 ,n3662);
    nand g969(n358 ,n167 ,n285);
    nor g970(n792 ,n12[3] ,n477);
    nor g971(n1714 ,n1703 ,n1702);
    nand g972(n3785 ,n3734 ,n3733);
    nand g973(n2736 ,n28[1] ,n26[2]);
    nand g974(n1602 ,n1048 ,n852);
    not g975(n3321 ,n3320);
    xnor g976(n3463 ,n3423 ,n3411);
    nand g977(n1571 ,n1046 ,n749);
    nand g978(n3055 ,n2877 ,n3044);
    nand g979(n41 ,n26[6] ,n38);
    nand g980(n1632 ,n912 ,n1193);
    or g981(n2659 ,n2620 ,n2647);
    nand g982(n752 ,n204 ,n490);
    nand g983(n1770 ,n1678 ,n1745);
    not g984(n2340 ,n2339);
    nor g985(n2535 ,n2429 ,n2498);
    nand g986(n1159 ,n22[10] ,n463);
    nor g987(n2538 ,n2451 ,n2488);
    or g988(n29[12] ,n3763 ,n3777);
    nand g989(n940 ,n19[4] ,n482);
    nand g990(n3306 ,n3183 ,n3254);
    nand g991(n3508 ,n3459 ,n3485);
    nand g992(n2091 ,n2005 ,n2030);
    nand g993(n146 ,n1878 ,n94);
    dff g994(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1424), .Q(n12[2]));
    nand g995(n2818 ,n28[1] ,n26[0]);
    nand g996(n1572 ,n1001 ,n1230);
    not g997(n2951 ,n2921);
    nor g998(n2465 ,n2406 ,n2417);
    nand g999(n3727 ,n3805 ,n3697);
    dff g1000(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n349), .Q(n25[0]));
    nor g1001(n2519 ,n2427 ,n2480);
    nand g1002(n2694 ,n2684 ,n2693);
    nand g1003(n356 ,n272 ,n314);
    nand g1004(n1347 ,n901 ,n531);
    xor g1005(n3851 ,n3588 ,n3579);
    nand g1006(n3792 ,n3718 ,n3770);
    nand g1007(n889 ,n23[14] ,n447);
    nand g1008(n599 ,n181 ,n483);
    dff g1009(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1528), .Q(n22[6]));
    nand g1010(n871 ,n17[1] ,n468);
    xnor g1011(n239 ,n115 ,n29[8]);
    dff g1012(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1472), .Q(n15[12]));
    nand g1013(n3603 ,n3591 ,n3602);
    dff g1014(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n391), .Q(n26[6]));
    xnor g1015(n2260 ,n2212 ,n2128);
    xnor g1016(n3322 ,n3229 ,n3131);
    nand g1017(n593 ,n180 ,n485);
    nand g1018(n2765 ,n28[3] ,n26[0]);
    not g1019(n2536 ,n2535);
    nand g1020(n1824 ,n29[15] ,n1787);
    or g1021(n3135 ,n3094 ,n3053);
    nand g1022(n2440 ,n2420 ,n2416);
    nand g1023(n2041 ,n3858 ,n1986);
    nand g1024(n720 ,n181 ,n480);
    nand g1025(n1499 ,n1133 ,n738);
    not g1026(n2364 ,n2363);
    nand g1027(n3468 ,n3410 ,n3445);
    nand g1028(n1864 ,n53 ,n52);
    nand g1029(n1630 ,n983 ,n1189);
    nand g1030(n2741 ,n27[1] ,n4[1]);
    nor g1031(n1985 ,n1953 ,n1963);
    or g1032(n1734 ,n1610 ,n1721);
    nand g1033(n1060 ,n16[13] ,n444);
    nor g1034(n2462 ,n2407 ,n2419);
    nand g1035(n1633 ,n1225 ,n1224);
    nor g1036(n2495 ,n2406 ,n2435);
    nand g1037(n1015 ,n19[14] ,n472);
    or g1038(n3319 ,n3240 ,n3270);
    nand g1039(n996 ,n19[2] ,n482);
    nor g1040(n3684 ,n3671 ,n2);
    nand g1041(n1594 ,n1074 ,n879);
    nand g1042(n2396 ,n2395 ,n2374);
    nand g1043(n431 ,n335 ,n384);
    nand g1044(n1116 ,n15[6] ,n443);
    nand g1045(n2081 ,n1978 ,n2032);
    nand g1046(n161 ,n24[3] ,n94);
    nand g1047(n1613 ,n1015 ,n1008);
    nor g1048(n2587 ,n2507 ,n2551);
    or g1049(n3496 ,n3424 ,n3482);
    dff g1050(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1494), .Q(n14[15]));
    dff g1051(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1479), .Q(n8[6]));
    nand g1052(n3759 ,n3838 ,n3685);
    nand g1053(n1809 ,n103 ,n1770);
    nand g1054(n1473 ,n1101 ,n717);
    nand g1055(n542 ,n182 ,n449);
    nand g1056(n887 ,n9[1] ,n496);
    nor g1057(n2567 ,n2486 ,n2539);
    nand g1058(n1262 ,n15[7] ,n493);
    nand g1059(n929 ,n13[6] ,n448);
    nand g1060(n1615 ,n1204 ,n1205);
    nand g1061(n1009 ,n12[2] ,n486);
    nand g1062(n2691 ,n2672 ,n2690);
    nand g1063(n3466 ,n3399 ,n3442);
    nand g1064(n152 ,n24[1] ,n94);
    nand g1065(n1203 ,n23[4] ,n465);
    nor g1066(n799 ,n14[3] ,n467);
    nor g1067(n1316 ,n840 ,n789);
    nor g1068(n2219 ,n2138 ,n2180);
    not g1069(n2709 ,n4[4]);
    nand g1070(n1634 ,n947 ,n1226);
    nand g1071(n717 ,n190 ,n488);
    nand g1072(n1269 ,n18[1] ,n456);
    nor g1073(n2515 ,n2459 ,n2479);
    nand g1074(n2435 ,n2421 ,n2412);
    nand g1075(n2756 ,n27[2] ,n4[7]);
    nand g1076(n679 ,n181 ,n442);
    nand g1077(n2030 ,n3853 ,n1985);
    or g1078(n3070 ,n3012 ,n3002);
    nand g1079(n265 ,n24[5] ,n201);
    nand g1080(n1110 ,n8[6] ,n489);
    or g1081(n2880 ,n2738 ,n2729);
    xnor g1082(n3832 ,n3515 ,n3573);
    nand g1083(n973 ,n9[15] ,n496);
    dff g1084(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1373), .Q(n21[2]));
    nand g1085(n127 ,n29[3] ,n94);
    xnor g1086(n3310 ,n3110 ,n3241);
    not g1087(n95 ,n29[1]);
    nand g1088(n753 ,n191 ,n490);
    nand g1089(n331 ,n26[15] ,n247);
    nor g1090(n2175 ,n2145 ,n2127);
    xnor g1091(n3112 ,n2980 ,n2779);
    nand g1092(n1424 ,n1009 ,n513);
    xnor g1093(n2284 ,n2140 ,n2239);
    nand g1094(n1481 ,n1115 ,n727);
    dff g1095(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1553), .Q(n8[15]));
    nand g1096(n3570 ,n3569 ,n3544);
    nor g1097(n2368 ,n2351 ,n2327);
    not g1098(n2450 ,n2449);
    nand g1099(n3564 ,n3553 ,n3563);
    nand g1100(n895 ,n23[7] ,n447);
    nor g1101(n3429 ,n3372 ,n3401);
    nand g1102(n953 ,n13[0] ,n448);
    dff g1103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1503), .Q(n10[0]));
    nand g1104(n3140 ,n2992 ,n3086);
    nor g1105(n405 ,n27[3] ,n363);
    nand g1106(n3237 ,n3063 ,n3177);
    nand g1107(n1599 ,n883 ,n1087);
    dff g1108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1478), .Q(n15[8]));
    nand g1109(n1771 ,n1681 ,n1756);
    nand g1110(n1114 ,n15[7] ,n443);
    nand g1111(n1515 ,n1151 ,n640);
    nand g1112(n2439 ,n2424 ,n2411);
    xnor g1113(n3830 ,n3549 ,n3569);
    nor g1114(n1715 ,n1706 ,n1705);
    nor g1115(n820 ,n16[9] ,n498);
    nand g1116(n2844 ,n27[3] ,n4[5]);
    not g1117(n2331 ,n2330);
    nand g1118(n1122 ,n15[2] ,n443);
    not g1119(n2707 ,n4[7]);
    dff g1120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1541), .Q(n9[7]));
    nand g1121(n319 ,n121 ,n242);
    dff g1122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1554), .Q(n18[12]));
    nand g1123(n244 ,n29[5] ,n200);
    xor g1124(n1952 ,n1936 ,n1914);
    nor g1125(n801 ,n13[3] ,n500);
    nand g1126(n3473 ,n3433 ,n3454);
    dff g1127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1324), .Q(n17[8]));
    nand g1128(n2769 ,n27[4] ,n4[4]);
    nand g1129(n2046 ,n1931 ,n1998);
    xnor g1130(n3865 ,n3638 ,n3647);
    nand g1131(n1490 ,n1123 ,n690);
    nand g1132(n303 ,n283 ,n248);
    xnor g1133(n30[11] ,n2657 ,n2700);
    nand g1134(n2039 ,n1930 ,n1996);
    xnor g1135(n3127 ,n2988 ,n2769);
    nand g1136(n936 ,n21[2] ,n454);
    nand g1137(n3766 ,n3715 ,n3748);
    nand g1138(n1133 ,n14[12] ,n491);
    nand g1139(n1500 ,n1135 ,n739);
    nor g1140(n2427 ,n2405 ,n2420);
    nand g1141(n510 ,n192 ,n485);
    nand g1142(n1807 ,n29[8] ,n1777);
    nand g1143(n2088 ,n2003 ,n2029);
    nand g1144(n1417 ,n940 ,n608);
    nor g1145(n2481 ,n2406 ,n2444);
    xnor g1146(n1736 ,n1662 ,n29[1]);
    nand g1147(n1218 ,n13[4] ,n501);
    nand g1148(n1228 ,n23[11] ,n465);
    nand g1149(n873 ,n10[1] ,n502);
    or g1150(n2116 ,n2071 ,n2069);
    nand g1151(n1382 ,n948 ,n575);
    nand g1152(n2841 ,n27[1] ,n4[4]);
    or g1153(n1732 ,n1596 ,n1711);
    dff g1154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1507), .Q(n14[6]));
    nand g1155(n1272 ,n23[6] ,n465);
    nand g1156(n2038 ,n1938 ,n2010);
    nor g1157(n2357 ,n2337 ,n2328);
    nor g1158(n2531 ,n2433 ,n2476);
    xnor g1159(n2236 ,n2165 ,n2129);
    nand g1160(n578 ,n191 ,n449);
    nand g1161(n739 ,n204 ,n480);
    nor g1162(n1798 ,n100 ,n1766);
    nand g1163(n1265 ,n11[13] ,n441);
    xnor g1164(n3121 ,n2973 ,n2838);
    xnor g1165(n2540 ,n2500 ,n2468);
    nand g1166(n1134 ,n14[11] ,n491);
    nand g1167(n3512 ,n3469 ,n3494);
    nand g1168(n1195 ,n23[14] ,n465);
    nand g1169(n2915 ,n2737 ,n2732);
    nand g1170(n311 ,n26[9] ,n247);
    or g1171(n2679 ,n2661 ,n2668);
    or g1172(n1839 ,n1825 ,n1831);
    xnor g1173(n2991 ,n2767 ,n2843);
    xnor g1174(n3440 ,n3387 ,n3369);
    nand g1175(n195 ,n123 ,n130);
    xnor g1176(n2215 ,n2158 ,n2119);
    nor g1177(n1312 ,n838 ,n814);
    nand g1178(n1066 ,n13[15] ,n501);
    nand g1179(n1979 ,n3851 ,n1959);
    nor g1180(n1747 ,n1581 ,n1730);
    nor g1181(n1745 ,n1611 ,n1734);
    nand g1182(n3219 ,n2872 ,n3149);
    xnor g1183(n3325 ,n3227 ,n3158);
    nand g1184(n1080 ,n22[14] ,n463);
    nand g1185(n2605 ,n2554 ,n2589);
    xnor g1186(n3104 ,n2956 ,n2768);
    nor g1187(n2482 ,n2408 ,n2439);
    nand g1188(n3696 ,n3864 ,n30[7]);
    xnor g1189(n2976 ,n2738 ,n2729);
    nand g1190(n1408 ,n974 ,n600);
    nand g1191(n1863 ,n51 ,n50);
    or g1192(n1856 ,n1806 ,n1851);
    nand g1193(n3729 ,n30[8] ,n3699);
    nor g1194(n1964 ,n1922 ,n1950);
    nand g1195(n1441 ,n1071 ,n759);
    nand g1196(n1364 ,n924 ,n554);
    nand g1197(n1401 ,n849 ,n611);
    nand g1198(n3579 ,n26[0] ,n4[0]);
    dff g1199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1438), .Q(n8[10]));
    nand g1200(n2339 ,n2282 ,n2306);
    nor g1201(n1806 ,n102 ,n1776);
    nand g1202(n3347 ,n3261 ,n3291);
    dff g1203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1370), .Q(n13[5]));
    nand g1204(n747 ,n178 ,n490);
    nand g1205(n2652 ,n2622 ,n2634);
    xnor g1206(n2207 ,n2097 ,n2151);
    or g1207(n3210 ,n3011 ,n3128);
    nand g1208(n1650 ,n874 ,n1257);
    dff g1209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1848), .Q(n5[14]));
    dff g1210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1535), .Q(n22[2]));
    dff g1211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1351), .Q(n13[13]));
    nand g1212(n1524 ,n1160 ,n647);
    nand g1213(n2778 ,n27[3] ,n4[6]);
    nand g1214(n1378 ,n941 ,n569);
    nand g1215(n559 ,n192 ,n455);
    xnor g1216(n3223 ,n3100 ,n3107);
    nand g1217(n3432 ,n3366 ,n3403);
    nand g1218(n2156 ,n1990 ,n2108);
    dff g1219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n223), .Q(n28[5]));
    nor g1220(n117 ,n28[5] ,n28[7]);
    nand g1221(n3351 ,n3213 ,n3290);
    xnor g1222(n2147 ,n1956 ,n2077);
    not g1223(n97 ,n29[4]);
    xnor g1224(n3312 ,n3160 ,n3238);
    nor g1225(n778 ,n8[9] ,n495);
    nor g1226(n3042 ,n2781 ,n2955);
    not g1227(n3114 ,n3113);
    nand g1228(n872 ,n11[1] ,n478);
    nand g1229(n1177 ,n22[11] ,n463);
    not g1230(n3123 ,n3122);
    nand g1231(n393 ,n311 ,n371);
    nand g1232(n860 ,n12[12] ,n486);
    nand g1233(n534 ,n178 ,n485);
    nand g1234(n2048 ,n3852 ,n2015);
    or g1235(n3333 ,n3190 ,n3300);
    nand g1236(n846 ,n17[6] ,n468);
    nand g1237(n1146 ,n14[4] ,n491);
    xor g1238(n3867 ,n3634 ,n3643);
    or g1239(n1729 ,n1572 ,n1723);
    xnor g1240(n3424 ,n3358 ,n3276);
    nand g1241(n1601 ,n1061 ,n1013);
    nand g1242(n850 ,n17[13] ,n484);
    nand g1243(n2833 ,n27[7] ,n4[3]);
    nand g1244(n1411 ,n981 ,n603);
    nand g1245(n417 ,n5[4] ,n359);
    or g1246(n29[13] ,n3722 ,n3775);
    or g1247(n2395 ,n2375 ,n2394);
    dff g1248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1482), .Q(n8[5]));
    nand g1249(n2837 ,n28[2] ,n26[0]);
    nor g1250(n1302 ,n821 ,n822);
    nand g1251(n3797 ,n3728 ,n3778);
    nand g1252(n3254 ,n3066 ,n3182);
    nand g1253(n270 ,n24[2] ,n201);
    xnor g1254(n2257 ,n2211 ,n2149);
    nor g1255(n762 ,n8[5] ,n495);
    nand g1256(n647 ,n183 ,n450);
    nand g1257(n3200 ,n3083 ,n3102);
    or g1258(n3184 ,n3083 ,n3102);
    xnor g1259(n3388 ,n3351 ,n3327);
    nand g1260(n1614 ,n864 ,n975);
    nand g1261(n657 ,n191 ,n450);
    not g1262(n456 ,n457);
    dff g1263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1322), .Q(n17[10]));
    xnor g1264(n2146 ,n2091 ,n1956);
    xnor g1265(n236 ,n153 ,n29[8]);
    nand g1266(n1359 ,n919 ,n598);
    nand g1267(n715 ,n179 ,n480);
    nor g1268(n131 ,n26[11] ,n26[12]);
    not g1269(n72 ,n71);
    nand g1270(n2500 ,n5[0] ,n2438);
    nand g1271(n1214 ,n12[12] ,n476);
    nor g1272(n3722 ,n3672 ,n3698);
    nand g1273(n1508 ,n1145 ,n747);
    nor g1274(n767 ,n17[2] ,n469);
    nand g1275(n566 ,n187 ,n483);
    not g1276(n2103 ,n2102);
    xnor g1277(n2642 ,n2613 ,n2552);
    nand g1278(n1460 ,n1091 ,n718);
    dff g1279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1537), .Q(n22[0]));
    nand g1280(n1513 ,n1148 ,n750);
    nand g1281(n1659 ,n1272 ,n1271);
    nand g1282(n2168 ,n2154 ,n2123);
    nor g1283(n2217 ,n2137 ,n2167);
    nand g1284(n651 ,n178 ,n450);
    or g1285(n1737 ,n1644 ,n1725);
    nand g1286(n639 ,n179 ,n450);
    nand g1287(n3182 ,n3077 ,n3121);
    nand g1288(n3027 ,n2853 ,n2943);
    nor g1289(n3009 ,n2725 ,n2904);
    nand g1290(n1543 ,n1184 ,n706);
    nand g1291(n751 ,n186 ,n490);
    or g1292(n1746 ,n1281 ,n1739);
    nand g1293(n678 ,n180 ,n442);
    dff g1294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1386), .Q(n20[9]));
    xnor g1295(n2995 ,n2840 ,n2754);
    nand g1296(n423 ,n5[6] ,n359);
    nand g1297(n684 ,n190 ,n442);
    nand g1298(n1501 ,n1134 ,n740);
    xor g1299(n1867 ,n26[15] ,n57);
    nand g1300(n1452 ,n1083 ,n624);
    nor g1301(n807 ,n13[2] ,n500);
    nand g1302(n1379 ,n944 ,n572);
    nand g1303(n673 ,n181 ,n440);
    nor g1304(n248 ,n125 ,n201);
    nand g1305(n1264 ,n13[7] ,n501);
    or g1306(n2191 ,n2154 ,n2123);
    nand g1307(n2942 ,n2741 ,n2792);
    xnor g1308(n3828 ,n3560 ,n3565);
    nand g1309(n2424 ,n3817 ,n4[7]);
    or g1310(n2671 ,n2654 ,n2656);
    nand g1311(n1169 ,n22[4] ,n451);
    nand g1312(n913 ,n21[15] ,n454);
    not g1313(n2848 ,n2847);
    xnor g1314(n240 ,n29[0] ,n116);
    dff g1315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1388), .Q(n20[8]));
    xnor g1316(n2149 ,n2090 ,n1956);
    or g1317(n1845 ,n1820 ,n1835);
    nand g1318(n1077 ,n13[0] ,n501);
    nand g1319(n691 ,n204 ,n440);
    xor g1320(n182 ,n4[11] ,n29[11]);
    xnor g1321(n3592 ,n4[2] ,n26[2]);
    nor g1322(n2552 ,n2471 ,n2537);
    dff g1323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1325), .Q(n17[7]));
    xnor g1324(n3393 ,n3274 ,n3325);
    or g1325(n44 ,n26[8] ,n42);
    xnor g1326(n2958 ,n2746 ,n2717);
    nor g1327(n2346 ,n2292 ,n2343);
    nor g1328(n2274 ,n1895 ,n2245);
    nand g1329(n1637 ,n925 ,n1229);
    nand g1330(n2058 ,n1983 ,n2023);
    xnor g1331(n3841 ,n2367 ,n2383);
    not g1332(n3111 ,n3110);
    nor g1333(n2190 ,n2126 ,n2124);
    dff g1334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1392), .Q(n20[5]));
    nand g1335(n1502 ,n1136 ,n741);
    nand g1336(n892 ,n188 ,n485);
    not g1337(n109 ,n28[1]);
    dff g1338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1501), .Q(n14[11]));
    nor g1339(n1691 ,n1649 ,n1648);
    nand g1340(n902 ,n23[0] ,n447);
    xnor g1341(n1870 ,n26[10] ,n76);
    or g1342(n2883 ,n2836 ,n2714);
    nand g1343(n3052 ,n2901 ,n2998);
    nand g1344(n3217 ,n3048 ,n3150);
    xnor g1345(n3833 ,n3478 ,n3575);
    nand g1346(n1399 ,n990 ,n516);
    xnor g1347(n2542 ,n2502 ,n2466);
    nand g1348(n380 ,n168 ,n289);
    nand g1349(n931 ,n17[11] ,n468);
    xnor g1350(n2137 ,n1955 ,n2075);
    nand g1351(n1838 ,n423 ,n1803);
    or g1352(n2874 ,n2834 ,n2825);
    xnor g1353(n3855 ,n3602 ,n3590);
    nand g1354(n3147 ,n3010 ,n3062);
    nand g1355(n1241 ,n15[10] ,n493);
    nand g1356(n741 ,n185 ,n490);
    nand g1357(n373 ,n281 ,n308);
    not g1358(n464 ,n465);
    not g1359(n2992 ,n2991);
    xnor g1360(n1963 ,n1942 ,n1934);
    nor g1361(n2318 ,n2271 ,n2294);
    or g1362(n1840 ,n1813 ,n1833);
    nand g1363(n2028 ,n3854 ,n1986);
    nor g1364(n2237 ,n2169 ,n2217);
    nand g1365(n1810 ,n104 ,n1771);
    xnor g1366(n3483 ,n3438 ,n3422);
    nor g1367(n1277 ,n793 ,n826);
    nor g1368(n1901 ,n28[1] ,n27[1]);
    not g1369(n458 ,n459);
    nand g1370(n897 ,n23[5] ,n447);
    xnor g1371(n2362 ,n2330 ,n2341);
    nor g1372(n2514 ,n2428 ,n2474);
    xnor g1373(n2280 ,n2244 ,n1895);
    not g1374(n2311 ,n2310);
    or g1375(n1744 ,n1636 ,n1724);
    nor g1376(n2478 ,n2406 ,n2446);
    nand g1377(n1266 ,n18[2] ,n456);
    or g1378(n2870 ,n2800 ,n2832);
    nand g1379(n1710 ,n1316 ,n1315);
    nand g1380(n1635 ,n995 ,n1227);
    nand g1381(n3255 ,n3158 ,n3207);
    nand g1382(n708 ,n187 ,n458);
    nor g1383(n2498 ,n2406 ,n2439);
    xnor g1384(n3132 ,n2995 ,n2946);
    xnor g1385(n2152 ,n2094 ,n1956);
    nand g1386(n1246 ,n18[11] ,n456);
    dff g1387(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1858), .Q(n5[15]));
    nand g1388(n1540 ,n1178 ,n703);
    nand g1389(n334 ,n1873 ,n245);
    xnor g1390(n3270 ,n3167 ,n3104);
    nand g1391(n3203 ,n3127 ,n3115);
    nand g1392(n932 ,n21[4] ,n454);
    nor g1393(n1791 ,n359 ,n1778);
    dff g1394(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1359), .Q(n21[11]));
    nand g1395(n3095 ,n2894 ,n3036);
    nand g1396(n3800 ,n3737 ,n3786);
    nor g1397(n2221 ,n2139 ,n2200);
    dff g1398(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1377), .Q(n20[15]));
    nand g1399(n2635 ,n2567 ,n2609);
    nand g1400(n3195 ,n3074 ,n3103);
    nand g1401(n1977 ,n3855 ,n1958);
    nand g1402(n1478 ,n1113 ,n683);
    not g1403(n484 ,n485);
    nand g1404(n898 ,n23[4] ,n447);
    nand g1405(n742 ,n191 ,n480);
    xnor g1406(n2212 ,n2107 ,n2133);
    nor g1407(n2232 ,n2098 ,n2215);
    nor g1408(n3610 ,n3837 ,n3821);
    or g1409(n2895 ,n2821 ,n2718);
    nand g1410(n2060 ,n1971 ,n2017);
    not g1411(n1897 ,n3855);
    nor g1412(n1934 ,n1909 ,n1913);
    xnor g1413(n3000 ,n2782 ,n2775);
    or g1414(n3179 ,n3057 ,n3104);
    xnor g1415(n1886 ,n26[6] ,n69);
    nor g1416(n2654 ,n2618 ,n2633);
    nand g1417(n275 ,n1865 ,n206);
    or g1418(n3361 ,n3287 ,n3336);
    nand g1419(n332 ,n1889 ,n245);
    nand g1420(n1367 ,n928 ,n556);
    nand g1421(n3500 ,n3457 ,n3484);
    nor g1422(n2316 ,n2240 ,n2298);
    xnor g1423(n3484 ,n3435 ,n3446);
    nand g1424(n1322 ,n855 ,n507);
    dff g1425(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n326), .Q(n24[7]));
    nor g1426(n2492 ,n2405 ,n2443);
    nand g1427(n1521 ,n1156 ,n619);
    nand g1428(n1350 ,n909 ,n538);
    nand g1429(n1358 ,n918 ,n548);
    nand g1430(n2004 ,n3851 ,n1963);
    nand g1431(n2933 ,n2836 ,n2714);
    nor g1432(n3342 ,n3278 ,n3276);
    nand g1433(n1968 ,n3852 ,n1959);
    nor g1434(n1753 ,n1573 ,n1729);
    not g1435(n3514 ,n3505);
    or g1436(n1843 ,n1818 ,n1838);
    nor g1437(n2295 ,n2172 ,n2263);
    xnor g1438(n3268 ,n3164 ,n3126);
    nand g1439(n723 ,n185 ,n480);
    nor g1440(n453 ,n135 ,n416);
    nor g1441(n835 ,n13[8] ,n500);
    nand g1442(n952 ,n20[9] ,n452);
    nand g1443(n904 ,n10[10] ,n502);
    nand g1444(n2793 ,n27[7] ,n4[7]);
    nand g1445(n1432 ,n1027 ,n667);
    nand g1446(n1124 ,n10[4] ,n481);
    nand g1447(n1158 ,n9[12] ,n459);
    nand g1448(n3419 ,n3364 ,n3405);
    nand g1449(n2008 ,n3858 ,n1958);
    xnor g1450(n2983 ,n2807 ,n2814);
    nand g1451(n1636 ,n1228 ,n931);
    nand g1452(n3569 ,n3568 ,n3556);
    xnor g1453(n3128 ,n2987 ,n2827);
    nand g1454(n734 ,n186 ,n480);
    nand g1455(n886 ,n19[11] ,n482);
    not g1456(n138 ,n139);
    not g1457(n448 ,n449);
    nand g1458(n323 ,n256 ,n264);
    nand g1459(n3188 ,n3052 ,n3146);
    nand g1460(n1239 ,n14[10] ,n466);
    nor g1461(n2227 ,n2156 ,n2166);
    nand g1462(n1862 ,n49 ,n48);
    nand g1463(n1466 ,n1098 ,n632);
    xnor g1464(n2979 ,n2781 ,n2792);
    nand g1465(n2803 ,n28[5] ,n26[3]);
    nand g1466(n3691 ,n3866 ,n30[5]);
    nand g1467(n3038 ,n2748 ,n2926);
    dff g1468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1495), .Q(n14[14]));
    nor g1469(n2468 ,n2406 ,n2422);
    dff g1470(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n342), .Q(n24[4]));
    xnor g1471(n30[5] ,n2677 ,n2685);
    nand g1472(n660 ,n180 ,n457);
    nand g1473(n2776 ,n27[0] ,n4[6]);
    dff g1474(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1379), .Q(n20[14]));
    nand g1475(n1533 ,n1169 ,n652);
    nor g1476(n809 ,n21[2] ,n470);
    nand g1477(n3063 ,n2875 ,n3018);
    nand g1478(n2747 ,n27[1] ,n4[7]);
    xnor g1479(n1923 ,n28[5] ,n27[5]);
    nand g1480(n733 ,n179 ,n490);
    dff g1481(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1442), .Q(n16[15]));
    nor g1482(n1296 ,n769 ,n825);
    nand g1483(n1978 ,n3851 ,n1958);
    dff g1484(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n324), .Q(n25[4]));
    nand g1485(n561 ,n187 ,n455);
    or g1486(n2189 ,n2133 ,n2128);
    nor g1487(n2556 ,n2465 ,n2536);
    nand g1488(n420 ,n5[8] ,n359);
    dff g1489(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1473), .Q(n8[7]));
    nand g1490(n1876 ,n43 ,n42);
    nor g1491(n321 ,n133 ,n251);
    nand g1492(n731 ,n192 ,n488);
    nor g1493(n3614 ,n3844 ,n3828);
    or g1494(n2684 ,n2658 ,n2667);
    nand g1495(n1013 ,n8[15] ,n494);
    nor g1496(n2905 ,n2846 ,n2858);
    dff g1497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1425), .Q(n12[3]));
    not g1498(n84 ,n83);
    nand g1499(n1181 ,n8[1] ,n489);
    nor g1500(n826 ,n13[5] ,n500);
    xor g1501(n1953 ,n1935 ,n1924);
    nand g1502(n858 ,n17[4] ,n468);
    dff g1503(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1428), .Q(n12[0]));
    xnor g1504(n3831 ,n3540 ,n3571);
    nor g1505(n3858 ,n3577 ,n3607);
    dff g1506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1489), .Q(n15[2]));
    nand g1507(n1090 ,n16[5] ,n444);
    nand g1508(n3427 ,n3416 ,n3395);
    xnor g1509(n2138 ,n2065 ,n1957);
    not g1510(n99 ,n29[0]);
    nand g1511(n955 ,n20[7] ,n452);
    nor g1512(n3074 ,n2882 ,n3020);
    nor g1513(n1759 ,n1653 ,n1738);
    xnor g1514(n30[9] ,n2688 ,n2696);
    xnor g1515(n386 ,n113 ,n284);
    nand g1516(n1104 ,n15[13] ,n443);
    xnor g1517(n3826 ,n3550 ,n3561);
    nand g1518(n3247 ,n3064 ,n3200);
    nand g1519(n2604 ,n2559 ,n2403);
    nor g1520(n2479 ,n2405 ,n2446);
    nand g1521(n635 ,n184 ,n457);
    nand g1522(n1174 ,n22[0] ,n451);
    xnor g1523(n2155 ,n2095 ,n1956);
    nand g1524(n2943 ,n2738 ,n2729);
    xnor g1525(n238 ,n155 ,n29[12]);
    or g1526(n3363 ,n3351 ,n3327);
    not g1527(n2501 ,n2500);
    nand g1528(n987 ,n9[12] ,n496);
    nor g1529(n3350 ,n3197 ,n3308);
    nand g1530(n340 ,n26[13] ,n247);
    not g1531(n2178 ,n2171);
    nand g1532(n2742 ,n28[0] ,n26[7]);
    xnor g1533(n3271 ,n3162 ,n3121);
    nand g1534(n3138 ,n2991 ,n3087);
    nand g1535(n1204 ,n20[13] ,n461);
    nand g1536(n3713 ,n30[10] ,n3699);
    nand g1537(n479 ,n207 ,n405);
    nand g1538(n851 ,n17[12] ,n484);
    not g1539(n3087 ,n3086);
    nand g1540(n1250 ,n18[8] ,n456);
    nand g1541(n1206 ,n23[13] ,n465);
    xnor g1542(n2330 ,n2234 ,n2279);
    nand g1543(n888 ,n23[15] ,n447);
    nand g1544(n2547 ,n2487 ,n2522);
    not g1545(n2761 ,n2710);
    dff g1546(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n228), .Q(n27[7]));
    nand g1547(n2800 ,n28[1] ,n26[4]);
    nor g1548(n3649 ,n3613 ,n3648);
    nand g1549(n1018 ,n10[6] ,n502);
    xnor g1550(n3856 ,n3586 ,n3604);
    xnor g1551(n3003 ,n2758 ,n2755);
    nor g1552(n2167 ,n2101 ,n2150);
    or g1553(n52 ,n26[12] ,n50);
    xnor g1554(n2668 ,n2644 ,n2622);
    nand g1555(n3698 ,n2 ,n3);
    nand g1556(n434 ,n5[7] ,n359);
    nand g1557(n1426 ,n962 ,n589);
    nor g1558(n1299 ,n823 ,n824);
    xnor g1559(n3230 ,n3116 ,n3129);
    nor g1560(n3678 ,n3861 ,n30[10]);
    xnor g1561(n3435 ,n3409 ,n3400);
    nand g1562(n1185 ,n9[4] ,n459);
    nand g1563(n160 ,n1876 ,n94);
    not g1564(n172 ,n171);
    dff g1565(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1455), .Q(n10[15]));
    nor g1566(n2521 ,n2458 ,n2493);
    nor g1567(n796 ,n23[5] ,n464);
    nand g1568(n2810 ,n28[4] ,n26[2]);
    xnor g1569(n2205 ,n2139 ,n2146);
    nand g1570(n2317 ,n2260 ,n2284);
    xnor g1571(n1916 ,n28[4] ,n27[4]);
    nand g1572(n1414 ,n963 ,n592);
    nand g1573(n1589 ,n1059 ,n1138);
    xnor g1574(n3122 ,n2964 ,n2759);
    nand g1575(n1212 ,n22[13] ,n463);
    nand g1576(n1240 ,n18[14] ,n456);
    not g1577(n2857 ,n2856);
    xor g1578(n2403 ,n2516 ,n2506);
    nand g1579(n3078 ,n2874 ,n3038);
    nand g1580(n1576 ,n1031 ,n992);
    not g1581(n2177 ,n1895);
    nor g1582(n793 ,n15[5] ,n492);
    nor g1583(n2507 ,n2467 ,n2502);
    nand g1584(n2909 ,n2713 ,n2822);
    nand g1585(n3719 ,n30[7] ,n3699);
    dff g1586(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1847), .Q(n5[10]));
    nand g1587(n3024 ,n2935 ,n2906);
    or g1588(n2866 ,n2713 ,n2822);
    nand g1589(n3669 ,n3618 ,n3668);
    xnor g1590(n2235 ,n2163 ,n2157);
    or g1591(n3235 ,n3114 ,n3185);
    nor g1592(n504 ,n128 ,n392);
    nand g1593(n2746 ,n28[6] ,n26[4]);
    dff g1594(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1556), .Q(n18[10]));
    nor g1595(n2393 ,n2392 ,n2378);
    nor g1596(n487 ,n140 ,n416);
    or g1597(n3553 ,n3535 ,n2705);
    or g1598(n2888 ,n2746 ,n2717);
    nand g1599(n2821 ,n28[0] ,n26[6]);
    nand g1600(n666 ,n178 ,n440);
    or g1601(n2486 ,n2407 ,n2440);
    nand g1602(n3556 ,n3536 ,n3542);
    nor g1603(n781 ,n17[5] ,n469);
    nor g1604(n2512 ,n2426 ,n2475);
    nor g1605(n825 ,n15[2] ,n492);
    dff g1606(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1550), .Q(n18[15]));
    nand g1607(n3522 ,n3502 ,n3507);
    nand g1608(n1423 ,n1002 ,n543);
    nand g1609(n941 ,n13[3] ,n448);
    nor g1610(n1973 ,n1897 ,n1961);
    nand g1611(n1493 ,n1127 ,n732);
    nand g1612(n469 ,n209 ,n413);
    xnor g1613(n2574 ,n2513 ,n2529);
    nor g1614(n1666 ,n1583 ,n1582);
    nor g1615(n2197 ,n2119 ,n2158);
    nand g1616(n3474 ,n3415 ,n3451);
    xnor g1617(n2960 ,n2811 ,n2716);
    nand g1618(n2026 ,n3855 ,n1985);
    nor g1619(n3304 ,n3174 ,n3251);
    dff g1620(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1326), .Q(n17[6]));
    xnor g1621(n3422 ,n3356 ,n3307);
    xor g1622(n1958 ,n1944 ,n1948);
    nand g1623(n572 ,n188 ,n453);
    xnor g1624(n2326 ,n2280 ,n2264);
    nand g1625(n313 ,n26[6] ,n247);
    nor g1626(n2464 ,n2405 ,n2423);
    nand g1627(n2779 ,n27[0] ,n4[7]);
    xnor g1628(n2344 ,n2310 ,n2242);
    nor g1629(n786 ,n10[9] ,n503);
    nand g1630(n1028 ,n18[15] ,n474);
    not g1631(n2612 ,n2611);
    nor g1632(n1692 ,n1651 ,n1650);
    nand g1633(n350 ,n268 ,n299);
    nor g1634(n1819 ,n97 ,n1782);
    nand g1635(n1557 ,n1244 ,n756);
    nand g1636(n252 ,n29[12] ,n202);
    nand g1637(n935 ,n19[9] ,n482);
    dff g1638(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1368), .Q(n21[5]));
    xnor g1639(n3638 ,n3838 ,n3822);
    or g1640(n46 ,n26[9] ,n44);
    nand g1641(n864 ,n19[13] ,n472);
    nor g1642(n3653 ,n3621 ,n3652);
    nand g1643(n1113 ,n15[8] ,n443);
    xnor g1644(n192 ,n97 ,n4[4]);
    nand g1645(n205 ,n94 ,n172);
    nand g1646(n473 ,n207 ,n413);
    nor g1647(n2247 ,n2194 ,n2222);
    nand g1648(n1803 ,n98 ,n1761);
    nand g1649(n2690 ,n2670 ,n2689);
    nand g1650(n2341 ,n2267 ,n2314);
    nand g1651(n1854 ,n419 ,n1814);
    nand g1652(n1772 ,n1684 ,n1754);
    nor g1653(n74 ,n59 ,n73);
    nand g1654(n1522 ,n1158 ,n698);
    nor g1655(n2218 ,n2134 ,n2178);
    nand g1656(n282 ,n25[7] ,n203);
    not g1657(n470 ,n471);
    xnor g1658(n2141 ,n2074 ,n2072);
    not g1659(n96 ,n29[7]);
    nand g1660(n637 ,n181 ,n457);
    xnor g1661(n3822 ,n3465 ,n3433);
    nand g1662(n3535 ,n3499 ,n3523);
    xnor g1663(n186 ,n100 ,n4[2]);
    dff g1664(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1513), .Q(n14[3]));
    xnor g1665(n3159 ,n2960 ,n3000);
    nand g1666(n1156 ,n22[11] ,n451);
    or g1667(n1857 ,n1796 ,n1853);
    nor g1668(n3683 ,n3860 ,n30[11]);
    or g1669(n1841 ,n1816 ,n1836);
    nand g1670(n985 ,n19[12] ,n472);
    dff g1671(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1320), .Q(n17[12]));
    dff g1672(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1444), .Q(n11[3]));
    xnor g1673(n2303 ,n2237 ,n2261);
    nor g1674(n2484 ,n2408 ,n2443);
    nand g1675(n1935 ,n1915 ,n1918);
    nand g1676(n687 ,n192 ,n442);
    nand g1677(n1837 ,n434 ,n1802);
    not g1678(n2839 ,n2838);
    nor g1679(n284 ,n29[0] ,n247);
    nand g1680(n2794 ,n28[5] ,n26[6]);
    nand g1681(n925 ,n11[11] ,n478);
    nand g1682(n2586 ,n2508 ,n2549);
    nand g1683(n1217 ,n13[12] ,n501);
    nor g1684(n3705 ,n3698 ,n3679);
    nand g1685(n627 ,n178 ,n445);
    not g1686(n2706 ,n27[3]);
    dff g1687(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1504), .Q(n14[9]));
    nor g1688(n3524 ,n3504 ,n3503);
    not g1689(n3287 ,n3286);
    nand g1690(n2002 ,n3856 ,n1963);
    nand g1691(n443 ,n139 ,n407);
    dff g1692(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1469), .Q(n21[3]));
    nor g1693(n1288 ,n801 ,n792);
    xnor g1694(n2968 ,n2712 ,n2824);
    nand g1695(n1413 ,n1019 ,n604);
    nand g1696(n644 ,n188 ,n457);
    xnor g1697(n3825 ,n3541 ,n3548);
    not g1698(n1765 ,n1764);
    not g1699(n2842 ,n2841);
    nor g1700(n1663 ,n1575 ,n1574);
    nand g1701(n2174 ,n2145 ,n2127);
    dff g1702(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1411), .Q(n19[8]));
    xnor g1703(n2208 ,n1956 ,n2134);
    nand g1704(n3050 ,n2947 ,n2995);
    nand g1705(n921 ,n21[10] ,n454);
    nand g1706(n354 ,n273 ,n341);
    nand g1707(n1390 ,n956 ,n582);
    dff g1708(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1412), .Q(n19[7]));
    xnor g1709(n2625 ,n2594 ,n2592);
    or g1710(n3180 ,n3108 ,n3106);
    dff g1711(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1382), .Q(n20[12]));
    xor g1712(n3161 ,n2990 ,n2844);
    nand g1713(n718 ,n188 ,n480);
    nand g1714(n2662 ,n2626 ,n2652);
    nand g1715(n3758 ,n3849 ,n3685);
    nor g1716(n776 ,n19[9] ,n473);
    nor g1717(n2499 ,n2408 ,n2444);
    or g1718(n391 ,n286 ,n346);
    dff g1719(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1348), .Q(n23[0]));
    nand g1720(n3433 ,n3383 ,n3406);
    nand g1721(n3236 ,n3110 ,n3189);
    nand g1722(n1058 ,n11[2] ,n441);
    nor g1723(n2229 ,n2144 ,n2196);
    nand g1724(n3413 ,n3315 ,n3377);
    nand g1725(n1723 ,n1695 ,n1694);
    nand g1726(n164 ,n1892 ,n94);
    nand g1727(n3430 ,n3409 ,n3400);
    nand g1728(n3566 ,n3565 ,n3551);
    not g1729(n498 ,n499);
    nand g1730(n2739 ,n27[2] ,n4[2]);
    nand g1731(n3407 ,n3316 ,n3378);
    nand g1732(n856 ,n11[7] ,n478);
    nand g1733(n326 ,n250 ,n263);
    nand g1734(n1720 ,n1674 ,n1673);
    nand g1735(n310 ,n1870 ,n245);
    nor g1736(n67 ,n58 ,n66);
    nand g1737(n2703 ,n27[0] ,n4[1]);
    dff g1738(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1391), .Q(n20[6]));
    xnor g1739(n1955 ,n1941 ,n1923);
    nand g1740(n1609 ,n1080 ,n1068);
    nor g1741(n2170 ,n1956 ,n2131);
    nor g1742(n3374 ,n3305 ,n3338);
    nor g1743(n207 ,n27[2] ,n175);
    nor g1744(n2113 ,n2068 ,n2067);
    not g1745(n3594 ,n3593);
    or g1746(n3554 ,n3536 ,n3542);
    nand g1747(n418 ,n5[10] ,n359);
    nand g1748(n2183 ,n2146 ,n2132);
    dff g1749(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1403), .Q(n19[14]));
    nand g1750(n3717 ,n3831 ,n3684);
    nand g1751(n3344 ,n3101 ,n3285);
    xnor g1752(n1888 ,n26[4] ,n66);
    nor g1753(n2879 ,n2719 ,n2819);
    dff g1754(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n13[8]));
    not g1755(n494 ,n495);
    nand g1756(n1595 ,n1075 ,n880);
    nand g1757(n928 ,n21[6] ,n454);
    dff g1758(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1319), .Q(n17[13]));
    nand g1759(n1462 ,n1094 ,n719);
    nand g1760(n1274 ,n23[9] ,n447);
    nand g1761(n1409 ,n935 ,n610);
    nand g1762(n1253 ,n18[6] ,n456);
    dff g1763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1331), .Q(n17[1]));
    nor g1764(n787 ,n10[2] ,n503);
    nor g1765(n1684 ,n1629 ,n1628);
    nand g1766(n1357 ,n916 ,n546);
    nand g1767(n1647 ,n1241 ,n903);
    or g1768(n2673 ,n2632 ,n2664);
    nand g1769(n1829 ,n421 ,n1810);
    nor g1770(n3457 ,n3360 ,n3429);
    dff g1771(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1418), .Q(n19[3]));
    not g1772(n3589 ,n3588);
    xnor g1773(n3107 ,n2957 ,n2732);
    or g1774(n1306 ,n776 ,n785);
    not g1775(n3080 ,n3079);
    nand g1776(n1430 ,n1025 ,n710);
    nand g1777(n2855 ,n28[2] ,n26[1]);
    nand g1778(n603 ,n184 ,n483);
    nand g1779(n1334 ,n889 ,n520);
    nand g1780(n3539 ,n3500 ,n3529);
    nand g1781(n1086 ,n10[15] ,n481);
    not g1782(n104 ,n29[13]);
    nand g1783(n2057 ,n3857 ,n1986);
    nand g1784(n1530 ,n1168 ,n651);
    nand g1785(n1646 ,n1006 ,n904);
    dff g1786(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n422), .Q(n26[14]));
    nand g1787(n2095 ,n2012 ,n2056);
    nor g1788(n1813 ,n29[3] ,n1783);
    nor g1789(n840 ,n16[8] ,n498);
    dff g1790(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1446), .Q(n16[13]));
    xnor g1791(n2345 ,n2312 ,n2277);
    nand g1792(n83 ,n26[13] ,n81);
    dff g1793(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1352), .Q(n13[12]));
    nor g1794(n1310 ,n836 ,n775);
    xnor g1795(n2328 ,n2276 ,n2259);
    xnor g1796(n3100 ,n2967 ,n2773);
    nand g1797(n2111 ,n1954 ,n2076);
    nand g1798(n2722 ,n28[5] ,n26[7]);
    nand g1799(n1631 ,n991 ,n943);
    nand g1800(n1184 ,n9[5] ,n459);
    nand g1801(n1938 ,n3858 ,n1922);
    nand g1802(n1797 ,n29[3] ,n1769);
    nand g1803(n2795 ,n27[7] ,n4[6]);
    nand g1804(n683 ,n184 ,n442);
    nand g1805(n2661 ,n2630 ,n2645);
    nand g1806(n395 ,n5[1] ,n359);
    nor g1807(n1990 ,n1946 ,n1962);
    dff g1808(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1339), .Q(n23[9]));
    xnor g1809(n30[8] ,n2687 ,n2694);
    xnor g1810(n231 ,n145 ,n29[0]);
    nand g1811(n2832 ,n27[2] ,n4[3]);
    nand g1812(n1483 ,n1116 ,n685);
    nand g1813(n2374 ,n2359 ,n2370);
    nand g1814(n3410 ,n3340 ,n3384);
    dff g1815(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n216), .Q(n28[6]));
    nor g1816(n2194 ,n2073 ,n2152);
    dff g1817(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n233), .Q(n28[2]));
    nand g1818(n3072 ,n2830 ,n2999);
    xnor g1819(n2135 ,n2082 ,n1957);
    or g1820(n2415 ,n3811 ,n4[1]);
    nand g1821(n881 ,n17[6] ,n484);
    nand g1822(n3665 ,n3619 ,n3664);
    nor g1823(n2114 ,n1945 ,n2067);
    nand g1824(n3256 ,n3114 ,n3185);
    nand g1825(n3574 ,n3506 ,n3573);
    nand g1826(n3202 ,n3108 ,n3106);
    dff g1827(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n431), .Q(n26[12]));
    or g1828(n1858 ,n1808 ,n1852);
    nor g1829(n2865 ,n2741 ,n2792);
    nor g1830(n2383 ,n2333 ,n2373);
    xnor g1831(n3842 ,n2361 ,n2385);
    nand g1832(n1471 ,n1107 ,n724);
    nand g1833(n3294 ,n3208 ,n3242);
    nand g1834(n3456 ,n3398 ,n3421);
    nand g1835(n2084 ,n2013 ,n2024);
    xnor g1836(n3864 ,n3640 ,n3649);
    or g1837(n128 ,n26[0] ,n26[1]);
    nand g1838(n1547 ,n1194 ,n755);
    xnor g1839(n221 ,n114 ,n29[2]);
    dff g1840(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1502), .Q(n14[10]));
    nand g1841(n1089 ,n8[8] ,n489);
    nand g1842(n616 ,n181 ,n485);
    or g1843(n3315 ,n3101 ,n3285);
    nand g1844(n632 ,n191 ,n445);
    xnor g1845(n2590 ,n2540 ,n2521);
    not g1846(n2796 ,n2795);
    nand g1847(n524 ,n183 ,n446);
    nand g1848(n713 ,n180 ,n440);
    or g1849(n31 ,n26[1] ,n26[0]);
    nand g1850(n3337 ,n3238 ,n3272);
    nor g1851(n811 ,n22[2] ,n462);
    nand g1852(n965 ,n20[3] ,n452);
    nor g1853(n116 ,n27[0] ,n1);
    nand g1854(n1929 ,n3856 ,n1922);
    nor g1855(n765 ,n11[3] ,n479);
    nand g1856(n1832 ,n417 ,n1799);
    nand g1857(n571 ,n186 ,n449);
    nand g1858(n3010 ,n2797 ,n2949);
    nand g1859(n3617 ,n3847 ,n3831);
    xnor g1860(n2158 ,n1956 ,n2092);
    xnor g1861(n2139 ,n1957 ,n2078);
    nand g1862(n251 ,n117 ,n197);
    nand g1863(n3732 ,n3832 ,n3684);
    nand g1864(n1123 ,n15[1] ,n443);
    nor g1865(n1987 ,n1952 ,n1959);
    or g1866(n2891 ,n2815 ,n2715);
    not g1867(n322 ,n317);
    nor g1868(n837 ,n22[8] ,n462);
    not g1869(n70 ,n69);
    nand g1870(n3716 ,n3828 ,n3684);
    xnor g1871(n2988 ,n2714 ,n2836);
    nand g1872(n700 ,n187 ,n440);
    nand g1873(n3394 ,n3288 ,n3375);
    nand g1874(n2910 ,n2799 ,n2731);
    xnor g1875(n1874 ,n26[14] ,n83);
    nand g1876(n1100 ,n10[11] ,n481);
    nand g1877(n1373 ,n936 ,n563);
    nand g1878(n1582 ,n1038 ,n966);
    nand g1879(n1372 ,n1102 ,n677);
    or g1880(n3193 ,n3060 ,n3126);
    nand g1881(n1850 ,n432 ,n1822);
    nand g1882(n2293 ,n2235 ,n2256);
    nand g1883(n3645 ,n3620 ,n3644);
    nor g1884(n822 ,n12[9] ,n477);
    nor g1885(n122 ,n29[1] ,n1884);
    nand g1886(n353 ,n257 ,n316);
    xnor g1887(n3355 ,n3273 ,n3187);
    nand g1888(n686 ,n178 ,n442);
    nand g1889(n278 ,n1867 ,n206);
    or g1890(n29[8] ,n3781 ,n3802);
    nand g1891(n1939 ,n1907 ,n1920);
    nor g1892(n3335 ,n3187 ,n3273);
    nand g1893(n1775 ,n1690 ,n1760);
    or g1894(n2267 ,n2233 ,n2236);
    dff g1895(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1845), .Q(n5[0]));
    or g1896(n2881 ,n2835 ,n2803);
    or g1897(n2894 ,n2721 ,n2790);
    nand g1898(n2715 ,n28[5] ,n26[2]);
    nand g1899(n170 ,n29[1] ,n1891);
    nand g1900(n550 ,n204 ,n483);
    nand g1901(n2944 ,n2824 ,n2712);
    nand g1902(n3013 ,n2785 ,n2915);
    nand g1903(n976 ,n8[13] ,n494);
    nand g1904(n3145 ,n3067 ,n3050);
    nor g1905(n1899 ,n28[5] ,n27[5]);
    nand g1906(n1154 ,n22[12] ,n451);
    or g1907(n2410 ,n3815 ,n4[5]);
    nor g1908(n2143 ,n1989 ,n2103);
    nand g1909(n3317 ,n3281 ,n3268);
    nor g1910(n804 ,n21[3] ,n470);
    dff g1911(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n437), .Q(n26[4]));
    or g1912(n3506 ,n3441 ,n3490);
    not g1913(n3776 ,n3764);
    nand g1914(n1323 ,n982 ,n605);
    nand g1915(n53 ,n26[12] ,n50);
    xnor g1916(n1912 ,n28[1] ,n27[1]);
    nor g1917(n457 ,n135 ,n409);
    nand g1918(n1271 ,n20[6] ,n461);
    not g1919(n2862 ,n2861);
    xnor g1920(n3238 ,n3132 ,n3067);
    nand g1921(n962 ,n12[13] ,n486);
    nand g1922(n2782 ,n28[3] ,n26[1]);
    not g1923(n1954 ,n1955);
    nand g1924(n3715 ,n3824 ,n3684);
    not g1925(n3082 ,n3081);
    nand g1926(n3371 ,n3262 ,n3318);
    nor g1927(n1311 ,n837 ,n815);
    xnor g1928(n2133 ,n2063 ,n1957);
    nand g1929(n754 ,n204 ,n488);
    nand g1930(n3746 ,n3847 ,n3685);
    nor g1931(n2428 ,n2408 ,n2423);
    nand g1932(n2017 ,n3852 ,n1986);
    nand g1933(n2768 ,n27[0] ,n4[5]);
    nand g1934(n3764 ,n3744 ,n3726);
    xnor g1935(n3274 ,n3166 ,n3102);
    nand g1936(n3583 ,n26[5] ,n4[5]);
    nand g1937(n2018 ,n3855 ,n1987);
    nand g1938(n2089 ,n2002 ,n2026);
    dff g1939(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1413), .Q(n12[7]));
    nand g1940(n519 ,n179 ,n446);
    or g1941(n3450 ,n3411 ,n3423);
    or g1942(n2558 ,n2509 ,n2527);
    or g1943(n1281 ,n797 ,n829);
    nand g1944(n1140 ,n10[0] ,n481);
    nand g1945(n3262 ,n3143 ,n3176);
    or g1946(n3597 ,n3592 ,n3596);
    nor g1947(n3251 ,n3129 ,n3220);
    nand g1948(n1025 ,n11[11] ,n441);
    nor g1949(n404 ,n27[3] ,n366);
    nand g1950(n1388 ,n954 ,n581);
    nand g1951(n901 ,n23[1] ,n447);
    nand g1952(n3303 ,n3199 ,n3255);
    dff g1953(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1490), .Q(n15[1]));
    nand g1954(n1391 ,n957 ,n584);
    nor g1955(n298 ,n122 ,n249);
    nand g1956(n3573 ,n3538 ,n3572);
    nand g1957(n2629 ,n2591 ,n2607);
    nor g1958(n2474 ,n2405 ,n2442);
    xnor g1959(n2576 ,n2527 ,n2509);
    nand g1960(n1558 ,n1249 ,n661);
    nand g1961(n1906 ,n28[6] ,n28[5]);
    nand g1962(n3477 ,n3432 ,n3439);
    nand g1963(n1033 ,n21[4] ,n471);
    not g1964(n2851 ,n2850);
    nand g1965(n1981 ,n3854 ,n1958);
    nand g1966(n3431 ,n3382 ,n3394);
    nor g1967(n841 ,n20[5] ,n460);
    nand g1968(n2843 ,n28[7] ,n26[0]);
    or g1969(n2636 ,n2581 ,n2614);
    nor g1970(n795 ,n14[5] ,n467);
    nor g1971(n142 ,n27[1] ,n27[6]);
    xnor g1972(n3593 ,n4[3] ,n26[3]);
    nor g1973(n1891 ,n63 ,n61);
    nand g1974(n2417 ,n3816 ,n4[6]);
    nor g1975(n2494 ,n2405 ,n2440);
    nand g1976(n80 ,n26[11] ,n79);
    nand g1977(n1620 ,n978 ,n1211);
    nor g1978(n3248 ,n3154 ,n3186);
    nand g1979(n1767 ,n1669 ,n1750);
    not g1980(n3308 ,n3294);
    dff g1981(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1567), .Q(n11[12]));
    not g1982(n444 ,n445);
    xor g1983(n3814 ,n28[4] ,n27[4]);
    nand g1984(n1402 ,n969 ,n595);
    nand g1985(n1164 ,n22[8] ,n451);
    nand g1986(n3581 ,n26[3] ,n4[3]);
    nand g1987(n363 ,n27[0] ,n320);
    dff g1988(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1464), .Q(n16[1]));
    dff g1989(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1497), .Q(n10[2]));
    nand g1990(n2826 ,n28[1] ,n26[6]);
    nand g1991(n697 ,n191 ,n458);
    nand g1992(n625 ,n190 ,n445);
    nand g1993(n946 ,n20[13] ,n452);
    dff g1994(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1451), .Q(n16[9]));
    nand g1995(n848 ,n17[14] ,n484);
    not g1996(n200 ,n201);
    nand g1997(n3795 ,n3713 ,n3762);
    nor g1998(n771 ,n8[8] ,n495);
    or g1999(n38 ,n26[5] ,n36);
    nor g2000(n2533 ,n2452 ,n2482);
    nand g2001(n1805 ,n101 ,n1775);
    dff g2002(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n237), .Q(n27[4]));
    nand g2003(n398 ,n5[14] ,n359);
    dff g2004(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n323), .Q(n24[6]));
    nand g2005(n1193 ,n21[15] ,n471);
    nand g2006(n870 ,n8[1] ,n494);
    dff g2007(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n377), .Q(n25[2]));
    xor g2008(n3313 ,n3190 ,n3263);
    not g2009(n2408 ,n5[1]);
    nand g2010(n2840 ,n28[5] ,n26[1]);
    nand g2011(n3043 ,n2780 ,n2914);
    nor g2012(n1812 ,n103 ,n1788);
    nand g2013(n3561 ,n3531 ,n3557);
    dff g2014(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1437), .Q(n11[6]));
    nand g2015(n721 ,n189 ,n488);
    nand g2016(n1049 ,n11[4] ,n441);
    xnor g2017(n3840 ,n2344 ,n2371);
    xnor g2018(n3225 ,n2733 ,n3128);
    nor g2019(n1309 ,n835 ,n834);
    nand g2020(n1433 ,n1029 ,n712);
    nand g2021(n1561 ,n1253 ,n663);
    dff g2022(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1521), .Q(n22[11]));
    nand g2023(n1001 ,n19[6] ,n472);
    not g2024(n2101 ,n2100);
    nand g2025(n2916 ,n2721 ,n2790);
    nand g2026(n947 ,n10[11] ,n502);
    nand g2027(n33 ,n26[2] ,n31);
    xnor g2028(n1871 ,n26[11] ,n78);
    nand g2029(n477 ,n212 ,n404);
    nand g2030(n729 ,n178 ,n480);
    nand g2031(n2419 ,n3811 ,n4[1]);
    xnor g2032(n2665 ,n2620 ,n2647);
    nand g2033(n1172 ,n9[10] ,n459);
    dff g2034(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1318), .Q(n17[14]));
    nor g2035(n775 ,n17[8] ,n469);
    nand g2036(n2824 ,n28[3] ,n26[4]);
    xnor g2037(n3129 ,n2969 ,n2776);
    nand g2038(n2931 ,n2722 ,n2820);
    nand g2039(n1507 ,n1143 ,n745);
    not g2040(n176 ,n175);
    nand g2041(n3093 ,n2876 ,n3029);
    nand g2042(n1199 ,n20[4] ,n461);
    xnor g2043(n2596 ,n2542 ,n2517);
    dff g2044(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1481), .Q(n10[7]));
    nand g2045(n3768 ,n3695 ,n3704);
    not g2046(n134 ,n135);
    dff g2047(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n224), .Q(n27[6]));
    nor g2048(n1304 ,n831 ,n819);
    not g2049(n413 ,n412);
    nand g2050(n1052 ,n16[1] ,n499);
    xnor g2051(n2361 ,n2332 ,n2318);
    nand g2052(n1007 ,n9[13] ,n496);
    nand g2053(n3411 ,n3349 ,n3376);
    nor g2054(n2461 ,n2407 ,n2418);
    xnor g2055(n2370 ,n2323 ,n2301);
    or g2056(n1762 ,n1698 ,n1746);
    nand g2057(n1237 ,n23[10] ,n465);
    nand g2058(n2864 ,n28[0] ,n26[0]);
    nand g2059(n521 ,n181 ,n446);
    xnor g2060(n2580 ,n2486 ,n2539);
    nand g2061(n2583 ,n2566 ,n2402);
    nand g2062(n596 ,n204 ,n453);
    nand g2063(n1628 ,n987 ,n986);
    nand g2064(n56 ,n26[13] ,n52);
    nand g2065(n400 ,n336 ,n372);
    nand g2066(n547 ,n180 ,n455);
    xnor g2067(n3097 ,n3002 ,n2805);
    not g2068(n406 ,n405);
    nand g2069(n309 ,n1871 ,n245);
    nor g2070(n2431 ,n2407 ,n2422);
    xor g2071(n1951 ,n1937 ,n1923);
    nand g2072(n2016 ,n3850 ,n1987);
    nand g2073(n1970 ,n3856 ,n1959);
    nand g2074(n258 ,n25[6] ,n203);
    nor g2075(n119 ,n29[4] ,n1888);
    nand g2076(n2927 ,n2811 ,n2716);
    dff g2077(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1461), .Q(n16[3]));
    dff g2078(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1395), .Q(n20[3]));
    nand g2079(n3260 ,n3141 ,n3181);
    nand g2080(n1560 ,n1251 ,n662);
    nor g2081(n813 ,n12[8] ,n477);
    nand g2082(n3642 ,n3622 ,n3632);
    nor g2083(n2522 ,n2432 ,n2496);
    not g2084(n442 ,n443);
    nor g2085(n2336 ,n2301 ,n2305);
    nand g2086(n1233 ,n20[10] ,n461);
    nand g2087(n2087 ,n2009 ,n2055);
    xnor g2088(n2106 ,n1945 ,n2037);
    dff g2089(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1452), .Q(n16[8]));
    nand g2090(n933 ,n21[3] ,n454);
    not g2091(n2180 ,n2174);
    nor g2092(n2592 ,n2544 ,n2584);
    not g2093(n2448 ,n2447);
    nor g2094(n2298 ,n2235 ,n2256);
    nand g2095(n3037 ,n2777 ,n2919);
    xnor g2096(n3624 ,n3842 ,n3826);
    xnor g2097(n2365 ,n2324 ,n2284);
    or g2098(n1728 ,n1626 ,n1727);
    nor g2099(n90 ,n27[1] ,n27[0]);
    nor g2100(n2518 ,n2431 ,n2477);
    nand g2101(n1504 ,n1137 ,n743);
    dff g2102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1443), .Q(n16[14]));
    xnor g2103(n2965 ,n2825 ,n2834);
    nand g2104(n2020 ,n3851 ,n1987);
    or g2105(n437 ,n290 ,n425);
    not g2106(n2568 ,n2560);
    nand g2107(n2562 ,n2529 ,n2513);
    nand g2108(n1045 ,n11[5] ,n441);
    xnor g2109(n3046 ,n2797 ,n2948);
    xnor g2110(n3559 ,n3535 ,n2705);
    dff g2111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1519), .Q(n22[12]));
    dff g2112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1518), .Q(n9[13]));
    nand g2113(n3724 ,n3804 ,n3699);
    dff g2114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1459), .Q(n16[4]));
    nand g2115(n1726 ,n1692 ,n1691);
    dff g2116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1427), .Q(n12[1]));
    nand g2117(n3736 ,n3808 ,n3697);
    not g2118(n486 ,n487);
    not g2119(n384 ,n373);
    nand g2120(n47 ,n26[9] ,n44);
    nor g2121(n3020 ,n2751 ,n2954);
    nand g2122(n1605 ,n1066 ,n1028);
    xnor g2123(n3421 ,n3357 ,n3282);
    nor g2124(n2454 ,n2408 ,n2418);
    nand g2125(n874 ,n10[7] ,n502);
    nand g2126(n1638 ,n1177 ,n1180);
    nand g2127(n1937 ,n1916 ,n1911);
    nand g2128(n3487 ,n3414 ,n3466);
    or g2129(n348 ,n199 ,n291);
    nand g2130(n518 ,n204 ,n487);
    nand g2131(n556 ,n189 ,n455);
    nor g2132(n1286 ,n799 ,n773);
    nand g2133(n2817 ,n28[5] ,n26[5]);
    nand g2134(n451 ,n134 ,n407);
    xnor g2135(n1956 ,n1939 ,n1924);
    nand g2136(n961 ,n20[4] ,n452);
    nand g2137(n724 ,n183 ,n480);
    nand g2138(n689 ,n186 ,n442);
    or g2139(n1786 ,n359 ,n1768);
    dff g2140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1393), .Q(n12[14]));
    nor g2141(n785 ,n11[9] ,n479);
    nor g2142(n113 ,n26[0] ,n1);
    nor g2143(n3681 ,n3864 ,n30[7]);
    dff g2144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1493), .Q(n10[3]));
    nand g2145(n2067 ,n1976 ,n2049);
    xnor g2146(n2610 ,n2577 ,n2589);
    nor g2147(n1685 ,n1633 ,n1631);
    nand g2148(n1024 ,n16[6] ,n499);
    nand g2149(n2035 ,n3853 ,n1987);
    nand g2150(n2721 ,n28[6] ,n26[7]);
    xnor g2151(n3327 ,n3228 ,n3119);
    nand g2152(n535 ,n191 ,n453);
    nor g2153(n2239 ,n2182 ,n2220);
    nand g2154(n1014 ,n12[0] ,n486);
    nand g2155(n1948 ,n1924 ,n1939);
    dff g2156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1844), .Q(n5[4]));
    or g2157(n2564 ,n2533 ,n2530);
    dff g2158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1383), .Q(n13[1]));
    nand g2159(n1427 ,n891 ,n518);
    nand g2160(n2908 ,n2736 ,n2808);
    nand g2161(n3769 ,n3688 ,n3701);
    nand g2162(n2775 ,n28[4] ,n26[0]);
    nand g2163(n1661 ,n1256 ,n671);
    xnor g2164(n3285 ,n3172 ,n3093);
    or g2165(n1730 ,n1580 ,n1717);
    nand g2166(n3301 ,n3180 ,n3257);
    nand g2167(n642 ,n180 ,n450);
    xnor g2168(n3560 ,n3543 ,n3532);
    nor g2169(n2480 ,n2406 ,n2440);
    nand g2170(n1396 ,n1003 ,n509);
    nand g2171(n3690 ,n3867 ,n30[4]);
    xnor g2172(n2163 ,n1988 ,n2103);
    nand g2173(n1380 ,n946 ,n573);
    nand g2174(n3667 ,n3617 ,n3666);
    nand g2175(n905 ,n8[10] ,n494);
    xnor g2176(n3152 ,n3004 ,n2731);
    nand g2177(n1020 ,n18[0] ,n456);
    xnor g2178(n2256 ,n2209 ,n2159);
    not g2179(n98 ,n29[6]);
    nand g2180(n3563 ,n3562 ,n3546);
    nor g2181(n387 ,n29[2] ,n353);
    nor g2182(n3709 ,n3698 ,n3681);
    nand g2183(n1079 ,n11[0] ,n441);
    nor g2184(n1820 ,n99 ,n1786);
    nand g2185(n1654 ,n856 ,n1263);
    nand g2186(n1270 ,n15[6] ,n493);
    xnor g2187(n2971 ,n2744 ,n2810);
    nand g2188(n267 ,n24[1] ,n201);
    nand g2189(n325 ,n244 ,n265);
    nand g2190(n3340 ,n3187 ,n3273);
    or g2191(n2413 ,n3814 ,n4[4]);
    xor g2192(n3850 ,n4[0] ,n26[0]);
    nand g2193(n269 ,n1860 ,n206);
    nand g2194(n914 ,n13[11] ,n448);
    nor g2195(n1686 ,n1635 ,n1634);
    nand g2196(n3415 ,n3333 ,n3379);
    dff g2197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1457), .Q(n8[8]));
    not g2198(n2015 ,n2014);
    or g2199(n1788 ,n359 ,n1770);
    xnor g2200(n2573 ,n2511 ,n2534);
    nand g2201(n1801 ,n99 ,n1768);
    nand g2202(n3298 ,n3201 ,n3252);
    nand g2203(n1566 ,n1108 ,n618);
    nand g2204(n1519 ,n1154 ,n643);
    nand g2205(n2720 ,n28[4] ,n26[5]);
    nand g2206(n1527 ,n1166 ,n649);
    nand g2207(n654 ,n187 ,n450);
    nand g2208(n430 ,n334 ,n368);
    nand g2209(n1075 ,n15[0] ,n493);
    nand g2210(n1484 ,n1118 ,n686);
    nor g2211(n2349 ,n2309 ,n2325);
    nand g2212(n2014 ,n27[7] ,n1961);
    nand g2213(n737 ,n187 ,n488);
    or g2214(n3201 ,n3152 ,n3156);
    nand g2215(n2735 ,n28[3] ,n26[7]);
    xnor g2216(n2363 ,n2322 ,n2275);
    not g2217(n107 ,n28[0]);
    nand g2218(n844 ,n306 ,n436);
    nor g2219(n1294 ,n780 ,n768);
    nand g2220(n977 ,n9[6] ,n496);
    nor g2221(n2334 ,n2242 ,n2311);
    nand g2222(n1107 ,n10[9] ,n481);
    dff g2223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n230), .Q(n27[1]));
    nor g2224(n2115 ,n1946 ,n2066);
    nand g2225(n1420 ,n996 ,n609);
    dff g2226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n219), .Q(n27[2]));
    dff g2227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1343), .Q(n23[5]));
    or g2228(n1748 ,n1289 ,n1740);
    nand g2229(n3073 ,n2927 ,n3001);
    nand g2230(n2674 ,n2659 ,n2663);
    xnor g2231(n3849 ,n2345 ,n2401);
    nor g2232(n2565 ,n2487 ,n2522);
    xnor g2233(n3109 ,n2968 ,n2771);
    nand g2234(n1451 ,n1076 ,n623);
    nand g2235(n736 ,n180 ,n490);
    nand g2236(n1428 ,n1014 ,n517);
    or g2237(n29[6] ,n3766 ,n3793);
    nor g2238(n499 ,n208 ,n415);
    nand g2239(n1534 ,n1170 ,n654);
    nand g2240(n1455 ,n1086 ,n715);
    nor g2241(n2272 ,n2115 ,n2247);
    nand g2242(n2854 ,n28[7] ,n26[2]);
    not g2243(n3077 ,n3076);
    nand g2244(n2064 ,n1977 ,n2028);
    not g2245(n210 ,n211);
    xor g2246(n3166 ,n3083 ,n3064);
    nand g2247(n3292 ,n3258 ,n3191);
    nand g2248(n2925 ,n2727 ,n2740);
    nand g2249(n3416 ,n3348 ,n3380);
    xnor g2250(n3110 ,n2963 ,n2778);
    nand g2251(n3546 ,n3537 ,n3520);
    nand g2252(n3551 ,n3532 ,n3543);
    nand g2253(n1227 ,n15[11] ,n493);
    nor g2254(n3701 ,n3698 ,n3674);
    not g2255(n3697 ,n3698);
    nand g2256(n3568 ,n3567 ,n3554);
    or g2257(n3609 ,n3835 ,n3819);
    or g2258(n439 ,n300 ,n424);
    nand g2259(n1552 ,n1243 ,n660);
    nor g2260(n808 ,n12[2] ,n477);
    nand g2261(n2823 ,n27[5] ,n4[6]);
    nand g2262(n971 ,n12[10] ,n486);
    nand g2263(n1406 ,n886 ,n514);
    nand g2264(n1153 ,n22[13] ,n451);
    or g2265(n2649 ,n2469 ,n2639);
    dff g2266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1506), .Q(n14[7]));
    or g2267(n2550 ,n2529 ,n2513);
    nand g2268(n1245 ,n18[12] ,n456);
    nand g2269(n1528 ,n1167 ,n650);
    nand g2270(n592 ,n189 ,n483);
    nand g2271(n2650 ,n2469 ,n2639);
    nand g2272(n1205 ,n14[13] ,n466);
    xnor g2273(n3501 ,n3463 ,n3460);
    nor g2274(n2453 ,n2405 ,n2419);
    xnor g2275(n3154 ,n2974 ,n2906);
    nor g2276(n1303 ,n777 ,n820);
    xnor g2277(n2109 ,n2041 ,n1955);
    nor g2278(n1669 ,n1591 ,n1590);
    nand g2279(n643 ,n181 ,n450);
    nor g2280(n2525 ,n2449 ,n2505);
    dff g2281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1839), .Q(n5[5]));
    nor g2282(n82 ,n26[13] ,n81);
    nor g2283(n816 ,n18[3] ,n475);
    nand g2284(n3748 ,n3840 ,n3685);
    nand g2285(n1575 ,n977 ,n1024);
    nor g2286(n2299 ,n2232 ,n2273);
    nand g2287(n3747 ,n3844 ,n3685);
    dff g2288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1456), .Q(n16[6]));
    nand g2289(n2693 ,n2683 ,n2692);
    dff g2290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1341), .Q(n23[7]));
    nor g2291(n389 ,n126 ,n344);
    not g2292(n2947 ,n2946);
    xnor g2293(n3002 ,n2786 ,n2854);
    nand g2294(n1171 ,n22[2] ,n451);
    xor g2295(n3835 ,n2108 ,n1990);
    nand g2296(n1162 ,n8[2] ,n489);
    not g2297(n3791 ,n3782);
    xnor g2298(n2108 ,n1946 ,n2046);
    xor g2299(n2982 ,n2863 ,n2817);
    not g2300(n2608 ,n2607);
    nor g2301(n3016 ,n2778 ,n2950);
    nand g2302(n570 ,n179 ,n453);
    nand g2303(n3548 ,n3495 ,n3539);
    xnor g2304(n2077 ,n1956 ,n1992);
    nor g2305(n1687 ,n1639 ,n1638);
    nand g2306(n2443 ,n2418 ,n2413);
    nand g2307(n2442 ,n2423 ,n2410);
    xnor g2308(n3806 ,n3663 ,n3627);
    nand g2309(n2941 ,n2815 ,n2715);
    nor g2310(n201 ,n1 ,n172);
    nand g2311(n1443 ,n1054 ,n638);
    nand g2312(n1463 ,n1095 ,n630);
    nand g2313(n513 ,n186 ,n487);
    nand g2314(n137 ,n28[0] ,n28[3]);
    nor g2315(n301 ,n1890 ,n246);
    nand g2316(n1044 ,n14[7] ,n466);
    nand g2317(n3207 ,n3153 ,n3155);
    xnor g2318(n2647 ,n2404 ,n2614);
    nand g2319(n1068 ,n16[14] ,n499);
    nand g2320(n93 ,n27[2] ,n92);
    nand g2321(n3412 ,n3339 ,n3367);
    nand g2322(n2065 ,n1979 ,n2016);
    nand g2323(n1555 ,n1246 ,n636);
    nor g2324(n2352 ,n2338 ,n2329);
    xnor g2325(n3845 ,n2380 ,n2392);
    nand g2326(n623 ,n183 ,n445);
    nand g2327(n960 ,n12[14] ,n486);
    nand g2328(n740 ,n182 ,n490);
    nand g2329(n1091 ,n10[14] ,n481);
    nand g2330(n703 ,n184 ,n458);
    nand g2331(n1095 ,n16[2] ,n444);
    not g2332(n2763 ,n2762);
    nand g2333(n379 ,n280 ,n332);
    nand g2334(n377 ,n260 ,n293);
    nand g2335(n563 ,n186 ,n455);
    nand g2336(n3056 ,n2889 ,n3019);
    not g2337(n2233 ,n2234);
    nand g2338(n1065 ,n16[12] ,n444);
    nor g2339(n1887 ,n68 ,n70);
    dff g2340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1544), .Q(n9[4]));
    xnor g2341(n2075 ,n1955 ,n1966);
    xnor g2342(n215 ,n97 ,n147);
    not g2343(n502 ,n503);
    nor g2344(n3041 ,n2787 ,n2951);
    dff g2345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1474), .Q(n15[11]));
    nand g2346(n1198 ,n15[14] ,n493);
    nand g2347(n624 ,n184 ,n445);
    nand g2348(n970 ,n17[15] ,n484);
    not g2349(n452 ,n453);
    dff g2350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1371), .Q(n21[4]));
    not g2351(n450 ,n451);
    nor g2352(n839 ,n21[8] ,n470);
    nand g2353(n964 ,n17[12] ,n468);
    nand g2354(n1109 ,n15[10] ,n443);
    nand g2355(n1366 ,n927 ,n555);
    nor g2356(n129 ,n29[5] ,n1887);
    not g2357(n1779 ,n1778);
    xnor g2358(n3482 ,n3434 ,n3368);
    not g2359(n212 ,n213);
    not g2360(n2772 ,n2771);
    nand g2361(n2788 ,n27[0] ,n4[0]);
    not g2362(n2505 ,n2504);
    dff g2363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1385), .Q(n20[10]));
    nor g2364(n2896 ,n2735 ,n2829);
    nand g2365(n2085 ,n2001 ,n2034);
    not g2366(n2243 ,n2242);
    nand g2367(n3720 ,n3825 ,n3684);
    nand g2368(n903 ,n9[10] ,n496);
    xnor g2369(n3172 ,n2795 ,n3084);
    nor g2370(n2618 ,n2592 ,n2595);
    nand g2371(n1225 ,n20[11] ,n461);
    dff g2372(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1323), .Q(n17[9]));
    nor g2373(n388 ,n29[3] ,n379);
    nand g2374(n3008 ,n2806 ,n2905);
    nand g2375(n1931 ,n3851 ,n1922);
    nand g2376(n756 ,n188 ,n488);
    nor g2377(n2551 ,n2524 ,n2517);
    nor g2378(n3675 ,n3869 ,n30[2]);
    nand g2379(n3149 ,n2923 ,n3096);
    xnor g2380(n2129 ,n2085 ,n1957);
    nand g2381(n3688 ,n3862 ,n30[9]);
    dff g2382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1369), .Q(n13[6]));
    nand g2383(n1442 ,n1051 ,n620);
    nand g2384(n1546 ,n1188 ,n709);
    nand g2385(n279 ,n25[3] ,n203);
    nand g2386(n2082 ,n1975 ,n2035);
    or g2387(n1733 ,n1603 ,n1720);
    xnor g2388(n2100 ,n1945 ,n2042);
    xnor g2389(n1719 ,n29[0] ,n1470);
    nand g2390(n497 ,n209 ,n405);
    nor g2391(n2475 ,n2408 ,n2437);
    xnor g2392(n3168 ,n3054 ,n3055);
    not g2393(n2068 ,n2069);
    nor g2394(n199 ,n1880 ,n171);
    nand g2395(n3526 ,n3492 ,n3508);
    nand g2396(n2714 ,n27[5] ,n4[3]);
    not g2397(n2953 ,n2936);
    xnor g2398(n30[2] ,n2606 ,n2565);
    nand g2399(n1718 ,n1668 ,n1667);
    nand g2400(n1404 ,n971 ,n614);
    nand g2401(n3177 ,n3057 ,n3104);
    nand g2402(n297 ,n200 ,n221);
    nand g2403(n602 ,n183 ,n455);
    or g2404(n29[7] ,n3773 ,n3794);
    nand g2405(n1551 ,n1240 ,n644);
    nand g2406(n3377 ,n3306 ,n3344);
    not g2407(n2398 ,n2397);
    nand g2408(n2825 ,n27[2] ,n4[6]);
    nand g2409(n1085 ,n16[0] ,n499);
    nand g2410(n2300 ,n2117 ,n2269);
    dff g2411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1547), .Q(n8[0]));
    not g2412(n2445 ,n2446);
    nand g2413(n2730 ,n27[4] ,n4[3]);
    nand g2414(n1653 ,n1261 ,n1262);
    nand g2415(n1940 ,n1906 ,n1919);
    not g2416(n2198 ,n2197);
    xnor g2417(n3276 ,n3169 ,n3103);
    xnor g2418(n185 ,n101 ,n4[10]);
    not g2419(n409 ,n408);
    xnor g2420(n3641 ,n3840 ,n3824);
    nand g2421(n598 ,n182 ,n455);
    nand g2422(n3692 ,n3860 ,n30[11]);
    not g2423(n492 ,n493);
    nand g2424(n3142 ,n3058 ,n3078);
    nand g2425(n3022 ,n2757 ,n2920);
    nand g2426(n852 ,n10[15] ,n502);
    xnor g2427(n3399 ,n3313 ,n3300);
    nand g2428(n527 ,n178 ,n446);
    xnor g2429(n3102 ,n2977 ,n2735);
    nand g2430(n939 ,n21[0] ,n454);
    nand g2431(n2630 ,n2590 ,n2608);
    nand g2432(n111 ,n1882 ,n94);
    nand g2433(n2685 ,n2660 ,n2674);
    nor g2434(n198 ,n1881 ,n171);
    nand g2435(n1494 ,n1126 ,n733);
    nand g2436(n3529 ,n3468 ,n3512);
    not g2437(n2255 ,n2254);
    nor g2438(n3194 ,n3112 ,n3109);
    dff g2439(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1480), .Q(n15[7]));
    nand g2440(n3723 ,n30[11] ,n3699);
    nand g2441(n711 ,n184 ,n440);
    nor g2442(n2764 ,n2706 ,n2709);
    or g2443(n1815 ,n29[9] ,n1793);
    xnor g2444(n2981 ,n2713 ,n2822);
    dff g2445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1543), .Q(n9[5]));
    nand g2446(n2939 ,n2802 ,n2801);
    nand g2447(n628 ,n192 ,n445);
    nor g2448(n828 ,n18[5] ,n475);
    nand g2449(n1651 ,n1042 ,n1044);
    or g2450(n2872 ,n2823 ,n2745);
    nand g2451(n1145 ,n14[5] ,n491);
    dff g2452(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1435), .Q(n11[7]));
    nand g2453(n2727 ,n28[4] ,n26[4]);
    dff g2454(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n238), .Q(n28[4]));
    nand g2455(n1368 ,n930 ,n558);
    nand g2456(n3460 ,n3402 ,n3428);
    xnor g2457(n3542 ,n3516 ,n3502);
    nor g2458(n766 ,n19[3] ,n473);
    nand g2459(n1348 ,n902 ,n532);
    not g2460(n2150 ,n2149);
    nand g2461(n3362 ,n3274 ,n3326);
    nand g2462(n694 ,n179 ,n458);
    nand g2463(n2752 ,n28[4] ,n26[6]);
    dff g2464(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1508), .Q(n14[5]));
    xnor g2465(n2613 ,n2578 ,n2538);
    nand g2466(n1975 ,n3854 ,n1959);
    nor g2467(n121 ,n27[4] ,n27[5]);
    nand g2468(n1178 ,n9[8] ,n459);
    nand g2469(n1127 ,n10[3] ,n481);
    xnor g2470(n3863 ,n3641 ,n3651);
    xnor g2471(n1944 ,n1905 ,n1916);
    nand g2472(n1324 ,n972 ,n508);
    nand g2473(n243 ,n29[4] ,n200);
    dff g2474(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1522), .Q(n9[12]));
    nand g2475(n1330 ,n1004 ,n613);
    nand g2476(n2423 ,n3815 ,n4[5]);
    or g2477(n3252 ,n3159 ,n3222);
    xnor g2478(n2160 ,n1955 ,n2076);
    not g2479(n2757 ,n2756);
    nand g2480(n1497 ,n1130 ,n734);
    nand g2481(n2640 ,n2600 ,n2617);
    nand g2482(n1439 ,n1045 ,n666);
    nand g2483(n1202 ,n14[14] ,n466);
    xnor g2484(n1885 ,n26[7] ,n71);
    not g2485(n208 ,n209);
    nand g2486(n1030 ,n18[14] ,n474);
    nand g2487(n351 ,n278 ,n339);
    xnor g2488(n3163 ,n3058 ,n3078);
    xnor g2489(n188 ,n103 ,n4[14]);
    nand g2490(n1583 ,n862 ,n861);
    nand g2491(n1998 ,n3850 ,n1964);
    nand g2492(n2731 ,n28[2] ,n26[2]);
    nand g2493(n507 ,n185 ,n485);
    nand g2494(n690 ,n204 ,n442);
    nand g2495(n425 ,n305 ,n380);
    nand g2496(n876 ,n17[5] ,n484);
    nand g2497(n2119 ,n1956 ,n2077);
    nand g2498(n1526 ,n1164 ,n648);
    nor g2499(n2222 ,n2074 ,n2192);
    nor g2500(n343 ,n195 ,n304);
    nand g2501(n1336 ,n506 ,n521);
    nand g2502(n667 ,n185 ,n440);
    dff g2503(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1423), .Q(n19[0]));
    xnor g2504(n3420 ,n3355 ,n3332);
    or g2505(n344 ,n198 ,n301);
    nand g2506(n1182 ,n8[15] ,n489);
    nand g2507(n3089 ,n2897 ,n3039);
    nand g2508(n701 ,n185 ,n458);
    nor g2509(n1679 ,n1615 ,n1614);
    nand g2510(n481 ,n141 ,n408);
    nand g2511(n585 ,n190 ,n455);
    nand g2512(n3028 ,n2862 ,n2925);
    nand g2513(n3738 ,n3803 ,n3699);
    xnor g2514(n2277 ,n2230 ,n2164);
    nand g2515(n2852 ,n28[4] ,n26[7]);
    nand g2516(n845 ,n20[1] ,n452);
    dff g2517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1353), .Q(n21[15]));
    xnor g2518(n3478 ,n3192 ,n3447);
    nand g2519(n569 ,n187 ,n449);
    nor g2520(n2292 ,n2238 ,n2261);
    nor g2521(n2172 ,n2097 ,n2151);
    nand g2522(n3375 ,n3302 ,n3320);
    nand g2523(n3510 ,n3419 ,n3491);
    nand g2524(n2729 ,n28[7] ,n26[4]);
    nand g2525(n1082 ,n22[0] ,n463);
    nand g2526(n1438 ,n1047 ,n760);
    nor g2527(n802 ,n15[3] ,n492);
    xnor g2528(n3465 ,n3420 ,n3350);
    nor g2529(n1279 ,n791 ,n841);
    nand g2530(n934 ,n13[5] ,n448);
    nand g2531(n2718 ,n27[1] ,n4[5]);
    xnor g2532(n2125 ,n2062 ,n1957);
    dff g2533(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n236), .Q(n28[0]));
    nand g2534(n3353 ,n3233 ,n3293);
    nor g2535(n3205 ,n3075 ,n3125);
    or g2536(n29[5] ,n3761 ,n3801);
    xnor g2537(n229 ,n161 ,n29[3]);
    dff g2538(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n21[14]));
    xnor g2539(n2993 ,n2855 ,n2765);
    dff g2540(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1568), .Q(n18[2]));
    not g2541(n2569 ,n2561);
    xnor g2542(n2657 ,n2639 ,n2469);
    dff g2543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1538), .Q(n9[10]));
    nand g2544(n1702 ,n1293 ,n1292);
    nand g2545(n3689 ,n3868 ,n30[3]);
    xor g2546(n3815 ,n28[5] ,n27[5]);
    nand g2547(n658 ,n191 ,n457);
    or g2548(n2409 ,n3813 ,n4[3]);
    xnor g2549(n2975 ,n2789 ,n2720);
    nand g2550(n958 ,n11[12] ,n478);
    nand g2551(n262 ,n25[0] ,n203);
    nand g2552(n1836 ,n420 ,n1807);
    nor g2553(n242 ,n27[7] ,n205);
    nand g2554(n1592 ,n877 ,n1070);
    nor g2555(n3703 ,n3698 ,n3676);
    nand g2556(n1622 ,n1214 ,n980);
    xnor g2557(n2687 ,n2668 ,n2661);
    nand g2558(n1010 ,n19[10] ,n482);
    nand g2559(n2737 ,n28[0] ,n26[3]);
    nand g2560(n937 ,n13[4] ,n448);
    nand g2561(n3406 ,n3385 ,n3373);
    nand g2562(n930 ,n21[5] ,n454);
    dff g2563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1454), .Q(n16[7]));
    not g2564(n440 ,n441);
    dff g2565(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1433), .Q(n11[9]));
    nand g2566(n475 ,n207 ,n414);
    nor g2567(n3682 ,n3859 ,n30[12]);
    xnor g2568(n219 ,n149 ,n29[2]);
    xnor g2569(n224 ,n159 ,n29[6]);
    nand g2570(n2118 ,n1957 ,n2078);
    nand g2571(n2623 ,n2564 ,n2605);
    nand g2572(n254 ,n29[14] ,n202);
    nand g2573(n1412 ,n984 ,n536);
    nand g2574(n1321 ,n853 ,n612);
    dff g2575(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1486), .Q(n15[4]));
    xor g2576(n178 ,n4[5] ,n29[5]);
    nand g2577(n581 ,n184 ,n453);
    nand g2578(n1802 ,n96 ,n1774);
    nand g2579(n2009 ,n3858 ,n1959);
    nand g2580(n1418 ,n993 ,n566);
    not g2581(n2238 ,n2237);
    xnor g2582(n3228 ,n3130 ,n3081);
    nand g2583(n2809 ,n28[2] ,n26[7]);
    nor g2584(n1313 ,n839 ,n772);
    nand g2585(n2185 ,n2133 ,n2128);
    nand g2586(n3076 ,n2899 ,n3045);
    or g2587(n1749 ,n1297 ,n1741);
    nand g2588(n1449 ,n1067 ,n691);
    not g2589(n364 ,n363);
    nand g2590(n702 ,n183 ,n458);
    nand g2591(n89 ,n28[2] ,n88);
    nand g2592(n3666 ,n3636 ,n3665);
    nor g2593(n3372 ,n3298 ,n3328);
    xor g2594(n3438 ,n3408 ,n3386);
    dff g2595(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1499), .Q(n14[12]));
    nand g2596(n1445 ,n1058 ,n672);
    nor g2597(n3300 ,n3211 ,n3245);
    nand g2598(n969 ,n12[11] ,n486);
    nor g2599(n814 ,n18[8] ,n475);
    dff g2600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1390), .Q(n12[15]));
    nand g2601(n1548 ,n1040 ,n692);
    nor g2602(n1689 ,n1643 ,n1642);
    dff g2603(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1334), .Q(n23[14]));
    nor g2604(n1986 ,n1951 ,n1958);
    not g2605(n3284 ,n3283);
    nor g2606(n120 ,n26[9] ,n26[10]);
    or g2607(n1758 ,n1314 ,n1743);
    nand g2608(n568 ,n191 ,n455);
    or g2609(n50 ,n26[11] ,n48);
    dff g2610(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n226), .Q(n28[3]));
    nor g2611(n797 ,n21[5] ,n470);
    nand g2612(n926 ,n21[7] ,n454);
    or g2613(n2886 ,n2826 ,n2730);
    not g2614(n371 ,n356);
    dff g2615(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1516), .Q(n22[13]));
    nand g2616(n546 ,n185 ,n449);
    nor g2617(n461 ,n213 ,n415);
    nand g2618(n3497 ,n3424 ,n3482);
    xnor g2619(n3445 ,n3390 ,n3401);
    dff g2620(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1434), .Q(n11[8]));
    nor g2621(n1690 ,n1647 ,n1646);
    nand g2622(n3538 ,n3501 ,n3528);
    dff g2623(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1505), .Q(n14[8]));
    nand g2624(n3025 ,n2753 ,n2913);
    dff g2625(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1539), .Q(n9[9]));
    nand g2626(n1565 ,n1103 ,n723);
    xor g2627(n2704 ,n3098 ,n3089);
    nand g2628(n1326 ,n881 ,n512);
    nor g2629(n3680 ,n3865 ,n30[6]);
    nand g2630(n163 ,n1894 ,n94);
    nand g2631(n114 ,n1883 ,n94);
    nand g2632(n1966 ,n3850 ,n1958);
    nor g2633(n2469 ,n2406 ,n2424);
    nand g2634(n268 ,n24[0] ,n201);
    nand g2635(n1617 ,n1258 ,n1207);
    xnor g2636(n1957 ,n1940 ,n1914);
    nand g2637(n3742 ,n30[12] ,n3699);
    xnor g2638(n2279 ,n2228 ,n2249);
    nand g2639(n1933 ,n3857 ,n1922);
    xnor g2640(n2973 ,n2820 ,n2722);
    nor g2641(n779 ,n17[3] ,n469);
    xnor g2642(n1893 ,n28[2] ,n87);
    or g2643(n1757 ,n1306 ,n1742);
    nand g2644(n2117 ,n2071 ,n2069);
    nand g2645(n1103 ,n10[10] ,n481);
    xnor g2646(n1890 ,n26[2] ,n62);
    nand g2647(n949 ,n20[11] ,n452);
    nand g2648(n394 ,n5[9] ,n359);
    xnor g2649(n2145 ,n2088 ,n1956);
    or g2650(n2414 ,n3816 ,n4[6]);
    nand g2651(n695 ,n188 ,n458);
    nand g2652(n2749 ,n27[5] ,n4[4]);
    nand g2653(n1168 ,n22[5] ,n451);
    not g2654(n2593 ,n2592);
    nand g2655(n3774 ,n3689 ,n3703);
    nor g2656(n2335 ,n2289 ,n2315);
    xnor g2657(n3264 ,n3154 ,n3186);
    nor g2658(n2509 ,n2460 ,n2489);
    nand g2659(n421 ,n5[13] ,n359);
    not g2660(n3302 ,n3301);
    nand g2661(n336 ,n26[8] ,n247);
    not g2662(n101 ,n29[10]);
    or g2663(n1731 ,n1588 ,n1718);
    nand g2664(n523 ,n185 ,n446);
    xnor g2665(n2097 ,n2040 ,n1946);
    xnor g2666(n2310 ,n2207 ,n2263);
    or g2667(n3576 ,n26[1] ,n4[1]);
    nand g2668(n257 ,n1881 ,n206);
    dff g2669(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1546), .Q(n9[2]));
    nand g2670(n1828 ,n398 ,n1809);
    xnor g2671(n3162 ,n3066 ,n3076);
    nand g2672(n3075 ,n2890 ,n3024);
    nor g2673(n3651 ,n3611 ,n3650);
    not g2674(n2302 ,n2293);
    nand g2675(n1036 ,n12[4] ,n476);
    nand g2676(n857 ,n9[7] ,n496);
    nor g2677(n3011 ,n2734 ,n2900);
    nand g2678(n675 ,n179 ,n440);
    xnor g2679(n2984 ,n2809 ,n2813);
    nand g2680(n577 ,n182 ,n453);
    or g2681(n36 ,n26[4] ,n34);
    not g2682(n2329 ,n2328);
    nand g2683(n1117 ,n10[6] ,n481);
    nand g2684(n1419 ,n994 ,n574);
    xor g2685(n3813 ,n28[3] ,n27[3]);
    not g2686(n1945 ,n1946);
    xnor g2687(n2230 ,n2162 ,n2111);
    dff g2688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1856), .Q(n5[9]));
    nand g2689(n629 ,n187 ,n445);
    nand g2690(n600 ,n183 ,n487);
    nor g2691(n2526 ,n2450 ,n2504);
    nand g2692(n2050 ,n3853 ,n2015);
    nor g2693(n2946 ,n2758 ,n2755);
    nor g2694(n3611 ,n3839 ,n3823);
    nand g2695(n1338 ,n1275 ,n523);
    xnor g2696(n2614 ,n2573 ,n2518);
    not g2697(n110 ,n7);
    nor g2698(n2291 ,n2237 ,n2262);
    nor g2699(n2151 ,n2110 ,n2120);
    nand g2700(n3786 ,n3693 ,n3708);
    xnor g2701(n2962 ,n2793 ,n2828);
    nand g2702(n710 ,n182 ,n440);
    or g2703(n3137 ,n2903 ,n3059);
    nand g2704(n2836 ,n28[3] ,n26[5]);
    nand g2705(n3458 ,n3381 ,n3418);
    nand g2706(n552 ,n184 ,n449);
    nand g2707(n1831 ,n403 ,n1811);
    or g2708(n1769 ,n1701 ,n1748);
    nand g2709(n612 ,n182 ,n485);
    nand g2710(n1774 ,n1693 ,n1759);
    nand g2711(n728 ,n189 ,n480);
    nand g2712(n743 ,n183 ,n490);
    nand g2713(n1096 ,n16[1] ,n444);
    or g2714(n1735 ,n1618 ,n1722);
    nor g2715(n2948 ,n2786 ,n2854);
    xnor g2716(n3323 ,n3226 ,n3127);
    nand g2717(n3208 ,n3107 ,n3100);
    nand g2718(n992 ,n10[4] ,n502);
    nand g2719(n924 ,n21[8] ,n454);
    xnor g2720(n3634 ,n3836 ,n3820);
    nand g2721(n211 ,n27[2] ,n176);
    nand g2722(n1621 ,n1212 ,n1007);
    nand g2723(n3601 ,n3585 ,n3600);
    dff g2724(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1340), .Q(n23[8]));
    nand g2725(n1919 ,n27[6] ,n1904);
    nand g2726(n2248 ,n2187 ,n2224);
    or g2727(n3267 ,n3258 ,n3191);
    nand g2728(n296 ,n200 ,n232);
    nand g2729(n1008 ,n11[14] ,n478);
    xnor g2730(n2322 ,n2287 ,n2254);
    nand g2731(n1190 ,n15[15] ,n493);
    nand g2732(n645 ,n185 ,n450);
    nand g2733(n2069 ,n1984 ,n2048);
    not g2734(n3279 ,n3278);
    or g2735(n2549 ,n2523 ,n2521);
    xnor g2736(n3515 ,n3441 ,n3490);
    nor g2737(n1823 ,n101 ,n1792);
    nand g2738(n875 ,n11[6] ,n478);
    nand g2739(n2079 ,n1972 ,n2025);
    nand g2740(n880 ,n10[0] ,n502);
    nor g2741(n1305 ,n818 ,n832);
    nand g2742(n1457 ,n1089 ,n714);
    nand g2743(n3029 ,n2839 ,n2931);
    nand g2744(n427 ,n267 ,n345);
    xnor g2745(n2140 ,n2069 ,n2067);
    nor g2746(n2581 ,n2566 ,n2402);
    nand g2747(n2664 ,n2631 ,n2651);
    dff g2748(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1414), .Q(n19[6]));
    nand g2749(n994 ,n12[5] ,n486);
    nor g2750(n833 ,n23[9] ,n464);
    nand g2751(n1229 ,n16[11] ,n499);
    nand g2752(n1700 ,n1287 ,n1286);
    nor g2753(n2376 ,n2340 ,n2364);
    dff g2754(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1439), .Q(n11[5]));
    nand g2755(n1697 ,n1279 ,n1278);
    not g2756(n3486 ,n3485);
    nor g2757(n2355 ,n2341 ,n2331);
    nand g2758(n1477 ,n1111 ,n761);
    dff g2759(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1509), .Q(n9[15]));
    nand g2760(n1221 ,n16[12] ,n499);
    nand g2761(n2921 ,n2735 ,n2829);
    nand g2762(n2815 ,n28[2] ,n26[5]);
    not g2763(n2860 ,n2859);
    nand g2764(n909 ,n13[14] ,n448);
    nand g2765(n745 ,n189 ,n490);
    not g2766(n3057 ,n3056);
    nor g2767(n2241 ,n2229 ,n2201);
    nand g2768(n194 ,n1884 ,n144);
    dff g2769(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1447), .Q(n16[12]));
    nand g2770(n1538 ,n1172 ,n701);
    nand g2771(n1047 ,n8[10] ,n489);
    xnor g2772(n3860 ,n3626 ,n3657);
    nor g2773(n823 ,n23[2] ,n464);
    xnor g2774(n3625 ,n3841 ,n3825);
    dff g2775(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1335), .Q(n23[13]));
    xnor g2776(n3640 ,n3839 ,n3823);
    nand g2777(n1655 ,n1026 ,n1264);
    not g2778(n2571 ,n2563);
    xnor g2779(n2632 ,n2579 ,n2599);
    nor g2780(n318 ,n283 ,n246);
    nand g2781(n2758 ,n28[4] ,n26[1]);
    nand g2782(n317 ,n26[1] ,n247);
    nand g2783(n665 ,n204 ,n457);
    nor g2784(n3700 ,n3698 ,n3673);
    xor g2785(n3869 ,n3834 ,n3818);
    not g2786(n2503 ,n2502);
    nand g2787(n656 ,n204 ,n450);
    xor g2788(n2978 ,n2766 ,n2743);
    dff g2789(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n325), .Q(n24[5]));
    not g2790(n143 ,n142);
    nand g2791(n3734 ,n3821 ,n3684);
    or g2792(n193 ,n1891 ,n144);
    nand g2793(n1510 ,n1146 ,n748);
    nand g2794(n1537 ,n1174 ,n657);
    xnor g2795(n2977 ,n2787 ,n2829);
    nand g2796(n1155 ,n14[1] ,n491);
    not g2797(n3636 ,n3635);
    dff g2798(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1321), .Q(n17[11]));
    nor g2799(n61 ,n26[1] ,n26[0]);
    nor g2800(n1293 ,n806 ,n787);
    nand g2801(n594 ,n190 ,n485);
    nand g2802(n3378 ,n3303 ,n3317);
    nand g2803(n3032 ,n2863 ,n2928);
    nor g2804(n2433 ,n2405 ,n2417);
    nand g2805(n540 ,n180 ,n449);
    nand g2806(n1421 ,n998 ,n553);
    nand g2807(n1006 ,n11[10] ,n478);
    nand g2808(n2563 ,n2534 ,n2511);
    nand g2809(n622 ,n185 ,n445);
    xnor g2810(n3848 ,n2362 ,n2399);
    nor g2811(n1760 ,n1645 ,n1737);
    dff g2812(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1419), .Q(n12[5]));
    nand g2813(n2856 ,n27[6] ,n4[7]);
    nand g2814(n1255 ,n18[5] ,n456);
    xnor g2815(n3273 ,n3170 ,n3059);
    nand g2816(n73 ,n26[7] ,n72);
    nand g2817(n1084 ,n16[7] ,n444);
    nand g2818(n1166 ,n22[7] ,n451);
    nand g2819(n281 ,n1864 ,n206);
    nand g2820(n51 ,n26[11] ,n48);
    nand g2821(n1607 ,n1195 ,n979);
    nor g2822(n2307 ,n2252 ,n2286);
    nand g2823(n1554 ,n1245 ,n637);
    xnor g2824(n3446 ,n3392 ,n3301);
    nand g2825(n2935 ,n2723 ,n2816);
    not g2826(n2073 ,n2072);
    nand g2827(n506 ,n23[12] ,n447);
    nand g2828(n626 ,n189 ,n445);
    nor g2829(n773 ,n8[3] ,n495);
    nand g2830(n1370 ,n934 ,n562);
    dff g2831(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1342), .Q(n23[6]));
    nand g2832(n869 ,n17[0] ,n484);
    nand g2833(n1611 ,n1200 ,n1030);
    nand g2834(n3567 ,n3552 ,n3566);
    nand g2835(n641 ,n185 ,n457);
    nand g2836(n699 ,n182 ,n458);
    nand g2837(n1226 ,n12[11] ,n476);
    xnor g2838(n3821 ,n3391 ,n3385);
    nand g2839(n3572 ,n3571 ,n3533);
    dff g2840(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1557), .Q(n8[14]));
    nand g2841(n2250 ,n2189 ,n2226);
    nand g2842(n923 ,n21[9] ,n454);
    or g2843(n1903 ,n28[4] ,n28[3]);
    nand g2844(n1590 ,n1062 ,n887);
    nand g2845(n3789 ,n3696 ,n3709);
    or g2846(n3471 ,n3417 ,n3446);
    nor g2847(n2945 ,n2849 ,n2837);
    nand g2848(n428 ,n5[12] ,n359);
    nand g2849(n2813 ,n28[5] ,n26[4]);
    nand g2850(n1598 ,n882 ,n1085);
    nor g2851(n2901 ,n2767 ,n2843);
    nand g2852(n951 ,n20[10] ,n452);
    nand g2853(n280 ,n1880 ,n206);
    dff g2854(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1551), .Q(n18[14]));
    nand g2855(n1835 ,n401 ,n1801);
    nor g2856(n2884 ,n2728 ,n2791);
    nand g2857(n333 ,n26[14] ,n247);
    nand g2858(n246 ,n174 ,n201);
    nand g2859(n1407 ,n1010 ,n601);
    xnor g2860(n3272 ,n3165 ,n3122);
    nand g2861(n3783 ,n3691 ,n3706);
    xnor g2862(n3516 ,n3491 ,n3419);
    xnor g2863(n3584 ,n4[4] ,n26[4]);
    nand g2864(n1263 ,n16[7] ,n499);
    nand g2865(n3148 ,n2795 ,n3085);
    dff g2866(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1570), .Q(n18[1]));
    nand g2867(n1211 ,n12[13] ,n476);
    nand g2868(n760 ,n185 ,n488);
    xnor g2869(n183 ,n102 ,n4[9]);
    nand g2870(n1532 ,n1181 ,n754);
    or g2871(n40 ,n26[6] ,n38);
    nor g2872(n2337 ,n2302 ,n2316);
    nand g2873(n1707 ,n1308 ,n1307);
    nand g2874(n2651 ,n2623 ,n2637);
    nand g2875(n2724 ,n27[5] ,n4[0]);
    nand g2876(n1337 ,n1276 ,n522);
    nor g2877(n1670 ,n1593 ,n1592);
    nand g2878(n1999 ,n3852 ,n1964);
    xnor g2879(n2204 ,n2123 ,n2154);
    nand g2880(n3157 ,n2867 ,n3073);
    nand g2881(n3067 ,n2893 ,n3031);
    nand g2882(n2086 ,n2008 ,n2057);
    not g2883(n2553 ,n2547);
    nand g2884(n49 ,n26[10] ,n46);
    nand g2885(n591 ,n178 ,n483);
    nand g2886(n2369 ,n2351 ,n2327);
    nand g2887(n1403 ,n885 ,n597);
    nand g2888(n1329 ,n866 ,n617);
    xnor g2889(n3133 ,n2993 ,n2945);
    nor g2890(n1683 ,n1625 ,n1624);
    nor g2891(n302 ,n201 ,n218);
    dff g2892(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1397), .Q(n20[1]));
    nand g2893(n1778 ,n1687 ,n1755);
    nand g2894(n3379 ,n3263 ,n3345);
    nor g2895(n3338 ,n3279 ,n3277);
    dff g2896(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1492), .Q(n15[0]));
    nand g2897(n345 ,n194 ,n298);
    nor g2898(n2426 ,n2407 ,n2417);
    nand g2899(n3049 ,n2946 ,n2996);
    nand g2900(n2701 ,n2649 ,n2700);
    nand g2901(n3339 ,n3259 ,n3297);
    nor g2902(n3336 ,n3260 ,n3282);
    not g2903(n478 ,n479);
    nand g2904(n3730 ,n30[2] ,n3699);
    nand g2905(n2697 ,n2682 ,n2696);
    xor g2906(n2404 ,n2402 ,n2566);
    nand g2907(n2797 ,n27[6] ,n4[4]);
    nand g2908(n1811 ,n29[5] ,n1762);
    not g2909(n362 ,n361);
    dff g2910(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1661), .Q(n11[14]));
    nand g2911(n538 ,n188 ,n449);
    not g2912(n2777 ,n2776);
    nor g2913(n3657 ,n3616 ,n3656);
    xnor g2914(n1924 ,n28[3] ,n27[3]);
    nand g2915(n3733 ,n30[3] ,n3699);
    nor g2916(n2458 ,n2405 ,n2418);
    nand g2917(n1851 ,n394 ,n1815);
    not g2918(n496 ,n497);
    nand g2919(n3765 ,n3686 ,n3700);
    nand g2920(n3209 ,n3152 ,n3156);
    nor g2921(n1695 ,n1659 ,n1658);
    nand g2922(n670 ,n192 ,n440);
    nand g2923(n1447 ,n1065 ,n633);
    nor g2924(n2457 ,n2408 ,n2419);
    xnor g2925(n3331 ,n3232 ,n3243);
    dff g2926(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1374), .Q(n21[1]));
    nor g2927(n768 ,n9[2] ,n497);
    nand g2928(n1161 ,n14[0] ,n491);
    nand g2929(n2827 ,n27[1] ,n4[0]);
    nor g2930(n2112 ,n2066 ,n2069);
    not g2931(n1773 ,n1772);
    nor g2932(n2378 ,n2350 ,n2366);
    nand g2933(n907 ,n13[15] ,n448);
    nand g2934(n620 ,n179 ,n445);
    nand g2935(n605 ,n183 ,n485);
    dff g2936(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1336), .Q(n23[12]));
    nand g2937(n2226 ,n2107 ,n2185);
    xnor g2938(n3118 ,n2979 ,n2741);
    xnor g2939(n3627 ,n3846 ,n3830);
    nand g2940(n533 ,n180 ,n446);
    nor g2941(n1665 ,n1579 ,n1578);
    nand g2942(n3212 ,n3093 ,n3148);
    xnor g2943(n2078 ,n1957 ,n1965);
    or g2944(n2282 ,n2214 ,n2259);
    nor g2945(n784 ,n8[2] ,n495);
    not g2946(n2366 ,n2365);
    xnor g2947(n2107 ,n1956 ,n2047);
    nand g2948(n1242 ,n12[14] ,n476);
    nand g2949(n1467 ,n1099 ,n676);
    or g2950(n3533 ,n3501 ,n3528);
    dff g2951(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1358), .Q(n21[12]));
    nor g2952(n1672 ,n1599 ,n1598);
    nand g2953(n2928 ,n2817 ,n2833);
    xnor g2954(n2970 ,n2801 ,n2802);
    nor g2955(n1680 ,n1617 ,n1616);
    nand g2956(n997 ,n12[8] ,n486);
    or g2957(n2873 ,n2809 ,n2813);
    xnor g2958(n3637 ,n3837 ,n3821);
    nand g2959(n256 ,n29[6] ,n200);
    nand g2960(n2738 ,n28[6] ,n26[5]);
    nand g2961(n1039 ,n11[7] ,n441);
    nand g2962(n432 ,n5[11] ,n359);
    nand g2963(n610 ,n183 ,n483);
    nor g2964(n1900 ,n28[7] ,n27[7]);
    nor g2965(n3699 ,n3670 ,n3);
    nand g2966(n2802 ,n28[2] ,n26[4]);
    not g2967(n92 ,n91);
    xnor g2968(n3155 ,n2982 ,n2833);
    nor g2969(n3211 ,n3082 ,n3119);
    dff g2970(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1405), .Q(n19[12]));
    nand g2971(n1219 ,n12[6] ,n476);
    nor g2972(n2598 ,n2546 ,n2585);
    nand g2973(n1037 ,n16[4] ,n499);
    nand g2974(n1658 ,n1270 ,n846);
    nand g2975(n3366 ,n3283 ,n3324);
    nand g2976(n1070 ,n12[0] ,n476);
    nand g2977(n2692 ,n2671 ,n2691);
    not g2978(n1913 ,n1912);
    nor g2979(n3613 ,n3838 ,n3822);
    nor g2980(n3215 ,n3079 ,n3123);
    nand g2981(n3364 ,n3275 ,n3325);
    nand g2982(n1099 ,n15[15] ,n443);
    nand g2983(n1509 ,n1142 ,n694);
    not g2984(n2286 ,n2285);
    nand g2985(n916 ,n13[10] ,n448);
    nand g2986(n2001 ,n3857 ,n1959);
    nand g2987(n1067 ,n11[1] ,n441);
    nand g2988(n3744 ,n3809 ,n3697);
    nand g2989(n1016 ,n8[7] ,n494);
    nor g2990(n2394 ,n2379 ,n2393);
    nor g2991(n3083 ,n2884 ,n3016);
    xnor g2992(n3171 ,n2991 ,n3086);
    or g2993(n29[3] ,n3785 ,n3799);
    nand g2994(n908 ,n19[10] ,n472);
    xnor g2995(n3004 ,n2762 ,n2799);
    nand g2996(n3045 ,n2766 ,n2932);
    nor g2997(n3305 ,n3214 ,n3246);
    nor g2998(n832 ,n14[9] ,n467);
    nand g2999(n112 ,n24[7] ,n94);
    nand g3000(n1071 ,n8[9] ,n489);
    nand g3001(n1175 ,n9[9] ,n459);
    xnor g3002(n3358 ,n3305 ,n3279);
    nand g3003(n29[14] ,n3745 ,n3791);
    nand g3004(n91 ,n27[1] ,n27[0]);
    nand g3005(n3741 ,n3827 ,n3684);
    nand g3006(n3793 ,n3714 ,n3765);
    nand g3007(n3176 ,n3061 ,n3137);
    nand g3008(n1612 ,n1201 ,n1248);
    not g3009(n460 ,n461);
    nand g3010(n2799 ,n28[0] ,n26[4]);
    xnor g3011(n3354 ,n3101 ,n3285);
    xnor g3012(n30[7] ,n2686 ,n2692);
    nand g3013(n64 ,n26[2] ,n63);
    nand g3014(n609 ,n186 ,n483);
    nor g3015(n2472 ,n2406 ,n2421);
    or g3016(n295 ,n203 ,n239);
    nand g3017(n615 ,n184 ,n487);
    nand g3018(n2835 ,n28[2] ,n26[6]);
    or g3019(n29[1] ,n3790 ,n3796);
    not g3020(n59 ,n26[8]);
    nand g3021(n2913 ,n2746 ,n2717);
    nand g3022(n2675 ,n2632 ,n2664);
    xnor g3023(n3503 ,n3464 ,n3432);
    nand g3024(n2812 ,n28[1] ,n26[3]);
    nor g3025(n2275 ,n2190 ,n2241);
    nor g3026(n3706 ,n3698 ,n3677);
    nand g3027(n1436 ,n1041 ,n758);
    nand g3028(n2314 ,n2300 ,n2265);
    dff g3029(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1406), .Q(n19[11]));
    dff g3030(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1840), .Q(n5[3]));
    nand g3031(n2421 ,n3810 ,n4[0]);
    nand g3032(n999 ,n19[1] ,n482);
    nand g3033(n966 ,n8[4] ,n494);
    dff g3034(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1475), .Q(n15[10]));
    nand g3035(n2759 ,n27[5] ,n4[1]);
    xnor g3036(n2096 ,n1957 ,n2043);
    nand g3037(n938 ,n21[1] ,n454);
    nor g3038(n463 ,n211 ,n415);
    xnor g3039(n2132 ,n2079 ,n1955);
    nand g3040(n1333 ,n888 ,n519);
    nand g3041(n1260 ,n20[7] ,n461);
    nand g3042(n1235 ,n21[10] ,n471);
    nor g3043(n2456 ,n2408 ,n2417);
    nor g3044(n1750 ,n1589 ,n1731);
    nand g3045(n1387 ,n953 ,n578);
    nand g3046(n541 ,n181 ,n449);
    nand g3047(n1055 ,n13[1] ,n501);
    nand g3048(n422 ,n333 ,n385);
    dff g3049(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1375), .Q(n13[4]));
    nand g3050(n1984 ,n3853 ,n1960);
    dff g3051(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n439), .Q(n26[7]));
    nand g3052(n2283 ,n2214 ,n2259);
    nand g3053(n3547 ,n3527 ,n3534);
    xnor g3054(n3808 ,n3667 ,n3629);
    nand g3055(n1967 ,n3856 ,n1960);
    nand g3056(n2791 ,n27[4] ,n4[5]);
    nand g3057(n693 ,n191 ,n442);
    nand g3058(n1118 ,n15[5] ,n443);
    xnor g3059(n2572 ,n2514 ,n2512);
    nor g3060(n836 ,n15[8] ,n492);
    nand g3061(n1129 ,n8[5] ,n489);
    nand g3062(n1879 ,n37 ,n36);
    nand g3063(n2044 ,n1928 ,n1999);
    xor g3064(n3868 ,n3631 ,n3622);
    or g3065(n3343 ,n3248 ,n3304);
    nand g3066(n3756 ,n3837 ,n3685);
    nand g3067(n402 ,n303 ,n347);
    nor g3068(n2766 ,n2708 ,n2707);
    nand g3069(n981 ,n19[8] ,n482);
    nand g3070(n744 ,n184 ,n490);
    not g3071(n368 ,n352);
    not g3072(n476 ,n477);
    dff g3073(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1401), .Q(n19[15]));
    nor g3074(n455 ,n137 ,n416);
    nor g3075(n3012 ,n2806 ,n2905);
    nand g3076(n3668 ,n3630 ,n3667);
    nand g3077(n1642 ,n908 ,n1236);
    nand g3078(n2814 ,n28[2] ,n26[3]);
    nand g3079(n3150 ,n3089 ,n3072);
    nor g3080(n827 ,n14[2] ,n467);
    nand g3081(n1425 ,n906 ,n539);
    nand g3082(n618 ,n187 ,n457);
    nand g3083(n259 ,n25[4] ,n203);
    not g3084(n2153 ,n2152);
    not g3085(n2199 ,n2181);
    nand g3086(n1657 ,n1268 ,n875);
    nor g3087(n805 ,n23[3] ,n464);
    nand g3088(n1191 ,n12[15] ,n476);
    nand g3089(n2929 ,n2814 ,n2807);
    not g3090(n472 ,n473);
    xnor g3091(n2278 ,n2234 ,n2236);
    nand g3092(n2861 ,n27[6] ,n4[2]);
    nand g3093(n2024 ,n3856 ,n1986);
    nor g3094(n1905 ,n28[3] ,n27[3]);
    nand g3095(n761 ,n184 ,n480);
    nor g3096(n501 ,n213 ,n406);
    nor g3097(n3246 ,n3092 ,n3215);
    nand g3098(n1618 ,n1208 ,n1209);
    nor g3099(n2463 ,n2407 ,n2423);
    dff g3100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1337), .Q(n23[11]));
    nand g3101(n3352 ,n3256 ,n3289);
    not g3102(n79 ,n78);
    nand g3103(n580 ,n183 ,n453);
    or g3104(n3495 ,n3457 ,n3484);
    xnor g3105(n2074 ,n1991 ,n1946);
    xnor g3106(n2264 ,n2206 ,n2138);
    nand g3107(n2508 ,n2468 ,n2501);
    xnor g3108(n177 ,n98 ,n1886);
    not g3109(n3585 ,n3584);
    xnor g3110(n1914 ,n27[7] ,n28[7]);
    dff g3111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1432), .Q(n11[10]));
    nor g3112(n2528 ,n2434 ,n2491);
    nor g3113(n3307 ,n3194 ,n3250);
    nand g3114(n3735 ,n3806 ,n3697);
    xor g3115(n218 ,n146 ,n29[5]);
    nor g3116(n3656 ,n3624 ,n3655);
    nand g3117(n1081 ,n20[0] ,n461);
    nand g3118(n2920 ,n2809 ,n2813);
    dff g3119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1566), .Q(n18[3]));
    nand g3120(n1332 ,n869 ,n511);
    or g3121(n1904 ,n28[6] ,n28[5]);
    not g3122(n462 ,n463);
    or g3123(n2619 ,n2556 ,n2599);
    nand g3124(n3385 ,n3295 ,n3347);
    dff g3125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1344), .Q(n23[4]));
    nor g3126(n203 ,n1 ,n174);
    nand g3127(n145 ,n24[0] ,n94);
    nand g3128(n3346 ,n3105 ,n3271);
    xnor g3129(n3357 ,n3260 ,n3286);
    not g3130(n3281 ,n3280);
    nand g3131(n1604 ,n1192 ,n1191);
    nand g3132(n1596 ,n1078 ,n1077);
    nand g3133(n3039 ,n2702 ,n2912);
    nand g3134(n3051 ,n2945 ,n2994);
    nand g3135(n2080 ,n1970 ,n2018);
    nand g3136(n668 ,n190 ,n440);
    nor g3137(n2294 ,n2274 ,n2264);
    xnor g3138(n1889 ,n26[3] ,n64);
    xnor g3139(n2134 ,n2080 ,n1957);
    nand g3140(n3017 ,n2761 ,n2941);
    or g3141(n2487 ,n2407 ,n2444);
    nand g3142(n1641 ,n1235 ,n1234);
    nand g3143(n3536 ,n3511 ,n3526);
    xnor g3144(n2678 ,n2656 ,n2654);
    nor g3145(n2584 ,n2518 ,n2571);
    dff g3146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1536), .Q(n22[1]));
    nand g3147(n1215 ,n23[12] ,n465);
    nand g3148(n677 ,n188 ,n442);
    nand g3149(n1563 ,n1255 ,n664);
    nand g3150(n2620 ,n2558 ,n2604);
    nand g3151(n726 ,n190 ,n490);
    nand g3152(n967 ,n20[0] ,n452);
    dff g3153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1436), .Q(n8[11]));
    nand g3154(n1625 ,n1197 ,n1196);
    dff g3155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1466), .Q(n16[0]));
    nand g3156(n158 ,n25[2] ,n94);
    nand g3157(n3253 ,n3161 ,n3203);
    nand g3158(n3725 ,n3819 ,n3684);
    xnor g3159(n3423 ,n3354 ,n3306);
    nor g3160(n2483 ,n2405 ,n2444);
    xnor g3161(n3590 ,n4[5] ,n26[5]);
    not g3162(n2998 ,n2997);
    nand g3163(n748 ,n192 ,n490);
    nand g3164(n1108 ,n18[3] ,n456);
    nand g3165(n530 ,n186 ,n446);
    xnor g3166(n3156 ,n2972 ,n2859);
    xnor g3167(n1872 ,n26[12] ,n80);
    nand g3168(n528 ,n192 ,n446);
    xnor g3169(n3265 ,n3219 ,n3105);
    nand g3170(n757 ,n179 ,n488);
    nand g3171(n3409 ,n3319 ,n3371);
    not g3172(n2161 ,n2160);
    nand g3173(n3428 ,n3352 ,n3396);
    nand g3174(n2936 ,n2864 ,n2788);
    nor g3175(n788 ,n9[8] ,n497);
    xnor g3176(n3847 ,n2372 ,n2396);
    nand g3177(n1706 ,n1304 ,n1303);
    nand g3178(n1487 ,n1120 ,n688);
    xnor g3179(n2655 ,n2625 ,n2615);
    nand g3180(n649 ,n190 ,n450);
    nor g3181(n819 ,n22[9] ,n462);
    xnor g3182(n3243 ,n3134 ,n3068);
    nand g3183(n1763 ,n1666 ,n1747);
    not g3184(n2798 ,n2797);
    xnor g3185(n2122 ,n2083 ,n1955);
    not g3186(n2532 ,n2531);
    dff g3187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1558), .Q(n18[9]));
    xnor g3188(n3391 ,n3217 ,n3330);
    nand g3189(n2072 ,n1982 ,n2054);
    xnor g3190(n3519 ,n3484 ,n3457);
    xnor g3191(n2615 ,n2575 ,n2520);
    nand g3192(n1355 ,n915 ,n545);
    nor g3193(n3662 ,n3633 ,n3661);
    not g3194(n2216 ,n2215);
    nand g3195(n1434 ,n1034 ,n711);
    xor g3196(n2165 ,n2070 ,n2109);
    not g3197(n206 ,n205);
    nand g3198(n43 ,n26[7] ,n40);
    or g3199(n2603 ,n2570 ,n2588);
    nand g3200(n663 ,n189 ,n457);
    dff g3201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1563), .Q(n18[5]));
    dff g3202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1417), .Q(n19[4]));
    nand g3203(n1865 ,n56 ,n55);
    nand g3204(n1699 ,n1285 ,n1284);
    nand g3205(n520 ,n188 ,n446);
    nand g3206(n706 ,n178 ,n458);
    nand g3207(n213 ,n27[2] ,n142);
    nand g3208(n424 ,n338 ,n358);
    nand g3209(n3454 ,n3350 ,n3420);
    nand g3210(n1397 ,n845 ,n596);
    nand g3211(n2934 ,n2744 ,n2810);
    nor g3212(n1755 ,n1637 ,n1744);
    nand g3213(n1069 ,n16[11] ,n444);
    xor g3214(n184 ,n4[8] ,n29[8]);
    dff g3215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1328), .Q(n17[4]));
    nand g3216(n3047 ,n2902 ,n2997);
    nand g3217(n1531 ,n1163 ,n699);
    dff g3218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n13[10]));
    not g3219(n2288 ,n2287);
    not g3220(n2200 ,n2183);
    dff g3221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1366), .Q(n13[7]));
    xnor g3222(n2324 ,n2260 ,n2289);
    xnor g3223(n3827 ,n3559 ,n3563);
    nand g3224(n1256 ,n11[14] ,n441);
    nand g3225(n3596 ,n3576 ,n3595);
    dff g3226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1346), .Q(n23[2]));
    nand g3227(n863 ,n17[7] ,n484);
    xor g3228(n2402 ,n2485 ,n2472);
    xnor g3229(n3356 ,n3297 ,n3259);
    nor g3230(n2557 ,n2447 ,n2532);
    xnor g3231(n3805 ,n3661 ,n3633);
    xnor g3232(n1943 ,n1899 ,n1917);
    nand g3233(n1394 ,n961 ,n588);
    nand g3234(n3475 ,n3407 ,n3440);
    nand g3235(n3694 ,n3859 ,n30[12]);
    nand g3236(n1150 ,n9[13] ,n459);
    nand g3237(n1541 ,n1179 ,n704);
    xnor g3238(n3165 ,n3080 ,n3092);
    nand g3239(n1564 ,n1259 ,n653);
    dff g3240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n427), .Q(n24[1]));
    nor g3241(n3676 ,n3868 ,n30[3]);
    nand g3242(n646 ,n179 ,n457);
    nand g3243(n995 ,n19[11] ,n472);
    nor g3244(n2658 ,n2628 ,n2646);
    xnor g3245(n227 ,n165 ,n29[9]);
    not g3246(n3398 ,n3397);
    xnor g3247(n2972 ,n2739 ,n2812);
    nand g3248(n575 ,n181 ,n453);
    nand g3249(n1059 ,n21[1] ,n471);
    nand g3250(n1354 ,n914 ,n542);
    not g3251(n60 ,n26[12]);
    nand g3252(n3622 ,n3834 ,n3818);
    nand g3253(n1143 ,n14[6] ,n491);
    nand g3254(n1137 ,n14[9] ,n491);
    or g3255(n3467 ,n3399 ,n3442);
    nand g3256(n3031 ,n2848 ,n2929);
    dff g3257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1430), .Q(n11[11]));
    or g3258(n3349 ,n3105 ,n3271);
    nand g3259(n972 ,n17[8] ,n484);
    nand g3260(n1701 ,n1291 ,n1290);
    dff g3261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1372), .Q(n15[14]));
    nor g3262(n2313 ,n2296 ,n2299);
    dff g3263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1360), .Q(n13[9]));
    nor g3264(n241 ,n26[15] ,n196);
    not g3265(n3632 ,n3631);
    nand g3266(n2354 ,n2318 ,n2332);
    nor g3267(n3803 ,n2407 ,n2435);
    nor g3268(n2358 ,n2321 ,n2335);
    nor g3269(n3658 ,n3626 ,n3657);
    dff g3270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1450), .Q(n16[10]));
    xnor g3271(n217 ,n96 ,n160);
    or g3272(n1844 ,n1819 ,n1832);
    dff g3273(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1421), .Q(n12[4]));
    nor g3274(n831 ,n21[9] ,n470);
    nand g3275(n1705 ,n1302 ,n1301);
    nand g3276(n576 ,n204 ,n449);
    nand g3277(n273 ,n1863 ,n206);
    nand g3278(n2021 ,n3854 ,n1987);
    nand g3279(n1724 ,n1686 ,n1685);
    nand g3280(n532 ,n191 ,n446);
    nand g3281(n1064 ,n22[1] ,n463);
    nor g3282(n3578 ,n26[6] ,n4[6]);
    xnor g3283(n3829 ,n3558 ,n3567);
    xnor g3284(n2677 ,n2653 ,n2655);
    nand g3285(n1768 ,n1672 ,n1751);
    nand g3286(n1559 ,n1250 ,n635);
    nand g3287(n584 ,n189 ,n453);
    dff g3288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1571), .Q(n8[13]));
    nand g3289(n1021 ,n18[6] ,n474);
    nand g3290(n1623 ,n1215 ,n1223);
    nand g3291(n2830 ,n28[0] ,n26[2]);
    nand g3292(n2789 ,n27[6] ,n4[3]);
    xnor g3293(n2285 ,n2121 ,n2250);
    nand g3294(n1170 ,n22[3] ,n451);
    nand g3295(n991 ,n9[11] ,n496);
    nand g3296(n865 ,n17[4] ,n484);
    nand g3297(n1053 ,n20[1] ,n461);
    nand g3298(n1011 ,n11[13] ,n478);
    nor g3299(n1676 ,n1607 ,n1606);
    nand g3300(n980 ,n8[12] ,n494);
    xnor g3301(n3853 ,n3593 ,n3598);
    xnor g3302(n2686 ,n2667 ,n2658);
    or g3303(n1783 ,n359 ,n1769);
    nand g3304(n2006 ,n3853 ,n1963);
    nor g3305(n2527 ,n2457 ,n2483);
    xnor g3306(n2609 ,n2576 ,n2403);
    nand g3307(n3761 ,n3712 ,n3711);
    nor g3308(n1307 ,n817 ,n786);
    nand g3309(n1520 ,n1155 ,n752);
    or g3310(n29[4] ,n3787 ,n3800);
    xnor g3311(n1918 ,n27[2] ,n27[1]);
    nand g3312(n2560 ,n2512 ,n2514);
    not g3313(n3324 ,n3323);
    xnor g3314(n2624 ,n2597 ,n2598);
    nand g3315(n3069 ,n2878 ,n3040);
    xnor g3316(n3101 ,n2989 ,n2856);
    nand g3317(n2186 ,n2125 ,n2130);
    nand g3318(n989 ,n12[6] ,n486);
    nor g3319(n2513 ,n2454 ,n2492);
    nand g3320(n491 ,n141 ,n407);
    nand g3321(n2696 ,n2681 ,n2695);
    nor g3322(n2473 ,n2406 ,n2442);
    nand g3323(n1516 ,n1153 ,n642);
    xnor g3324(n3105 ,n2981 ,n2850);
    nand g3325(n1017 ,n19[7] ,n472);
    dff g3326(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1332), .Q(n17[0]));
    nand g3327(n1698 ,n1283 ,n1282);
    nand g3328(n554 ,n184 ,n455);
    nand g3329(n2386 ,n2354 ,n2385);
    nand g3330(n156 ,n24[5] ,n94);
    nor g3331(n2543 ,n2448 ,n2531);
    nor g3332(n1821 ,n96 ,n1780);
    xnor g3333(n3541 ,n3488 ,n3521);
    nor g3334(n2343 ,n2297 ,n2313);
    nor g3335(n2488 ,n2405 ,n2439);
    dff g3336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1491), .Q(n10[4]));
    xnor g3337(n3229 ,n3112 ,n3109);
    xnor g3338(n2251 ,n2215 ,n2099);
    xnor g3339(n180 ,n104 ,n4[13]);
    or g3340(n3290 ,n3205 ,n3243);
    xnor g3341(n3824 ,n3519 ,n3529);
    nor g3342(n2491 ,n2405 ,n2435);
    nand g3343(n3288 ,n3179 ,n3237);
    nand g3344(n1384 ,n949 ,n577);
    dff g3345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1399), .Q(n19[13]));
    nand g3346(n943 ,n8[11] ,n494);
    nand g3347(n337 ,n26[10] ,n247);
    nor g3348(n2588 ,n2526 ,n2555);
    nand g3349(n2919 ,n2821 ,n2718);
    nor g3350(n287 ,n129 ,n246);
    xor g3351(n2705 ,n3517 ,n3503);
    nor g3352(n2297 ,n2198 ,n2258);
    nand g3353(n2743 ,n27[7] ,n4[4]);
    nand g3354(n1608 ,n1202 ,n1242);
    xnor g3355(n223 ,n166 ,n29[13]);
    nor g3356(n3250 ,n3131 ,n3221);
    nand g3357(n2034 ,n3856 ,n1987);
    dff g3358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1540), .Q(n9[8]));
    nand g3359(n3511 ,n3458 ,n3486);
    dff g3360(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n227), .Q(n28[1]));
    nor g3361(n2373 ,n2334 ,n2371);
    nand g3362(n495 ,n209 ,n404);
    nor g3363(n3648 ,n3638 ,n3647);
    nand g3364(n2819 ,n28[3] ,n26[2]);
    nor g3365(n2347 ,n2320 ,n2326);
    nand g3366(n1535 ,n1171 ,n655);
    dff g3367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1330), .Q(n17[2]));
    nand g3368(n548 ,n181 ,n455);
    xnor g3369(n3320 ,n3230 ,n3117);
    xnor g3370(n237 ,n157 ,n29[4]);
    nand g3371(n1709 ,n1312 ,n1311);
    nand g3372(n680 ,n182 ,n442);
    nand g3373(n433 ,n309 ,n369);
    nand g3374(n327 ,n253 ,n261);
    nand g3375(n1057 ,n18[1] ,n474);
    nand g3376(n1976 ,n3852 ,n1960);
    nand g3377(n3455 ,n3411 ,n3423);
    nand g3378(n2808 ,n27[2] ,n4[1]);
    nand g3379(n900 ,n23[2] ,n447);
    nand g3380(n288 ,n177 ,n245);
    or g3381(n1297 ,n809 ,n808);
    nand g3382(n3714 ,n30[6] ,n3699);
    nor g3383(n2451 ,n2408 ,n2424);
    nand g3384(n1949 ,n1923 ,n1941);
    not g3385(n174 ,n173);
    xnor g3386(n232 ,n111 ,n29[3]);
    nand g3387(n3788 ,n3741 ,n3739);
    nand g3388(n1249 ,n18[9] ,n456);
    nand g3389(n854 ,n19[12] ,n482);
    dff g3390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1532), .Q(n8[1]));
    nand g3391(n459 ,n139 ,n410);
    nand g3392(n1197 ,n21[12] ,n471);
    dff g3393(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1527), .Q(n22[7]));
    or g3394(n2600 ,n2528 ,n2580);
    nand g3395(n3257 ,n3157 ,n3202);
    nand g3396(n698 ,n181 ,n458);
    nand g3397(n277 ,n25[1] ,n203);
    nand g3398(n3426 ,n3267 ,n3413);
    nand g3399(n983 ,n11[15] ,n478);
    nand g3400(n1004 ,n17[2] ,n484);
    nor g3401(n2391 ,n2390 ,n2377);
    xnor g3402(n3153 ,n2958 ,n2752);
    or g3403(n3199 ,n3153 ,n3155);
    nand g3404(n3745 ,n3848 ,n3685);
    nand g3405(n1220 ,n18[12] ,n474);
    or g3406(n436 ,n387 ,n389);
    nand g3407(n3749 ,n3841 ,n3685);
    nand g3408(n3395 ,n3322 ,n3368);
    nand g3409(n2639 ,n2548 ,n2619);
    nand g3410(n1180 ,n18[11] ,n474);
    nand g3411(n1742 ,n1305 ,n1715);
    not g3412(n2996 ,n2995);
    nor g3413(n144 ,n95 ,n1);
    xnor g3414(n3540 ,n3528 ,n3501);
    xnor g3415(n2136 ,n1957 ,n2087);
    dff g3416(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1402), .Q(n12[11]));
    nor g3417(n2466 ,n2406 ,n2420);
    nand g3418(n1739 ,n1280 ,n1712);
    nor g3419(n115 ,n28[0] ,n1);
    nor g3420(n483 ,n137 ,n409);
    nand g3421(n1586 ,n872 ,n873);
    nand g3422(n2631 ,n2552 ,n2613);
    nor g3423(n1826 ,n104 ,n1789);
    or g3424(n3499 ,n3444 ,n3483);
    or g3425(n1738 ,n1652 ,n1726);
    nand g3426(n3802 ,n3753 ,n3768);
    nand g3427(n1570 ,n1269 ,n665);
    nand g3428(n1186 ,n9[3] ,n459);
    nand g3429(n3801 ,n3731 ,n3789);
    nand g3430(n3068 ,n2907 ,n3043);
    nor g3431(n123 ,n26[5] ,n26[6]);
    not g3432(n2750 ,n2749);
    dff g3433(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1317), .Q(n17[15]));
    nand g3434(n2726 ,n27[6] ,n4[0]);
    nand g3435(n1853 ,n428 ,n1827);
    nor g3436(n3650 ,n3640 ,n3649);
    nand g3437(n2698 ,n2680 ,n2697);
    nand g3438(n1518 ,n1150 ,n696);
    nor g3439(n3710 ,n3698 ,n3682);
    nor g3440(n810 ,n16[2] ,n498);
    nand g3441(n3753 ,n3842 ,n3685);
    nor g3442(n2485 ,n2407 ,n2443);
    nand g3443(n950 ,n13[1] ,n448);
    or g3444(n1847 ,n1823 ,n1830);
    nand g3445(n335 ,n26[12] ,n247);
    nand g3446(n196 ,n120 ,n131);
    nor g3447(n118 ,n29[7] ,n1885);
    nand g3448(n2265 ,n2233 ,n2236);
    nand g3449(n727 ,n190 ,n480);
    nand g3450(n1038 ,n14[4] ,n466);
    nand g3451(n583 ,n190 ,n453);
    nand g3452(n3799 ,n3756 ,n3783);
    nand g3453(n1363 ,n922 ,n552);
    nand g3454(n1498 ,n1132 ,n731);
    nand g3455(n349 ,n262 ,n295);
    nand g3456(n3173 ,n3060 ,n3126);
    nand g3457(n539 ,n187 ,n487);
    nand g3458(n1072 ,n18[0] ,n474);
    nand g3459(n1878 ,n39 ,n38);
    nand g3460(n1643 ,n1237 ,n1165);
    not g3461(n2405 ,n5[2]);
    dff g3462(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1534), .Q(n22[3]));
    not g3463(n3120 ,n3119);
    xnor g3464(n2967 ,n2808 ,n2736);
    nand g3465(n166 ,n25[5] ,n94);
    or g3466(n438 ,n302 ,n426);
    nand g3467(n1251 ,n18[7] ,n456);
    xnor g3468(n2589 ,n2470 ,n2537);
    nor g3469(n2308 ,n2287 ,n2255);
    nand g3470(n1410 ,n997 ,n615);
    nand g3471(n998 ,n12[4] ,n486);
    nand g3472(n3528 ,n3475 ,n3509);
    nor g3473(n1756 ,n1619 ,n1735);
    nand g3474(n2672 ,n2654 ,n2656);
    or g3475(n2889 ,n2812 ,n2739);
    xnor g3476(n2098 ,n1945 ,n2044);
    nand g3477(n2717 ,n28[7] ,n26[3]);
    xnor g3478(n225 ,n148 ,n29[15]);
    nand g3479(n988 ,n19[5] ,n482);
    xnor g3480(n3103 ,n2985 ,n2815);
    nand g3481(n3751 ,n3834 ,n3685);
    xor g3482(n3817 ,n28[7] ,n27[7]);
    not g3483(n202 ,n203);
    nand g3484(n253 ,n29[13] ,n202);
    nand g3485(n1252 ,n11[15] ,n441);
    dff g3486(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1356), .Q(n21[13]));
    nand g3487(n2601 ,n2528 ,n2580);
    xnor g3488(n2669 ,n2642 ,n2623);
    nand g3489(n927 ,n13[7] ,n448);
    nand g3490(n1157 ,n22[10] ,n451);
    nand g3491(n3345 ,n3190 ,n3300);
    or g3492(n29[2] ,n3780 ,n3797);
    nand g3493(n1580 ,n1035 ,n1199);
    dff g3494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1477), .Q(n10[8]));
    nand g3495(n3470 ,n3386 ,n3452);
    nand g3496(n1351 ,n910 ,n540);
    nand g3497(n151 ,n25[6] ,n94);
    xnor g3498(n2956 ,n2719 ,n2819);
    nor g3499(n2356 ,n2342 ,n2330);
    nand g3500(n847 ,n17[14] ,n468);
    xnor g3501(n2259 ,n2203 ,n2229);
    nand g3502(n3721 ,n3829 ,n3684);
    nand g3503(n604 ,n190 ,n487);
    nand g3504(n910 ,n13[13] ,n448);
    nand g3505(n587 ,n178 ,n453);
    nand g3506(n441 ,n139 ,n408);
    nand g3507(n1383 ,n950 ,n576);
    nand g3508(n1083 ,n16[8] ,n444);
    not g3509(n385 ,n374);
    nand g3510(n529 ,n187 ,n446);
    nor g3511(n2231 ,n2099 ,n2216);
    dff g3512(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n327), .Q(n25[5]));
    nand g3513(n2829 ,n27[5] ,n4[5]);
    xnor g3514(n2611 ,n2574 ,n2588);
    nand g3515(n3244 ,n3090 ,n3173);
    nor g3516(n1712 ,n1697 ,n1696);
    or g3517(n1902 ,n28[2] ,n28[1]);
    nand g3518(n1491 ,n1124 ,n730);
    dff g3519(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1400), .Q(n20[0]));
    nand g3520(n1992 ,n3850 ,n1963);
    nand g3521(n894 ,n23[8] ,n447);
    nand g3522(n1930 ,n3852 ,n1922);
    nand g3523(n2007 ,n3852 ,n1963);
    nand g3524(n1243 ,n18[13] ,n456);
    nand g3525(n1431 ,n1022 ,n716);
    dff g3526(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n399), .Q(n26[10]));
    nand g3527(n1523 ,n1157 ,n645);
    nor g3528(n798 ,n16[3] ,n498);
    nor g3529(n1674 ,n1630 ,n1602);
    nor g3530(n75 ,n26[9] ,n74);
    or g3531(n1846 ,n1817 ,n1834);
    nand g3532(n3296 ,n3193 ,n3244);
    nand g3533(n1000 ,n17[10] ,n468);
    nand g3534(n261 ,n25[5] ,n203);
    or g3535(n2195 ,n2070 ,n2129);
    or g3536(n2867 ,n2811 ,n2716);
    or g3537(n2545 ,n2512 ,n2514);
    nand g3538(n1244 ,n8[14] ,n489);
    nand g3539(n1717 ,n1665 ,n1664);
    nand g3540(n3787 ,n3740 ,n3759);
    nand g3541(n378 ,n279 ,n292);
    nand g3542(n3023 ,n2750 ,n2918);
    nor g3543(n3053 ,n2945 ,n2994);
    nand g3544(n2940 ,n2828 ,n2793);
    nand g3545(n1098 ,n16[0] ,n444);
    nand g3546(n525 ,n190 ,n446);
    nor g3547(n2430 ,n2408 ,n2420);
    dff g3548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1389), .Q(n20[7]));
    nor g3549(n1894 ,n88 ,n86);
    nand g3550(n650 ,n189 ,n450);
    xor g3551(n2986 ,n2764 ,n2730);
    nand g3552(n3778 ,n3690 ,n3705);
    nand g3553(n1094 ,n10[13] ,n481);
    nand g3554(n1034 ,n11[8] ,n441);
    nand g3555(n608 ,n192 ,n483);
    nor g3556(n2240 ,n2175 ,n2219);
    nand g3557(n2831 ,n28[3] ,n26[3]);
    nand g3558(n1969 ,n3854 ,n1960);
    nand g3559(n2422 ,n3813 ,n4[3]);
    or g3560(n2384 ,n2347 ,n2383);
    xor g3561(n3164 ,n3060 ,n3090);
    nand g3562(n315 ,n26[5] ,n247);
    nand g3563(n2811 ,n27[3] ,n4[1]);
    nor g3564(n2904 ,n2782 ,n2775);
    nor g3565(n360 ,n27[6] ,n319);
    or g3566(n1781 ,n359 ,n1762);
    nand g3567(n993 ,n19[3] ,n482);
    nand g3568(n1997 ,n3853 ,n1964);
    or g3569(n3136 ,n3054 ,n3055);
    nand g3570(n3492 ,n3456 ,n3477);
    nand g3571(n1051 ,n16[15] ,n444);
    xnor g3572(n1883 ,n27[2] ,n91);
    xnor g3573(n3442 ,n3393 ,n3353);
    nor g3574(n2489 ,n2408 ,n2440);
    nor g3575(n790 ,n9[3] ,n497);
    not g3576(n2471 ,n2470);
    nor g3577(n2425 ,n2405 ,n2421);
    nand g3578(n1035 ,n18[4] ,n474);
    nand g3579(n1907 ,n28[2] ,n28[1]);
    nor g3580(n3607 ,n3587 ,n3606);
    nand g3581(n1980 ,n3856 ,n1958);
    nand g3582(n1105 ,n15[12] ,n443);
    nand g3583(n168 ,n29[4] ,n1888);
    not g3584(n3220 ,n3204);
    xnor g3585(n2162 ,n2059 ,n2096);
    nand g3586(n944 ,n20[14] ,n452);
    dff g3587(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n329), .Q(n25[7]));
    nand g3588(n512 ,n189 ,n485);
    nor g3589(n3702 ,n3698 ,n3675);
    xnor g3590(n3836 ,n2210 ,n2156);
    nand g3591(n859 ,n19[4] ,n472);
    nand g3592(n595 ,n182 ,n487);
    nor g3593(n3408 ,n3342 ,n3374);
    nand g3594(n536 ,n190 ,n483);
    nand g3595(n2723 ,n27[1] ,n4[6]);
    nand g3596(n3780 ,n3730 ,n3755);
    nand g3597(n3602 ,n3580 ,n3601);
    nand g3598(n1640 ,n1000 ,n1233);
    nor g3599(n2493 ,n2406 ,n2443);
    nand g3600(n2849 ,n28[1] ,n26[1]);
    nor g3601(n1716 ,n1709 ,n1708);
    not g3602(n369 ,n354);
    nand g3603(n272 ,n1861 ,n206);
    nand g3604(n712 ,n183 ,n440);
    nand g3605(n1365 ,n926 ,n585);
    nand g3606(n555 ,n190 ,n449);
    nand g3607(n1741 ,n1296 ,n1714);
    nand g3608(n551 ,n185 ,n455);
    dff g3609(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1545), .Q(n9[3]));
    nor g3610(n1776 ,n1707 ,n1757);
    dff g3611(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1846), .Q(n5[1]));
    nor g3612(n2375 ,n2359 ,n2370);
    nor g3613(n3679 ,n3867 ,n30[4]);
    xnor g3614(n3332 ,n3231 ,n3159);
    nor g3615(n1300 ,n770 ,n812);
    nand g3616(n263 ,n24[7] ,n201);
    nand g3617(n1446 ,n1060 ,n634);
    nand g3618(n661 ,n183 ,n457);
    nand g3619(n1115 ,n10[7] ,n481);
    nor g3620(n2470 ,n2406 ,n2418);
    nand g3621(n1062 ,n23[1] ,n465);
    xnor g3622(n3191 ,n2962 ,n3095);
    nand g3623(n553 ,n192 ,n487);
    nor g3624(n2379 ,n2349 ,n2365);
    nand g3625(n29[15] ,n3758 ,n3776);
    nor g3626(n3334 ,n3259 ,n3297);
    nand g3627(n3502 ,n3467 ,n3487);
    nand g3628(n562 ,n178 ,n449);
    dff g3629(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1542), .Q(n9[6]));
    nor g3630(n1667 ,n1585 ,n1584);
    nand g3631(n1784 ,n360 ,n1766);
    not g3632(n3275 ,n3274);
    not g3633(n2258 ,n2257);
    xnor g3634(n2102 ,n1945 ,n2038);
    nand g3635(n1489 ,n1122 ,n689);
    nor g3636(n3616 ,n3842 ,n3826);
    nand g3637(n1429 ,n1020 ,n658);
    xnor g3638(n2327 ,n2278 ,n2300);
    nand g3639(n2783 ,n27[2] ,n4[4]);
    nand g3640(n2838 ,n27[5] ,n4[7]);
    nor g3641(n3033 ,n2768 ,n2952);
    dff g3642(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1381), .Q(n13[2]));
    xnor g3643(n228 ,n112 ,n29[7]);
    xnor g3644(n3485 ,n3436 ,n3442);
    nand g3645(n1026 ,n23[7] ,n465);
    nand g3646(n1983 ,n3853 ,n1959);
    nor g3647(n1873 ,n82 ,n84);
    not g3648(n2955 ,n2942);
    xnor g3649(n2594 ,n2541 ,n2519);
    nor g3650(n3417 ,n3409 ,n3400);
    nand g3651(n853 ,n17[11] ,n484);
    or g3652(n29[9] ,n3788 ,n3798);
    nand g3653(n3739 ,n30[9] ,n3699);
    nand g3654(n3619 ,n3846 ,n3830);
    nor g3655(n3605 ,n3586 ,n3604);
    nand g3656(n429 ,n5[15] ,n359);
    nand g3657(n2801 ,n27[4] ,n4[2]);
    or g3658(n3545 ,n3537 ,n3520);
    not g3659(n2338 ,n2337);
    xor g3660(n1866 ,n26[14] ,n54);
    nand g3661(n573 ,n180 ,n453);
    nor g3662(n769 ,n19[2] ,n473);
    nand g3663(n1503 ,n1140 ,n742);
    nand g3664(n963 ,n19[6] ,n482);
    nor g3665(n2496 ,n2408 ,n2435);
    or g3666(n2871 ,n2737 ,n2732);
    dff g3667(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1440), .Q(n11[4]));
    or g3668(n2682 ,n2662 ,n2669);
    nor g3669(n1283 ,n781 ,n828);
    nand g3670(n2092 ,n2004 ,n2022);
    nand g3671(n692 ,n204 ,n458);
    nand g3672(n1881 ,n33 ,n32);
    or g3673(n3472 ,n3407 ,n3440);
    xnor g3674(n2332 ,n2281 ,n2256);
    nand g3675(n906 ,n12[3] ,n486);
    nand g3676(n1398 ,n860 ,n560);
    xnor g3677(n3834 ,n1945 ,n1962);
    nand g3678(n2249 ,n2195 ,n2223);
    not g3679(n2148 ,n2147);
    nand g3680(n614 ,n185 ,n487);
    nand g3681(n891 ,n12[1] ,n486);
    nand g3682(n447 ,n136 ,n407);
    not g3683(n2597 ,n2596);
    dff g3684(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1467), .Q(n15[15]));
    nand g3685(n707 ,n192 ,n458);
    nand g3686(n2444 ,n2419 ,n2415);
    nand g3687(n1860 ,n45 ,n44);
    nand g3688(n361 ,n109 ,n321);
    nand g3689(n2385 ,n2348 ,n2384);
    not g3690(n2099 ,n2098);
    nand g3691(n2083 ,n1980 ,n2036);
    nor g3692(n777 ,n9[9] ,n497);
    nand g3693(n153 ,n25[0] ,n94);
    nand g3694(n3365 ,n3284 ,n3323);
    nand g3695(n1496 ,n1131 ,n736);
    nor g3696(n824 ,n20[2] ,n460);
    xnor g3697(n3425 ,n3359 ,n3303);
    nand g3698(n1112 ,n15[9] ,n443);
    xnor g3699(n3113 ,n2978 ,n2794);
    dff g3700(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1338), .Q(n23[10]));
    nor g3701(n1301 ,n830 ,n778);
    or g3702(n3396 ,n3296 ,n3369);
    nand g3703(n294 ,n202 ,n234);
    nand g3704(n1971 ,n3853 ,n1958);
    not g3705(n466 ,n467);
    nand g3706(n2911 ,n2812 ,n2739);
    nand g3707(n2056 ,n3857 ,n1985);
    nand g3708(n3505 ,n3443 ,n3489);
    nand g3709(n849 ,n19[15] ,n482);
    nor g3710(n2539 ,n2462 ,n2499);
    nand g3711(n3488 ,n3430 ,n3471);
    not g3712(n2262 ,n2261);
    or g3713(n3507 ,n3419 ,n3491);
    nand g3714(n671 ,n188 ,n440);
    dff g3715(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1471), .Q(n10[9]));
    nand g3716(n890 ,n23[13] ,n447);
    dff g3717(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1719), .Q(n6));
    nand g3718(n1261 ,n21[7] ,n471);
    nand g3719(n2224 ,n2159 ,n2186);
    nor g3720(n3685 ,n2 ,n3);
    nand g3721(n1996 ,n3851 ,n1964);
    not g3722(n2725 ,n2724);
    nand g3723(n2716 ,n27[4] ,n4[0]);
    dff g3724(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1487), .Q(n15[3]));
    nand g3725(n1662 ,n504 ,n1470);
    xnor g3726(n3558 ,n3542 ,n3536);
    nand g3727(n2052 ,n3855 ,n2015);
    nand g3728(n974 ,n12[9] ,n486);
    nor g3729(n1766 ,n1704 ,n1749);
    not g3730(n2774 ,n2773);
    nand g3731(n1216 ,n20[12] ,n461);
    nand g3732(n1276 ,n23[11] ,n447);
    not g3733(n2253 ,n2252);
    nor g3734(n197 ,n28[6] ,n173);
    nand g3735(n1236 ,n16[10] ,n499);
    nand g3736(n1476 ,n1112 ,n682);
    nand g3737(n664 ,n178 ,n457);
    dff g3738(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1376), .Q(n21[0]));
    xnor g3739(n3866 ,n3637 ,n3645);
    nand g3740(n2713 ,n28[6] ,n26[6]);
    nor g3741(n2530 ,n2456 ,n2490);
    nand g3742(n1200 ,n13[14] ,n501);
    nand g3743(n1479 ,n1110 ,n721);
    nand g3744(n2622 ,n2545 ,n2602);
    nand g3745(n1377 ,n942 ,n570);
    nand g3746(n621 ,n182 ,n445);
    nor g3747(n1818 ,n98 ,n1795);
    not g3748(n2342 ,n2341);
    nand g3749(n383 ,n28[1] ,n321);
    nand g3750(n148 ,n25[7] ,n94);
    nand g3751(n652 ,n192 ,n450);
    dff g3752(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1420), .Q(n19[2]));
    nand g3753(n2859 ,n27[1] ,n4[3]);
    xnor g3754(n191 ,n99 ,n4[0]);
    nand g3755(n1012 ,n17[15] ,n468);
    nor g3756(n3532 ,n3514 ,n3524);
    nor g3757(n3092 ,n2879 ,n3033);
    xnor g3758(n3282 ,n3163 ,n3065);
    nand g3759(n601 ,n185 ,n483);
    nand g3760(n3206 ,n3112 ,n3109);
    or g3761(n3175 ,n3127 ,n3115);
    nand g3762(n574 ,n178 ,n487);
    xnor g3763(n3387 ,n3296 ,n3352);
    or g3764(n2634 ,n2586 ,n2610);
    not g3765(n366 ,n365);
    nor g3766(n408 ,n28[2] ,n383);
    nor g3767(n2546 ,n2510 ,n2515);
    not g3768(n2436 ,n2437);
    nand g3769(n2059 ,n1993 ,n2053);
    nand g3770(n1485 ,n1117 ,n728);
    nand g3771(n2036 ,n3855 ,n1986);
    nor g3772(n2459 ,n2408 ,n2422);
    nor g3773(n2490 ,n2405 ,n2437);
    xnor g3774(n3820 ,n3309 ,n3261);
    xnor g3775(n3167 ,n3063 ,n3056);
    or g3776(n2411 ,n3817 ,n4[7]);
    nand g3777(n1342 ,n896 ,n526);
    nand g3778(n1536 ,n1173 ,n656);
    nand g3779(n3418 ,n3363 ,n3412);
    xor g3780(n3816 ,n28[6] ,n27[6]);
    nand g3781(n2689 ,n2666 ,n2685);
    nand g3782(n1974 ,n3855 ,n1959);
    nand g3783(n2744 ,n28[1] ,n26[5]);
    nand g3784(n2932 ,n2794 ,n2743);
    xnor g3785(n3588 ,n4[1] ,n26[1]);
    nand g3786(n381 ,n169 ,n287);
    nand g3787(n3081 ,n2883 ,n3034);
    nand g3788(n1459 ,n1092 ,n628);
    nand g3789(n2781 ,n27[0] ,n4[2]);
    nand g3790(n2937 ,n2831 ,n2726);
    nand g3791(n2710 ,n27[5] ,n4[2]);
    nand g3792(n3297 ,n3196 ,n3234);
    nor g3793(n791 ,n19[5] ,n473);
    or g3794(n32 ,n26[2] ,n31);
    dff g3795(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1367), .Q(n21[6]));
    not g3796(n2179 ,n2173);
    nand g3797(n1092 ,n16[4] ,n444);
    not g3798(n2950 ,n2917);
    not g3799(n370 ,n355);
    nand g3800(n135 ,n28[3] ,n107);
    nor g3801(n1796 ,n29[12] ,n1773);
    nor g3802(n842 ,n26[4] ,n505);
    xnor g3803(n1946 ,n1912 ,n1909);
    nor g3804(n3659 ,n3615 ,n3658);
    dff g3805(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1449), .Q(n11[1]));
    nand g3806(n157 ,n24[4] ,n94);
    nand g3807(n1619 ,n1011 ,n1210);
    dff g3808(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n400), .Q(n26[8]));
    nor g3809(n2903 ,n2855 ,n2765);
    not g3810(n3591 ,n3590);
    not g3811(n88 ,n87);
    nor g3812(n2182 ,n2155 ,n2122);
    nand g3813(n3580 ,n26[4] ,n4[4]);
    nand g3814(n1852 ,n429 ,n1824);
    dff g3815(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1387), .Q(n13[0]));
    not g3816(n505 ,n504);
    nor g3817(n2051 ,n1898 ,n2014);
    nand g3818(n2042 ,n1927 ,n1997);
    nand g3819(n162 ,n1893 ,n94);
    or g3820(n2887 ,n2817 ,n2833);
    not g3821(n2320 ,n2319);
    dff g3822(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1496), .Q(n14[13]));
    nand g3823(n1921 ,n27[4] ,n1903);
    nand g3824(n260 ,n25[2] ,n203);
    dff g3825(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n433), .Q(n26[11]));
    nand g3826(n3476 ,n3450 ,n3460);
    nand g3827(n342 ,n243 ,n274);
    nand g3828(n1639 ,n1231 ,n1232);
    nand g3829(n2683 ,n2658 ,n2667);
    nand g3830(n3178 ,n3065 ,n3151);
    nor g3831(n1804 ,n29[11] ,n1779);
    or g3832(n1849 ,n1826 ,n1829);
    nand g3833(n1050 ,n11[3] ,n441);
    xnor g3834(n3633 ,n3845 ,n3829);
    nand g3835(n1224 ,n14[11] ,n466);
    nand g3836(n2181 ,n2155 ,n2122);
    nor g3837(n289 ,n119 ,n246);
    nor g3838(n2390 ,n2357 ,n2389);
    xnor g3839(n233 ,n158 ,n29[10]);
    nand g3840(n2680 ,n2662 ,n2669);
    xnor g3841(n30[6] ,n2678 ,n2690);
    nor g3842(n2301 ,n2112 ,n2270);
    nand g3843(n1201 ,n21[14] ,n471);
    nand g3844(n3575 ,n3513 ,n3574);
    nand g3845(n1703 ,n1295 ,n1294);
    nand g3846(n3086 ,n2869 ,n3026);
    nand g3847(n1450 ,n1073 ,n622);
    dff g3848(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1515), .Q(n22[14]));
    nand g3849(n1474 ,n1106 ,n680);
    nor g3850(n2196 ,n2143 ,n2157);
    nand g3851(n1610 ,n1198 ,n884);
    nand g3852(n3014 ,n2774 ,n2908);
    nand g3853(n503 ,n207 ,n404);
    nand g3854(n755 ,n191 ,n488);
    nand g3855(n862 ,n11[4] ,n478);
    nor g3856(n125 ,n94 ,n29[1]);
    nor g3857(n2534 ,n2430 ,n2494);
    nand g3858(n37 ,n26[4] ,n34);
    nor g3859(n830 ,n15[9] ,n492);
    nand g3860(n688 ,n187 ,n442);
    nand g3861(n1469 ,n933 ,n561);
    nand g3862(n607 ,n179 ,n485);
    nand g3863(n1652 ,n1260 ,n857);
    nand g3864(n1764 ,n1675 ,n1752);
    xor g3865(n187 ,n4[3] ,n29[3]);
    nand g3866(n722 ,n182 ,n480);
    nand g3867(n3498 ,n3444 ,n3483);
    nand g3868(n3531 ,n3488 ,n3521);
    nand g3869(n45 ,n26[8] ,n42);
    not g3870(n3671 ,n3);
    nand g3871(n171 ,n3 ,n106);
    nand g3872(n283 ,n170 ,n193);
    xnor g3873(n1950 ,n1926 ,n1912);
    nand g3874(n2063 ,n1974 ,n2021);
    nand g3875(n1920 ,n27[2] ,n1902);
    nand g3876(n2093 ,n2006 ,n2027);
    nand g3877(n1040 ,n9[1] ,n459);
    xnor g3878(n3401 ,n3314 ,n3270);
    or g3879(n1842 ,n1821 ,n1837);
    nand g3880(n674 ,n191 ,n440);
    nand g3881(n1141 ,n14[7] ,n491);
    nand g3882(n514 ,n182 ,n483);
    nand g3883(n633 ,n181 ,n445);
    nand g3884(n1588 ,n1056 ,n1057);
    dff g3885(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n844), .Q(n26[2]));
    nand g3886(n1833 ,n396 ,n1797);
    or g3887(n48 ,n26[10] ,n46);
    or g3888(n2869 ,n2831 ,n2726);
    nand g3889(n586 ,n188 ,n487);
    nand g3890(n509 ,n186 ,n453);
    nand g3891(n376 ,n277 ,n294);
    nand g3892(n3604 ,n3583 ,n3603);
    nor g3893(n130 ,n26[7] ,n26[8]);
    nand g3894(n1088 ,n16[6] ,n444);
    nand g3895(n3040 ,n2784 ,n2934);
    nor g3896(n2319 ,n2179 ,n2295);
    or g3897(n3404 ,n3322 ,n3368);
    nand g3898(n1393 ,n960 ,n586);
    nand g3899(n1400 ,n967 ,n535);
    nand g3900(n3018 ,n2763 ,n2910);
    nand g3901(n2054 ,n3850 ,n2015);
    nor g3902(n209 ,n27[2] ,n143);
    nand g3903(n3772 ,n3738 ,n3751);
    nor g3904(n2497 ,n2408 ,n2442);
    nand g3905(n292 ,n202 ,n220);
    or g3906(n2897 ,n2818 ,n2827);
    nor g3907(n2392 ,n2376 ,n2391);
    xnor g3908(n3480 ,n3444 ,n3461);
    dff g3909(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n393), .Q(n26[9]));
    nand g3910(n1209 ,n16[13] ,n499);
    nor g3911(n3677 ,n3866 ,n30[5]);
    xnor g3912(n2213 ,n2141 ,n2152);
    nand g3913(n1488 ,n1121 ,n729);
    nand g3914(n2446 ,n2422 ,n2409);
    nor g3915(n2585 ,n2520 ,n2569);
    dff g3916(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1378), .Q(n13[3]));
    nand g3917(n1147 ,n9[14] ,n459);
    nand g3918(n1525 ,n1161 ,n753);
    dff g3919(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1350), .Q(n13[14]));
    nand g3920(n508 ,n184 ,n485);
    nand g3921(n3782 ,n3736 ,n3732);
    nor g3922(n81 ,n60 ,n80);
    xnor g3923(n3444 ,n3389 ,n3331);
    nand g3924(n1356 ,n917 ,n547);
    nor g3925(n3673 ,n3863 ,n30[8]);
    nand g3926(n3066 ,n2880 ,n3027);
    nand g3927(n2554 ,n2533 ,n2530);
    nand g3928(n1320 ,n851 ,n616);
    nand g3929(n306 ,n26[2] ,n247);
    nand g3930(n30[12] ,n2650 ,n2701);
    nor g3931(n3216 ,n3081 ,n3120);
    nand g3932(n1743 ,n1313 ,n1716);
    xnor g3933(n3587 ,n4[7] ,n26[7]);
    nand g3934(n1579 ,n1203 ,n859);
    or g3935(n1794 ,n359 ,n1777);
    nor g3936(n2523 ,n2468 ,n2501);
    nand g3937(n582 ,n179 ,n487);
    or g3938(n3530 ,n3488 ,n3521);
    or g3939(n299 ,n201 ,n240);
    or g3940(n2416 ,n3812 ,n4[2]);
    dff g3941(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n350), .Q(n24[0]));
    nor g3942(n2176 ,n2104 ,n2147);
    nand g3943(n2043 ,n3858 ,n1987);
    xnor g3944(n2990 ,n2835 ,n2803);
    nand g3945(n2917 ,n2728 ,n2791);
    nand g3946(n1078 ,n21[0] ,n471);
    nand g3947(n2914 ,n2742 ,n2804);
    nor g3948(n365 ,n27[0] ,n319);
    xnor g3949(n3859 ,n3639 ,n3659);
    xnor g3950(n2360 ,n2329 ,n2337);
    xnor g3951(n2276 ,n2213 ,n2248);
    nor g3952(n2164 ,n2161 ,n2136);
    nand g3953(n1361 ,n921 ,n551);
    nand g3954(n3743 ,n3830 ,n3684);
    xnor g3955(n2252 ,n2208 ,n2131);
    xnor g3956(n3115 ,n2966 ,n2861);
    nand g3957(n1568 ,n1266 ,n659);
    nand g3958(n2055 ,n3857 ,n1987);
    nand g3959(n982 ,n17[9] ,n484);
    nand g3960(n2223 ,n2109 ,n2193);
    nand g3961(n1994 ,n3856 ,n1964);
    nand g3962(n1335 ,n890 ,n533);
    nand g3963(n3218 ,n3006 ,n3147);
    nor g3964(n2377 ,n2339 ,n2363);
    dff g3965(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n13[15]));
    nor g3966(n465 ,n211 ,n412);
    not g3967(n2806 ,n2805);
    xnor g3968(n3283 ,n3168 ,n3091);
    nand g3969(n3213 ,n3075 ,n3125);
    nand g3970(n564 ,n192 ,n449);
    not g3971(n2780 ,n2779);
    nand g3972(n3762 ,n3694 ,n3710);
    not g3973(n2845 ,n2844);
    nor g3974(n300 ,n201 ,n217);
    not g3975(n2952 ,n2930);
    xnor g3976(n214 ,n156 ,n29[5]);
    nor g3977(n783 ,n9[5] ,n497);
    xnor g3978(n1915 ,n28[2] ,n27[2]);
    nor g3979(n1308 ,n833 ,n774);
    nand g3980(n1192 ,n16[15] ,n499);
    nand g3981(n1188 ,n9[2] ,n459);
    nor g3982(n2544 ,n2534 ,n2511);
    dff g3983(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1465), .Q(n10[12]));
    nand g3984(n2420 ,n3812 ,n4[2]);
    nand g3985(n957 ,n20[6] ,n452);
    nand g3986(n1512 ,n1144 ,n737);
    nand g3987(n1176 ,n12[10] ,n476);
    dff g3988(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1483), .Q(n15[6]));
    nand g3989(n2807 ,n27[4] ,n4[1]);
    xnor g3990(n3809 ,n3623 ,n3669);
    nand g3991(n1761 ,n1663 ,n1753);
    nand g3992(n274 ,n24[4] ,n201);
    dff g3993(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1855), .Q(n5[11]));
    nand g3994(n412 ,n27[3] ,n364);
    nand g3995(n611 ,n179 ,n483);
    nor g3996(n3612 ,n3845 ,n3829);
    xnor g3997(n2963 ,n2791 ,n2728);
    nand g3998(n2850 ,n27[7] ,n4[5]);
    xnor g3999(n3389 ,n3323 ,n3283);
    xnor g4000(n3549 ,n3527 ,n3534);
    nand g4001(n1727 ,n1683 ,n1682);
    nor g4002(n1678 ,n1613 ,n1612);
    xnor g4003(n1892 ,n28[3] ,n89);
    nand g4004(n878 ,n17[0] ,n468);
    nand g4005(n307 ,n1874 ,n245);
    nand g4006(n1649 ,n1017 ,n868);
    nand g4007(n3263 ,n3142 ,n3178);
    or g4008(n133 ,n28[4] ,n1);
    xnor g4009(n2281 ,n2235 ,n2240);
    nand g4010(n2049 ,n3851 ,n2015);
    xnor g4011(n204 ,n95 ,n4[1]);
    nand g4012(n1486 ,n1119 ,n687);
    nand g4013(n617 ,n187 ,n485);
    or g4014(n2878 ,n2744 ,n2810);
    xnor g4015(n2641 ,n2607 ,n2590);
    nand g4016(n2719 ,n28[0] ,n26[5]);
    xnor g4017(n2964 ,n2726 ,n2831);
    nor g4018(n3621 ,n3840 ,n3824);
    nand g4019(n1711 ,n1671 ,n1670);
    nor g4020(n2144 ,n1988 ,n2102);
    nand g4021(n2670 ,n2653 ,n2655);
    nand g4022(n597 ,n188 ,n483);
    nand g4023(n685 ,n189 ,n442);
    nand g4024(n662 ,n190 ,n457);
    nand g4025(n1696 ,n1277 ,n1300);
    xnor g4026(n220 ,n164 ,n29[11]);
    or g4027(n1289 ,n766 ,n802);
    nand g4028(n264 ,n24[6] ,n201);
    nand g4029(n2029 ,n3854 ,n1985);
    nor g4030(n410 ,n28[2] ,n361);
    nor g4031(n1673 ,n1601 ,n1600);
    xnor g4032(n3309 ,n2704 ,n3118);
    or g4033(n3071 ,n3009 ,n3003);
    nand g4034(n1468 ,n1100 ,n722);
    nand g4035(n3737 ,n3822 ,n3684);
    nand g4036(n1539 ,n1175 ,n702);
    nand g4037(n396 ,n5[3] ,n359);
    xnor g4038(n3124 ,n2965 ,n2747);
    dff g4039(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n23[3]));
    nand g4040(n1965 ,n3850 ,n1959);
    nand g4041(n1627 ,n964 ,n1221);
    nor g4042(n1713 ,n1700 ,n1699);
    nand g4043(n3509 ,n3472 ,n3493);
    nand g4044(n85 ,n26[14] ,n84);
    not g4045(n103 ,n29[14]);
    nand g4046(n1437 ,n1043 ,n669);
    nor g4047(n141 ,n28[0] ,n28[3]);
    nand g4048(n2754 ,n28[6] ,n26[0]);
    nand g4049(n1567 ,n1273 ,n673);
    nand g4050(n2437 ,n2417 ,n2414);
    nor g4051(n2184 ,n2146 ,n2132);
    not g4052(n2785 ,n2711);
    nand g4053(n919 ,n21[11] ,n454);
    dff g4054(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1530), .Q(n22[5]));
    nand g4055(n511 ,n191 ,n485);
    xnor g4056(n2203 ,n2124 ,n2126);
    or g4057(n29[11] ,n3779 ,n3771);
    nand g4058(n1578 ,n1033 ,n858);
    nand g4059(n2732 ,n27[3] ,n4[0]);
    nor g4060(n794 ,n22[5] ,n462);
    xnor g4061(n3586 ,n4[6] ,n26[6]);
    nand g4062(n749 ,n180 ,n488);
    nand g4063(n35 ,n26[3] ,n32);
    nand g4064(n1340 ,n894 ,n515);
    not g4065(n482 ,n483);
    xnor g4066(n3631 ,n3835 ,n3819);
    nand g4067(n66 ,n26[3] ,n65);
    nand g4068(n1148 ,n14[3] ,n491);
    xnor g4069(n2688 ,n2669 ,n2662);
    xnor g4070(n2382 ,n2358 ,n2370);
    xnor g4071(n3479 ,n3410 ,n3445);
    nor g4072(n2628 ,n2597 ,n2611);
    nor g4073(n3707 ,n3698 ,n3683);
    nand g4074(n954 ,n20[8] ,n452);
    xnor g4075(n1911 ,n27[4] ,n27[3]);
    nand g4076(n3740 ,n30[4] ,n3699);
    nand g4077(n3054 ,n2891 ,n3017);
    nor g4078(n2516 ,n2425 ,n2495);
    xnor g4079(n3266 ,n3185 ,n3113);
    nand g4080(n2266 ,n2228 ,n2233);
    xnor g4081(n3368 ,n3264 ,n3304);
    or g4082(n2602 ,n2568 ,n2587);
    nand g4083(n346 ,n313 ,n288);
    nand g4084(n1032 ,n15[4] ,n493);
    not g4085(n102 ,n29[9]);
    nor g4086(n780 ,n11[2] ,n479);
    nand g4087(n312 ,n1868 ,n245);
    nand g4088(n2773 ,n27[1] ,n4[2]);
    nand g4089(n669 ,n189 ,n440);
    nand g4090(n2711 ,n27[0] ,n4[3]);
    nand g4091(n1644 ,n1159 ,n905);
    nand g4092(n1584 ,n1052 ,n870);
    not g4093(n468 ,n469);
    nand g4094(n843 ,n330 ,n435);
    nand g4095(n896 ,n23[6] ,n447);
    nand g4096(n3595 ,n3579 ,n3589);
    xnor g4097(n3131 ,n2986 ,n2826);
    nand g4098(n3341 ,n3260 ,n3282);
    nand g4099(n2312 ,n2266 ,n2290);
    nand g4100(n2918 ,n2720 ,n2789);
    dff g4101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n843), .Q(n26[3]));
    nand g4102(n3249 ,n3154 ,n3186);
    nand g4103(n1128 ,n14[14] ,n491);
    xnor g4104(n3126 ,n2976 ,n2852);
    nor g4105(n1282 ,n783 ,n763);
    nor g4106(n2315 ,n2260 ,n2284);
    nor g4107(n3608 ,n3841 ,n3825);
    nand g4108(n704 ,n190 ,n458);
    nand g4109(n3382 ,n3301 ,n3321);
    nand g4110(n3490 ,n3455 ,n3476);
    nand g4111(n1042 ,n22[7] ,n463);
    nor g4112(n2510 ,n2461 ,n2484);
    nand g4113(n3146 ,n3068 ,n3047);
    nor g4114(n390 ,n127 ,n348);
    dff g4115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1404), .Q(n12[10]));
    nor g4116(n2455 ,n2405 ,n2422);
    dff g4117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n402), .Q(n26[1]));
    nand g4118(n1125 ,n15[0] ,n443);
    nand g4119(n2846 ,n28[6] ,n26[2]);
    nand g4120(n1056 ,n15[1] ,n493);
    not g4121(n3277 ,n3276);
    nand g4122(n2617 ,n2565 ,n2601);
    nand g4123(n1542 ,n1183 ,n705);
    nand g4124(n392 ,n124 ,n343);
    xnor g4125(n2974 ,n2723 ,n2816);
    nand g4126(n3693 ,n3865 ,n30[6]);
    nand g4127(n2699 ,n2673 ,n2698);
    nand g4128(n1139 ,n14[8] ,n491);
    nor g4129(n285 ,n118 ,n246);
    nand g4130(n1721 ,n1677 ,n1676);
    nand g4131(n3293 ,n3241 ,n3236);
    nor g4132(n2476 ,n2406 ,n2437);
    nor g4133(n2399 ,n2398 ,n2368);
    nand g4134(n3686 ,n3863 ,n30[8]);
    dff g4135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1460), .Q(n10[14]));
    nand g4136(n1231 ,n21[11] ,n471);
    xnor g4137(n2228 ,n2160 ,n2136);
    xnor g4138(n3098 ,n2999 ,n2830);
    nor g4139(n2582 ,n2538 ,n2557);
    dff g4140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1365), .Q(n21[7]));
    nor g4141(n2460 ,n2407 ,n2420);
    not g4142(n94 ,n1);
    xnor g4143(n3518 ,n3458 ,n3485);
    dff g4144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1416), .Q(n12[6]));
    nor g4145(n1280 ,n796 ,n762);
    nand g4146(n1230 ,n13[6] ,n501);
    xnor g4147(n2304 ,n2258 ,n2197);
    xnor g4148(n3481 ,n3407 ,n3440);
    nor g4149(n286 ,n201 ,n222);
    nor g4150(n2400 ,n2355 ,n2399);
    nor g4151(n139 ,n107 ,n28[3]);
    nand g4152(n557 ,n189 ,n449);
    xnor g4153(n3462 ,n3431 ,n3424);
    xnor g4154(n1961 ,n1947 ,n1900);
    nand g4155(n1002 ,n19[0] ,n482);
    nand g4156(n1440 ,n1049 ,n670);
    nand g4157(n489 ,n141 ,n410);
    nand g4158(n3493 ,n3449 ,n3474);
    xnor g4159(n2263 ,n2205 ,n2132);
    not g4160(n3125 ,n3124);
    not g4161(n3326 ,n3325);
    nor g4162(n2388 ,n2387 ,n2353);
    nand g4163(n2816 ,n27[2] ,n4[5]);
    dff g4164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1531), .Q(n9[11]));
    or g4165(n435 ,n388 ,n390);
    nand g4166(n2792 ,n27[2] ,n4[0]);
    not g4167(n2902 ,n2901);
    nand g4168(n956 ,n12[15] ,n486);
    or g4169(n29[0] ,n3772 ,n3792);
    nand g4170(n1422 ,n999 ,n550);
    nand g4171(n3643 ,n3609 ,n3642);
    dff g4172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1429), .Q(n18[0]));
    nor g4173(n2429 ,n2405 ,n2424);
    nand g4174(n3489 ,n3448 ,n3470);
    xnor g4175(n2541 ,n2504 ,n2449);
    nand g4176(n537 ,n179 ,n449);
    nand g4177(n126 ,n29[2] ,n94);
    nand g4178(n71 ,n26[6] ,n70);
    nand g4179(n339 ,n1875 ,n245);
    nor g4180(n1298 ,n811 ,n810);
    nor g4181(n2353 ,n2318 ,n2332);
    nand g4182(n3760 ,n3826 ,n3684);
    nand g4183(n1993 ,n3857 ,n1960);
    nand g4184(n1054 ,n16[14] ,n444);
    or g4185(n3367 ,n3307 ,n3334);
    nand g4186(n1371 ,n932 ,n559);
    nor g4187(n838 ,n23[8] ,n464);
endmodule
