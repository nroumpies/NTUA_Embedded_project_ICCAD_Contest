module top (n0, n1, n3, n4, n5, n6, n8, n9, n2, n7, n10, n11, n12, n13, n14, n15, n16, n17);
    input n0, n1, n2;
    input [31:0] n3, n4, n5;
    input [3:0] n6, n7;
    input [1:0] n8;
    input [7:0] n9;
    output [3:0] n10;
    output [31:0] n11, n12, n13, n14;
    output [15:0] n15, n16;
    output [7:0] n17;
    wire n0, n1, n2;
    wire [31:0] n3, n4, n5;
    wire [3:0] n6, n7;
    wire [1:0] n8;
    wire [7:0] n9;
    wire [3:0] n10;
    wire [31:0] n11, n12, n13, n14;
    wire [15:0] n15, n16;
    wire [7:0] n17;
    wire [1:0] n18;
    wire [31:0] n19;
    wire [31:0] n20;
    wire [31:0] n21;
    wire [7:0] n22;
    wire [3:0] n23;
    wire [31:0] n24;
    wire [31:0] n25;
    wire [31:0] n26;
    wire [3:0] n27;
    wire [31:0] n28;
    wire [31:0] n29;
    wire [31:0] n30;
    wire [31:0] n31;
    wire [31:0] n32;
    wire [31:0] n33;
    wire [31:0] n34;
    wire [31:0] n35;
    wire [3:0] n36;
    wire n37, n38, n39, n40, n41, n42, n43, n44;
    wire n45, n46, n47, n48, n49, n50, n51, n52;
    wire n53, n54, n55, n56, n57, n58, n59, n60;
    wire n61, n62, n63, n64, n65, n66, n67, n68;
    wire n69, n70, n71, n72, n73, n74, n75, n76;
    wire n77, n78, n79, n80, n81, n82, n83, n84;
    wire n85, n86, n87, n88, n89, n90, n91, n92;
    wire n93, n94, n95, n96, n97, n98, n99, n100;
    wire n101, n102, n103, n104, n105, n106, n107, n108;
    wire n109, n110, n111, n112, n113, n114, n115, n116;
    wire n117, n118, n119, n120, n121, n122, n123, n124;
    wire n125, n126, n127, n128, n129, n130, n131, n132;
    wire n133, n134, n135, n136, n137, n138, n139, n140;
    wire n141, n142, n143, n144, n145, n146, n147, n148;
    wire n149, n150, n151, n152, n153, n154, n155, n156;
    wire n157, n158, n159, n160, n161, n162, n163, n164;
    wire n165, n166, n167, n168, n169, n170, n171, n172;
    wire n173, n174, n175, n176, n177, n178, n179, n180;
    wire n181, n182, n183, n184, n185, n186, n187, n188;
    wire n189, n190, n191, n192, n193, n194, n195, n196;
    wire n197, n198, n199, n200, n201, n202, n203, n204;
    wire n205, n206, n207, n208, n209, n210, n211, n212;
    wire n213, n214, n215, n216, n217, n218, n219, n220;
    wire n221, n222, n223, n224, n225, n226, n227, n228;
    wire n229, n230, n231, n232, n233, n234, n235, n236;
    wire n237, n238, n239, n240, n241, n242, n243, n244;
    wire n245, n246, n247, n248, n249, n250, n251, n252;
    wire n253, n254, n255, n256, n257, n258, n259, n260;
    wire n261, n262, n263, n264, n265, n266, n267, n268;
    wire n269, n270, n271, n272, n273, n274, n275, n276;
    wire n277, n278, n279, n280, n281, n282, n283, n284;
    wire n285, n286, n287, n288, n289, n290, n291, n292;
    wire n293, n294, n295, n296, n297, n298, n299, n300;
    wire n301, n302, n303, n304, n305, n306, n307, n308;
    wire n309, n310, n311, n312, n313, n314, n315, n316;
    wire n317, n318, n319, n320, n321, n322, n323, n324;
    wire n325, n326, n327, n328, n329, n330, n331, n332;
    wire n333, n334, n335, n336, n337, n338, n339, n340;
    wire n341, n342, n343, n344, n345, n346, n347, n348;
    wire n349, n350, n351, n352, n353, n354, n355, n356;
    wire n357, n358, n359, n360, n361, n362, n363, n364;
    wire n365, n366, n367, n368, n369, n370, n371, n372;
    wire n373, n374, n375, n376, n377, n378, n379, n380;
    wire n381, n382, n383, n384, n385, n386, n387, n388;
    wire n389, n390, n391, n392, n393, n394, n395, n396;
    wire n397, n398, n399, n400, n401, n402, n403, n404;
    wire n405, n406, n407, n408, n409, n410, n411, n412;
    wire n413, n414, n415, n416, n417, n418, n419, n420;
    wire n421, n422, n423, n424, n425, n426, n427, n428;
    wire n429, n430, n431, n432, n433, n434, n435, n436;
    wire n437, n438, n439, n440, n441, n442, n443, n444;
    wire n445, n446, n447, n448, n449, n450, n451, n452;
    wire n453, n454, n455, n456, n457, n458, n459, n460;
    wire n461, n462, n463, n464, n465, n466, n467, n468;
    wire n469, n470, n471, n472, n473, n474, n475, n476;
    wire n477, n478, n479, n480, n481, n482, n483, n484;
    wire n485, n486, n487, n488, n489, n490, n491, n492;
    wire n493, n494, n495, n496, n497, n498, n499, n500;
    wire n501, n502, n503, n504, n505, n506, n507, n508;
    wire n509, n510, n511, n512, n513, n514, n515, n516;
    wire n517, n518, n519, n520, n521, n522, n523, n524;
    wire n525, n526, n527, n528, n529, n530, n531, n532;
    wire n533, n534, n535, n536, n537, n538, n539, n540;
    wire n541, n542, n543, n544, n545, n546, n547, n548;
    wire n549, n550, n551, n552, n553, n554, n555, n556;
    wire n557, n558, n559, n560, n561, n562, n563, n564;
    wire n565, n566, n567, n568, n569, n570, n571, n572;
    wire n573, n574, n575, n576, n577, n578, n579, n580;
    wire n581, n582, n583, n584, n585, n586, n587, n588;
    wire n589, n590, n591, n592, n593, n594, n595, n596;
    wire n597, n598, n599, n600, n601, n602, n603, n604;
    wire n605, n606, n607, n608, n609, n610, n611, n612;
    wire n613, n614, n615, n616, n617, n618, n619, n620;
    wire n621, n622, n623, n624, n625, n626, n627, n628;
    wire n629, n630, n631, n632, n633, n634, n635, n636;
    wire n637, n638, n639, n640, n641, n642, n643, n644;
    wire n645, n646, n647, n648, n649, n650, n651, n652;
    wire n653, n654, n655, n656, n657, n658, n659, n660;
    wire n661, n662, n663, n664, n665, n666, n667, n668;
    wire n669, n670, n671, n672, n673, n674, n675, n676;
    wire n677, n678, n679, n680, n681, n682, n683, n684;
    wire n685, n686, n687, n688, n689, n690, n691, n692;
    wire n693, n694, n695, n696, n697, n698, n699, n700;
    wire n701, n702, n703, n704, n705, n706, n707, n708;
    wire n709, n710, n711, n712, n713, n714, n715, n716;
    wire n717, n718, n719, n720, n721, n722, n723, n724;
    wire n725, n726, n727, n728, n729, n730, n731, n732;
    wire n733, n734, n735, n736, n737, n738, n739, n740;
    wire n741, n742, n743, n744, n745, n746, n747, n748;
    wire n749, n750, n751, n752, n753, n754, n755, n756;
    wire n757, n758, n759, n760, n761, n762, n763, n764;
    wire n765, n766, n767, n768, n769, n770, n771, n772;
    wire n773, n774, n775, n776, n777, n778, n779, n780;
    wire n781, n782, n783, n784, n785, n786, n787, n788;
    wire n789, n790, n791, n792, n793, n794, n795, n796;
    wire n797, n798, n799, n800, n801, n802, n803, n804;
    wire n805, n806, n807, n808, n809, n810, n811, n812;
    wire n813, n814, n815, n816, n817, n818, n819, n820;
    wire n821, n822, n823, n824, n825, n826, n827, n828;
    wire n829, n830, n831, n832, n833, n834, n835, n836;
    wire n837, n838, n839, n840, n841, n842, n843, n844;
    wire n845, n846, n847, n848, n849, n850, n851, n852;
    wire n853, n854, n855, n856, n857, n858, n859, n860;
    wire n861, n862, n863, n864, n865, n866, n867, n868;
    wire n869, n870, n871, n872, n873, n874, n875, n876;
    wire n877, n878, n879, n880, n881, n882, n883, n884;
    wire n885, n886, n887, n888, n889, n890, n891, n892;
    wire n893, n894, n895, n896, n897, n898, n899, n900;
    wire n901, n902, n903, n904, n905, n906, n907, n908;
    wire n909, n910, n911, n912, n913, n914, n915, n916;
    wire n917, n918, n919, n920, n921, n922, n923, n924;
    wire n925, n926, n927, n928, n929, n930, n931, n932;
    wire n933, n934, n935, n936, n937, n938, n939, n940;
    wire n941, n942, n943, n944, n945, n946, n947, n948;
    wire n949, n950, n951, n952, n953, n954, n955, n956;
    wire n957, n958, n959, n960, n961, n962, n963, n964;
    wire n965, n966, n967, n968, n969, n970, n971, n972;
    wire n973, n974, n975, n976, n977, n978, n979, n980;
    wire n981, n982, n983, n984, n985, n986, n987, n988;
    wire n989, n990, n991, n992, n993, n994, n995, n996;
    wire n997, n998, n999, n1000, n1001, n1002, n1003, n1004;
    wire n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012;
    wire n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
    wire n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
    wire n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
    wire n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044;
    wire n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
    wire n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060;
    wire n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068;
    wire n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076;
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084;
    wire n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092;
    wire n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100;
    wire n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108;
    wire n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116;
    wire n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124;
    wire n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132;
    wire n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140;
    wire n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148;
    wire n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156;
    wire n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164;
    wire n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172;
    wire n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180;
    wire n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188;
    wire n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196;
    wire n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204;
    wire n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
    wire n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220;
    wire n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228;
    wire n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236;
    wire n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244;
    wire n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252;
    wire n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260;
    wire n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268;
    wire n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276;
    wire n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284;
    wire n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292;
    wire n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300;
    wire n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308;
    wire n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;
    wire n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;
    wire n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332;
    wire n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340;
    wire n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348;
    wire n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356;
    wire n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364;
    wire n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372;
    wire n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380;
    wire n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388;
    wire n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;
    wire n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404;
    wire n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412;
    wire n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;
    wire n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428;
    wire n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436;
    wire n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444;
    wire n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452;
    wire n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;
    wire n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468;
    wire n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476;
    wire n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
    wire n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492;
    wire n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500;
    wire n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508;
    wire n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516;
    wire n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524;
    wire n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532;
    wire n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540;
    wire n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548;
    wire n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556;
    wire n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564;
    wire n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572;
    wire n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580;
    wire n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588;
    wire n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596;
    wire n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604;
    wire n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612;
    wire n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620;
    wire n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628;
    wire n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636;
    wire n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644;
    wire n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652;
    wire n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660;
    wire n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668;
    wire n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676;
    wire n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684;
    wire n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692;
    wire n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700;
    wire n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708;
    wire n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716;
    wire n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724;
    wire n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732;
    wire n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740;
    wire n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748;
    wire n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756;
    wire n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764;
    wire n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772;
    wire n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780;
    wire n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788;
    wire n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796;
    wire n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804;
    wire n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812;
    wire n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820;
    wire n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828;
    wire n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836;
    wire n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844;
    wire n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852;
    wire n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860;
    wire n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868;
    wire n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876;
    wire n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884;
    wire n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892;
    wire n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900;
    wire n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908;
    wire n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916;
    wire n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924;
    wire n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932;
    wire n1933;
    nand g0(n172 ,n21[28] ,n24[28]);
    dff g1(.RN(n1), .SN(1'b1), .CK(n0), .D(n1485), .Q(n28[19]));
    or g2(n469 ,n328 ,n351);
    dff g3(.RN(n1), .SN(1'b1), .CK(n0), .D(n1705), .Q(n21[0]));
    nand g4(n158 ,n22[5] ,n32[5]);
    nand g5(n1429 ,n168 ,n368);
    nand g6(n1906 ,n1902 ,n1876);
    nand g7(n1108 ,n33[21] ,n355);
    nand g8(n1296 ,n624 ,n485);
    not g9(n350 ,n52);
    nand g10(n1125 ,n28[16] ,n46);
    nand g11(n1765 ,n1269 ,n1718);
    dff g12(.RN(n1), .SN(1'b1), .CK(n0), .D(n1609), .Q(n33[25]));
    nand g13(n153 ,n27[0] ,n27[1]);
    or g14(n1919 ,n1904 ,n1909);
    nand g15(n590 ,n21[26] ,n52);
    nand g16(n1515 ,n844 ,n1182);
    nand g17(n1681 ,n1244 ,n936);
    nand g18(n1374 ,n1088 ,n391);
    nand g19(n1777 ,n1228 ,n1641);
    nand g20(n1533 ,n219 ,n463);
    nand g21(n1475 ,n1114 ,n593);
    nand g22(n1447 ,n730 ,n1085);
    nor g23(n1837 ,n27[0] ,n1517);
    nand g24(n233 ,n31[15] ,n34[15]);
    nand g25(n1330 ,n1018 ,n436);
    nor g26(n478 ,n66 ,n50);
    xnor g27(n252 ,n29[29] ,n30[29]);
    nor g28(n86 ,n29[0] ,n30[0]);
    nand g29(n1204 ,n30[13] ,n351);
    dff g30(.RN(n1), .SN(1'b1), .CK(n0), .D(n1529), .Q(n26[10]));
    nand g31(n160 ,n30[2] ,n23[2]);
    not g32(n345 ,n44);
    nand g33(n1059 ,n26[4] ,n45);
    nand g34(n1211 ,n35[21] ,n346);
    or g35(n822 ,n308 ,n345);
    nand g36(n679 ,n11[29] ,n50);
    nand g37(n726 ,n35[20] ,n356);
    dff g38(.RN(n1), .SN(1'b1), .CK(n0), .D(n1370), .Q(n32[25]));
    nand g39(n722 ,n11[0] ,n345);
    nand g40(n1658 ,n1231 ,n914);
    nand g41(n1746 ,n187 ,n445);
    nand g42(n669 ,n33[18] ,n49);
    nand g43(n230 ,n26[25] ,n33[21]);
    nand g44(n812 ,n35[4] ,n356);
    nand g45(n1343 ,n972 ,n504);
    nor g46(n127 ,n28[16] ,n32[16]);
    nand g47(n1814 ,n1098 ,n1458);
    nand g48(n173 ,n21[27] ,n24[27]);
    dff g49(.RN(n1), .SN(1'b1), .CK(n0), .D(n1556), .Q(n34[19]));
    dff g50(.RN(n1), .SN(1'b1), .CK(n0), .D(n1749), .Q(n13[3]));
    dff g51(.RN(n1), .SN(1'b1), .CK(n0), .D(n1685), .Q(n22[0]));
    nand g52(n1183 ,n30[22] ,n351);
    nor g53(n88 ,n26[7] ,n33[3]);
    xnor g54(n282 ,n26[17] ,n33[13]);
    nand g55(n1245 ,n24[17] ,n51);
    nand g56(n1155 ,n30[31] ,n54);
    nand g57(n1468 ,n1110 ,n589);
    nand g58(n1909 ,n1894 ,n1877);
    nand g59(n1150 ,n28[1] ,n46);
    buf g60(n12[27], n11[27]);
    nand g61(n1213 ,n30[10] ,n47);
    nand g62(n1639 ,n648 ,n889);
    nor g63(n54 ,n153 ,n37);
    dff g64(.RN(n1), .SN(1'b1), .CK(n0), .D(n1755), .Q(n13[12]));
    nand g65(n1060 ,n26[3] ,n45);
    nand g66(n1167 ,n30[27] ,n351);
    nand g67(n1333 ,n800 ,n455);
    dff g68(.RN(n1), .SN(1'b1), .CK(n0), .D(n1468), .Q(n28[27]));
    buf g69(n12[24], n11[24]);
    nand g70(n564 ,n22[4] ,n347);
    nand g71(n1149 ,n33[10] ,n55);
    nand g72(n942 ,n9[6] ,n349);
    xnor g73(n313 ,n36[2] ,n33[30]);
    nand g74(n1832 ,n1023 ,n1392);
    nor g75(n132 ,n30[2] ,n23[2]);
    nand g76(n1805 ,n770 ,n1500);
    nand g77(n1826 ,n1071 ,n1443);
    nand g78(n1217 ,n35[17] ,n45);
    not g79(n1870 ,n24[17]);
    dff g80(.RN(n1), .SN(1'b1), .CK(n0), .D(n1318), .Q(n31[30]));
    nand g81(n793 ,n35[19] ,n42);
    dff g82(.RN(n1), .SN(1'b1), .CK(n0), .D(n1541), .Q(n34[28]));
    nand g83(n1528 ,n218 ,n458);
    nor g84(n62 ,n21[9] ,n24[9]);
    dff g85(.RN(n1), .SN(1'b1), .CK(n0), .D(n1544), .Q(n34[26]));
    dff g86(.RN(n1), .SN(1'b1), .CK(n0), .D(n1593), .Q(n26[4]));
    nand g87(n1021 ,n26[31] ,n346);
    dff g88(.RN(n1), .SN(1'b1), .CK(n0), .D(n1354), .Q(n13[15]));
    nor g89(n108 ,n21[28] ,n24[28]);
    nand g90(n1191 ,n30[19] ,n48);
    dff g91(.RN(n1), .SN(1'b1), .CK(n0), .D(n1484), .Q(n28[20]));
    dff g92(.RN(n1), .SN(1'b1), .CK(n0), .D(n1412), .Q(n15[1]));
    dff g93(.RN(n1), .SN(1'b1), .CK(n0), .D(n1340), .Q(n33[7]));
    xnor g94(n317 ,n21[2] ,n24[2]);
    nand g95(n1697 ,n208 ,n496);
    nand g96(n956 ,n5[5] ,n349);
    nand g97(n1382 ,n1229 ,n480);
    nand g98(n1428 ,n710 ,n1053);
    nand g99(n1585 ,n1188 ,n849);
    nand g100(n580 ,n21[1] ,n348);
    nand g101(n657 ,n21[5] ,n51);
    nand g102(n861 ,n34[0] ,n353);
    xnor g103(n259 ,n29[20] ,n30[20]);
    dff g104(.RN(n1), .SN(1'b1), .CK(n0), .D(n1297), .Q(n30[0]));
    dff g105(.RN(n1), .SN(1'b1), .CK(n0), .D(n1605), .Q(n33[27]));
    nand g106(n601 ,n21[15] ,n52);
    dff g107(.RN(n1), .SN(1'b1), .CK(n0), .D(n1564), .Q(n34[15]));
    nand g108(n866 ,n32[14] ,n53);
    nand g109(n1896 ,n21[11] ,n21[10]);
    nand g110(n1098 ,n32[13] ,n46);
    nand g111(n985 ,n35[28] ,n356);
    nand g112(n791 ,n32[22] ,n53);
    dff g113(.RN(n1), .SN(1'b1), .CK(n0), .D(n1472), .Q(n26[21]));
    dff g114(.RN(n1), .SN(1'b1), .CK(n0), .D(n1686), .Q(n24[15]));
    dff g115(.RN(n1), .SN(1'b1), .CK(n0), .D(n1582), .Q(n21[23]));
    nand g116(n1097 ,n28[31] ,n46);
    xnor g117(n308 ,n33[1] ,n26[5]);
    nand g118(n974 ,n13[29] ,n345);
    nor g119(n346 ,n40 ,n38);
    nand g120(n1040 ,n26[17] ,n346);
    nand g121(n1653 ,n962 ,n666);
    buf g122(n14[28], n12[28]);
    buf g123(n16[5], n15[1]);
    nand g124(n1146 ,n33[12] ,n55);
    not g125(n352 ,n54);
    dff g126(.RN(n1), .SN(1'b1), .CK(n0), .D(n1754), .Q(n13[10]));
    nand g127(n952 ,n4[0] ,n43);
    nand g128(n1176 ,n30[24] ,n48);
    nand g129(n1196 ,n30[16] ,n351);
    nand g130(n1339 ,n667 ,n822);
    nand g131(n611 ,n21[5] ,n52);
    nand g132(n1717 ,n969 ,n555);
    nand g133(n702 ,n26[31] ,n354);
    nor g134(n387 ,n63 ,n46);
    or g135(n1933 ,n1932 ,n1931);
    dff g136(.RN(n1), .SN(1'b1), .CK(n0), .D(n1768), .Q(n29[29]));
    not g137(n44 ,n50);
    nand g138(n194 ,n26[29] ,n33[25]);
    nand g139(n190 ,n21[21] ,n24[21]);
    nand g140(n1557 ,n1167 ,n832);
    xnor g141(n341 ,n28[15] ,n32[15]);
    nand g142(n1140 ,n28[7] ,n350);
    xnor g143(n289 ,n26[22] ,n33[18]);
    nand g144(n1472 ,n739 ,n1108);
    nand g145(n222 ,n31[5] ,n34[5]);
    nand g146(n1353 ,n993 ,n522);
    nor g147(n70 ,n31[21] ,n34[21]);
    nor g148(n498 ,n117 ,n47);
    or g149(n532 ,n243 ,n49);
    nand g150(n1288 ,n203 ,n443);
    or g151(n460 ,n272 ,n356);
    nand g152(n1619 ,n1213 ,n875);
    nor g153(n546 ,n86 ,n353);
    nand g154(n1424 ,n703 ,n1047);
    xnor g155(n280 ,n31[10] ,n34[10]);
    nand g156(n606 ,n21[10] ,n52);
    nand g157(n1762 ,n975 ,n1722);
    dff g158(.RN(n1), .SN(1'b1), .CK(n0), .D(n1790), .Q(n35[12]));
    nand g159(n632 ,n21[16] ,n51);
    nand g160(n1558 ,n835 ,n1168);
    nand g161(n1616 ,n1210 ,n695);
    dff g162(.RN(n1), .SN(1'b1), .CK(n0), .D(n1597), .Q(n33[31]));
    nand g163(n1747 ,n887 ,n1222);
    nand g164(n156 ,n22[7] ,n32[7]);
    dff g165(.RN(n1), .SN(1'b1), .CK(n0), .D(n1557), .Q(n30[27]));
    nand g166(n1932 ,n1928 ,n1929);
    nand g167(n911 ,n26[1] ,n354);
    dff g168(.RN(n1), .SN(1'b1), .CK(n0), .D(n1712), .Q(n18[1]));
    nand g169(n1514 ,n191 ,n506);
    nand g170(n761 ,n31[25] ,n352);
    nand g171(n1545 ,n1187 ,n766);
    nand g172(n1924 ,n1912 ,n1916);
    nand g173(n1501 ,n1135 ,n606);
    nand g174(n1512 ,n226 ,n503);
    nand g175(n1466 ,n736 ,n1094);
    nand g176(n609 ,n21[7] ,n52);
    nand g177(n957 ,n5[4] ,n349);
    dff g178(.RN(n1), .SN(1'b1), .CK(n0), .D(n1424), .Q(n11[12]));
    nand g179(n1228 ,n30[5] ,n47);
    buf g180(n14[15], n11[15]);
    nand g181(n1559 ,n1285 ,n1171);
    dff g182(.RN(n1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n13[14]));
    xnor g183(n322 ,n21[18] ,n24[18]);
    dff g184(.RN(n1), .SN(1'b1), .CK(n0), .D(n1447), .Q(n26[25]));
    dff g185(.RN(n1), .SN(1'b1), .CK(n0), .D(n1822), .Q(n32[22]));
    nand g186(n1269 ,n29[27] ,n48);
    nand g187(n241 ,n29[28] ,n30[28]);
    not g188(n1868 ,n21[14]);
    nand g189(n887 ,n33[13] ,n49);
    nor g190(n421 ,n93 ,n352);
    nor g191(n526 ,n64 ,n50);
    dff g192(.RN(n1), .SN(1'b1), .CK(n0), .D(n1507), .Q(n28[6]));
    nand g193(n1845 ,n150 ,n1841);
    nand g194(n1700 ,n1258 ,n955);
    xnor g195(n285 ,n26[30] ,n33[26]);
    nand g196(n915 ,n9[7] ,n349);
    nor g197(n139 ,n30[3] ,n23[3]);
    nand g198(n1483 ,n578 ,n748);
    dff g199(.RN(n1), .SN(1'b1), .CK(n0), .D(n1489), .Q(n26[17]));
    dff g200(.RN(n1), .SN(1'b1), .CK(n0), .D(n1801), .Q(n35[26]));
    nand g201(n1847 ,n147 ,n1844);
    nand g202(n1791 ,n799 ,n1525);
    nand g203(n859 ,n32[29] ,n53);
    nand g204(n1885 ,n21[15] ,n1868);
    or g205(n514 ,n286 ,n50);
    dff g206(.RN(n1), .SN(1'b1), .CK(n0), .D(n1426), .Q(n11[10]));
    nand g207(n1118 ,n28[21] ,n350);
    nand g208(n867 ,n34[29] ,n353);
    nor g209(n368 ,n123 ,n351);
    nor g210(n101 ,n28[13] ,n32[13]);
    dff g211(.RN(n1), .SN(1'b1), .CK(n0), .D(n1676), .Q(n21[5]));
    nand g212(n1770 ,n1251 ,n1690);
    nand g213(n615 ,n32[7] ,n46);
    nor g214(n401 ,n82 ,n46);
    nor g215(n140 ,n26[14] ,n33[10]);
    nand g216(n1614 ,n658 ,n711);
    nand g217(n1181 ,n30[23] ,n351);
    nor g218(n68 ,n22[5] ,n35[5]);
    dff g219(.RN(n1), .SN(1'b1), .CK(n0), .D(n1692), .Q(n21[1]));
    dff g220(.RN(n1), .SN(1'b1), .CK(n0), .D(n1680), .Q(n24[19]));
    nor g221(n394 ,n110 ,n42);
    nor g222(n131 ,n31[4] ,n34[4]);
    nor g223(n144 ,n28[18] ,n32[18]);
    nand g224(n951 ,n10[0] ,n356);
    nand g225(n987 ,n35[31] ,n356);
    dff g226(.RN(n1), .SN(1'b1), .CK(n0), .D(n1494), .Q(n28[15]));
    nand g227(n1718 ,n225 ,n502);
    buf g228(n12[5], n11[5]);
    or g229(n381 ,n336 ,n46);
    nand g230(n1753 ,n1283 ,n1734);
    nand g231(n1234 ,n24[27] ,n348);
    or g232(n414 ,n267 ,n42);
    nand g233(n1128 ,n33[16] ,n55);
    nand g234(n1164 ,n30[29] ,n351);
    dff g235(.RN(n1), .SN(1'b1), .CK(n0), .D(n1689), .Q(n24[13]));
    dff g236(.RN(n1), .SN(1'b1), .CK(n0), .D(n1604), .Q(n21[19]));
    dff g237(.RN(n1), .SN(1'b1), .CK(n0), .D(n1640), .Q(n33[8]));
    or g238(n488 ,n17[1] ,n357);
    nand g239(n621 ,n32[1] ,n350);
    nor g240(n91 ,n22[5] ,n32[5]);
    nand g241(n1931 ,n1930 ,n1927);
    not g242(n1853 ,n24[23]);
    xnor g243(n298 ,n31[14] ,n34[14]);
    nand g244(n1711 ,n1267 ,n961);
    dff g245(.RN(n1), .SN(1'b1), .CK(n0), .D(n1369), .Q(n29[4]));
    xnor g246(n300 ,n21[16] ,n24[16]);
    nand g247(n240 ,n26[8] ,n33[4]);
    nand g248(n700 ,n11[14] ,n49);
    nand g249(n1086 ,n32[20] ,n350);
    nand g250(n1308 ,n798 ,n453);
    nand g251(n1828 ,n1055 ,n1429);
    xnor g252(n306 ,n32[4] ,n28[4]);
    nor g253(n99 ,n27[0] ,n27[1]);
    nand g254(n1154 ,n30[15] ,n54);
    nand g255(n781 ,n35[30] ,n356);
    nand g256(n1804 ,n978 ,n1509);
    nand g257(n1366 ,n1065 ,n467);
    nand g258(n576 ,n23[2] ,n51);
    nand g259(n1719 ,n971 ,n552);
    nand g260(n839 ,n34[14] ,n353);
    nand g261(n964 ,n8[0] ,n43);
    buf g262(n14[18], n11[18]);
    xor g263(n19[6] ,n21[6] ,n22[6]);
    nand g264(n1133 ,n28[11] ,n350);
    nand g265(n1504 ,n1139 ,n608);
    nand g266(n991 ,n13[17] ,n49);
    dff g267(.RN(n1), .SN(1'b1), .CK(n0), .D(n1766), .Q(n29[28]));
    nand g268(n1272 ,n29[26] ,n48);
    nand g269(n681 ,n11[27] ,n345);
    dff g270(.RN(n1), .SN(1'b1), .CK(n0), .D(n1329), .Q(n31[15]));
    nand g271(n778 ,n26[13] ,n354);
    nand g272(n1690 ,n210 ,n474);
    nand g273(n1324 ,n767 ,n427);
    dff g274(.RN(n1), .SN(1'b1), .CK(n0), .D(n1782), .Q(n31[0]));
    nand g275(n1347 ,n977 ,n510);
    dff g276(.RN(n1), .SN(1'b1), .CK(n0), .D(n1607), .Q(n33[26]));
    dff g277(.RN(n1), .SN(1'b1), .CK(n0), .D(n1808), .Q(n31[28]));
    nor g278(n539 ,n127 ,n351);
    nand g279(n1549 ,n1164 ,n859);
    nand g280(n342 ,n7[0] ,n154);
    xnor g281(n320 ,n21[3] ,n23[3]);
    buf g282(n14[29], n12[29]);
    nand g283(n1683 ,n1245 ,n938);
    nand g284(n1081 ,n29[3] ,n48);
    nor g285(n365 ,n101 ,n47);
    nand g286(n1691 ,n1250 ,n901);
    nand g287(n1745 ,n782 ,n1146);
    dff g288(.RN(n1), .SN(1'b1), .CK(n0), .D(n1555), .Q(n34[20]));
    nand g289(n1776 ,n899 ,n1643);
    xnor g290(n247 ,n26[21] ,n33[17]);
    nand g291(n1617 ,n684 ,n1211);
    dff g292(.RN(n1), .SN(1'b1), .CK(n0), .D(n1666), .Q(n24[27]));
    dff g293(.RN(n1), .SN(1'b1), .CK(n0), .D(n1394), .Q(n12[29]));
    nand g294(n640 ,n21[27] ,n348);
    nand g295(n1624 ,n755 ,n1217);
    nand g296(n1897 ,n20[3] ,n20[2]);
    nor g297(n118 ,n31[12] ,n34[12]);
    dff g298(.RN(n1), .SN(1'b1), .CK(n0), .D(n1804), .Q(n35[29]));
    nand g299(n754 ,n31[28] ,n352);
    dff g300(.RN(n1), .SN(1'b1), .CK(n0), .D(n1636), .Q(n33[10]));
    dff g301(.RN(n1), .SN(1'b1), .CK(n0), .D(n1575), .Q(n34[25]));
    nand g302(n1326 ,n773 ,n431);
    dff g303(.RN(n1), .SN(1'b1), .CK(n0), .D(n1398), .Q(n11[30]));
    dff g304(.RN(n1), .SN(1'b1), .CK(n0), .D(n1551), .Q(n21[28]));
    nand g305(n1444 ,n173 ,n378);
    nand g306(n1073 ,n32[27] ,n350);
    nand g307(n947 ,n5[11] ,n43);
    not g308(n1863 ,n24[24]);
    xnor g309(n286 ,n26[27] ,n33[23]);
    dff g310(.RN(n1), .SN(1'b1), .CK(n0), .D(n1401), .Q(n15[3]));
    nand g311(n844 ,n34[10] ,n353);
    nand g312(n1632 ,n156 ,n500);
    nor g313(n446 ,n136 ,n353);
    nand g314(n843 ,n35[26] ,n42);
    nor g315(n1912 ,n1898 ,n1882);
    nand g316(n779 ,n31[15] ,n352);
    dff g317(.RN(n1), .SN(1'b1), .CK(n0), .D(n1672), .Q(n24[23]));
    xnor g318(n318 ,n21[1] ,n24[1]);
    nand g319(n1220 ,n35[14] ,n45);
    xnor g320(n243 ,n26[13] ,n33[9]);
    nand g321(n1491 ,n211 ,n421);
    xnor g322(n262 ,n29[16] ,n30[16]);
    dff g323(.RN(n1), .SN(1'b1), .CK(n0), .D(n1310), .Q(n35[8]));
    not g324(n360 ,n359);
    nand g325(n1400 ,n679 ,n628);
    nand g326(n1355 ,n997 ,n367);
    nand g327(n854 ,n34[27] ,n352);
    nand g328(n685 ,n11[25] ,n344);
    dff g329(.RN(n1), .SN(1'b1), .CK(n0), .D(n1815), .Q(n32[14]));
    dff g330(.RN(n1), .SN(1'b1), .CK(n0), .D(n1747), .Q(n33[13]));
    nand g331(n801 ,n26[10] ,n354);
    nand g332(n1318 ,n752 ,n417);
    nand g333(n873 ,n34[30] ,n353);
    nor g334(n75 ,n28[22] ,n32[22]);
    nand g335(n1302 ,n967 ,n438);
    nand g336(n745 ,n26[19] ,n354);
    nand g337(n1809 ,n622 ,n1477);
    buf g338(n14[23], n11[23]);
    dff g339(.RN(n1), .SN(1'b1), .CK(n0), .D(n1376), .Q(n32[17]));
    or g340(n374 ,n247 ,n49);
    nor g341(n543 ,n88 ,n50);
    nand g342(n1560 ,n1159 ,n827);
    nor g343(n90 ,n31[29] ,n34[29]);
    dff g344(.RN(n1), .SN(1'b1), .CK(n0), .D(n1716), .Q(n14[2]));
    dff g345(.RN(n1), .SN(1'b1), .CK(n0), .D(n1694), .Q(n21[2]));
    xnor g346(n270 ,n28[17] ,n32[17]);
    nand g347(n1435 ,n716 ,n1060);
    nor g348(n95 ,n29[23] ,n30[23]);
    dff g349(.RN(n1), .SN(1'b1), .CK(n0), .D(n1309), .Q(n35[9]));
    nand g350(n1672 ,n1238 ,n926);
    nand g351(n1023 ,n29[14] ,n48);
    dff g352(.RN(n1), .SN(1'b1), .CK(n0), .D(n1567), .Q(n26[7]));
    dff g353(.RN(n1), .SN(1'b1), .CK(n0), .D(n1817), .Q(n32[15]));
    or g354(n433 ,n262 ,n352);
    nand g355(n225 ,n28[27] ,n32[27]);
    nand g356(n573 ,n18[1] ,n361);
    nand g357(n733 ,n33[30] ,n50);
    nand g358(n1380 ,n1148 ,n444);
    dff g359(.RN(n1), .SN(1'b1), .CK(n0), .D(n1385), .Q(n29[23]));
    nor g360(n1927 ,n1921 ,n1919);
    dff g361(.RN(n1), .SN(1'b1), .CK(n0), .D(n1626), .Q(n30[8]));
    nand g362(n1506 ,n1140 ,n609);
    nand g363(n1044 ,n26[15] ,n346);
    dff g364(.RN(n1), .SN(1'b1), .CK(n0), .D(n1348), .Q(n13[23]));
    nand g365(n1531 ,n216 ,n461);
    nand g366(n1193 ,n30[27] ,n54);
    dff g367(.RN(n1), .SN(1'b1), .CK(n0), .D(n1843), .Q(n28[1]));
    buf g368(n14[24], n11[24]);
    nor g369(n130 ,n31[6] ,n34[6]);
    buf g370(n12[20], n11[20]);
    nand g371(n1016 ,n35[17] ,n356);
    nand g372(n1291 ,n618 ,n408);
    dff g373(.RN(n1), .SN(1'b1), .CK(n0), .D(n1307), .Q(n35[17]));
    nand g374(n1589 ,n1191 ,n850);
    nand g375(n966 ,n14[3] ,n50);
    or g376(n476 ,n245 ,n351);
    nand g377(n1151 ,n33[9] ,n55);
    nand g378(n769 ,n31[20] ,n352);
    nand g379(n981 ,n13[24] ,n345);
    xnor g380(n276 ,n29[14] ,n30[14]);
    dff g381(.RN(n1), .SN(1'b1), .CK(n0), .D(n1823), .Q(n32[26]));
    nand g382(n751 ,n26[18] ,n354);
    nand g383(n1276 ,n29[24] ,n47);
    nand g384(n1802 ,n959 ,n1510);
    nand g385(n1174 ,n30[25] ,n351);
    dff g386(.RN(n1), .SN(1'b1), .CK(n0), .D(n1720), .Q(n25[30]));
    nand g387(n1688 ,n1248 ,n943);
    nand g388(n642 ,n21[22] ,n348);
    nand g389(n1496 ,n196 ,n425);
    nand g390(n1571 ,n786 ,n1180);
    nand g391(n898 ,n4[11] ,n349);
    nor g392(n486 ,n129 ,n48);
    dff g393(.RN(n1), .SN(1'b1), .CK(n0), .D(n1439), .Q(n11[0]));
    nand g394(n1231 ,n24[31] ,n51);
    or g395(n520 ,n289 ,n345);
    nor g396(n105 ,n31[26] ,n34[26]);
    nand g397(n195 ,n31[19] ,n34[19]);
    nand g398(n1328 ,n776 ,n433);
    nand g399(n1189 ,n30[5] ,n54);
    dff g400(.RN(n1), .SN(1'b1), .CK(n0), .D(n1497), .Q(n28[13]));
    nand g401(n1502 ,n1137 ,n607);
    nand g402(n673 ,n12[29] ,n49);
    nor g403(n120 ,n28[30] ,n32[30]);
    nand g404(n984 ,n3[28] ,n349);
    dff g405(.RN(n1), .SN(1'b1), .CK(n0), .D(n487), .Q(n17[2]));
    not g406(n48 ,n53);
    nand g407(n1604 ,n633 ,n732);
    nand g408(n553 ,n22[3] ,n346);
    nand g409(n1818 ,n1087 ,n1453);
    nand g410(n169 ,n28[20] ,n32[20]);
    dff g411(.RN(n1), .SN(1'b1), .CK(n0), .D(n1677), .Q(n22[2]));
    nand g412(n630 ,n36[2] ,n45);
    nand g413(n591 ,n21[25] ,n52);
    not g414(n347 ,n43);
    xnor g415(n336 ,n21[25] ,n24[25]);
    xnor g416(n275 ,n31[0] ,n34[0]);
    nand g417(n1584 ,n760 ,n1189);
    nand g418(n1821 ,n1083 ,n1450);
    nor g419(n484 ,n102 ,n50);
    nand g420(n990 ,n13[18] ,n344);
    nand g421(n1327 ,n775 ,n432);
    nand g422(n704 ,n32[12] ,n53);
    dff g423(.RN(n1), .SN(1'b1), .CK(n0), .D(n1691), .Q(n24[12]));
    nand g424(n1323 ,n765 ,n426);
    nand g425(n1643 ,n198 ,n478);
    buf g426(n14[8], n11[8]);
    nand g427(n785 ,n35[25] ,n356);
    nand g428(n1266 ,n24[1] ,n347);
    dff g429(.RN(n1), .SN(1'b1), .CK(n0), .D(n1368), .Q(n32[30]));
    nand g430(n1822 ,n1082 ,n1448);
    nand g431(n680 ,n11[28] ,n345);
    not g432(n58 ,n27[1]);
    buf g433(n14[25], n11[25]);
    nand g434(n1391 ,n671 ,n1021);
    nand g435(n214 ,n22[1] ,n35[1]);
    nand g436(n1307 ,n1016 ,n535);
    nand g437(n1735 ,n1001 ,n661);
    not g438(n50 ,n346);
    nand g439(n1535 ,n175 ,n466);
    dff g440(.RN(n1), .SN(1'b1), .CK(n0), .D(n1553), .Q(n34[21]));
    buf g441(n17[5], 1'b0);
    nand g442(n1566 ,n839 ,n1175);
    nand g443(n1408 ,n688 ,n1032);
    dff g444(.RN(n1), .SN(1'b1), .CK(n0), .D(n1571), .Q(n34[11]));
    nor g445(n385 ,n85 ,n46);
    nand g446(n1687 ,n582 ,n908);
    nand g447(n1438 ,n719 ,n1057);
    dff g448(.RN(n1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n13[29]));
    nor g449(n437 ,n90 ,n356);
    nand g450(n1129 ,n28[13] ,n46);
    nand g451(n1684 ,n1246 ,n891);
    nand g452(n980 ,n33[15] ,n345);
    or g453(n402 ,n301 ,n350);
    xnor g454(n309 ,n36[1] ,n33[29]);
    dff g455(.RN(n1), .SN(1'b1), .CK(n0), .D(n1671), .Q(n22[4]));
    nand g456(n1437 ,n718 ,n1063);
    nand g457(n1002 ,n13[11] ,n49);
    xnor g458(n324 ,n18[1] ,n33[1]);
    dff g459(.RN(n1), .SN(1'b1), .CK(n0), .D(n1589), .Q(n30[19]));
    nand g460(n697 ,n33[23] ,n50);
    buf g461(n15[14], 1'b0);
    nand g462(n1144 ,n33[5] ,n55);
    nand g463(n1299 ,n987 ,n435);
    buf g464(n16[0], n15[8]);
    dff g465(.RN(n1), .SN(1'b1), .CK(n0), .D(n1759), .Q(n13[22]));
    xnor g466(n263 ,n29[15] ,n30[15]);
    dff g467(.RN(n1), .SN(1'b1), .CK(n0), .D(n1473), .Q(n28[25]));
    dff g468(.RN(n1), .SN(1'b1), .CK(n0), .D(n1356), .Q(n13[13]));
    nand g469(n199 ,n29[19] ,n30[19]);
    nand g470(n1705 ,n583 ,n952);
    dff g471(.RN(n1), .SN(1'b1), .CK(n0), .D(n1633), .Q(n21[14]));
    nand g472(n1027 ,n26[27] ,n44);
    nand g473(n649 ,n21[12] ,n51);
    dff g474(.RN(n1), .SN(1'b1), .CK(n0), .D(n1620), .Q(n33[19]));
    nand g475(n711 ,n4[17] ,n349);
    not g476(n1869 ,n24[28]);
    nand g477(n1248 ,n24[14] ,n348);
    nand g478(n1623 ,n632 ,n876);
    nand g479(n1664 ,n1242 ,n932);
    not g480(n59 ,n7[3]);
    nand g481(n1693 ,n1252 ,n947);
    nand g482(n1399 ,n166 ,n365);
    nand g483(n1808 ,n754 ,n1488);
    nand g484(n1904 ,n1879 ,n1878);
    nand g485(n1142 ,n28[6] ,n46);
    nand g486(n176 ,n21[22] ,n24[22]);
    nand g487(n1292 ,n619 ,n410);
    buf g488(n14[22], n11[22]);
    dff g489(.RN(n1), .SN(1'b1), .CK(n0), .D(n1638), .Q(n33[9]));
    nand g490(n1701 ,n1259 ,n956);
    nand g491(n1893 ,n24[20] ,n1857);
    nor g492(n466 ,n126 ,n356);
    nand g493(n1344 ,n973 ,n472);
    nand g494(n1820 ,n1084 ,n1449);
    nand g495(n1169 ,n33[6] ,n355);
    or g496(n536 ,n270 ,n48);
    nand g497(n1722 ,n227 ,n507);
    nand g498(n1223 ,n35[11] ,n44);
    nand g499(n209 ,n29[0] ,n30[0]);
    nand g500(n1100 ,n28[30] ,n350);
    nor g501(n142 ,n26[8] ,n33[4]);
    nand g502(n1224 ,n30[6] ,n47);
    nand g503(n1143 ,n30[9] ,n54);
    nand g504(n1469 ,n741 ,n1115);
    nand g505(n1301 ,n784 ,n377);
    nand g506(n765 ,n31[22] ,n352);
    not g507(n354 ,n55);
    buf g508(n15[12], 1'b0);
    nand g509(n1253 ,n24[10] ,n347);
    not g510(n1857 ,n24[21]);
    nand g511(n1678 ,n1241 ,n918);
    nand g512(n563 ,n22[0] ,n55);
    xnor g513(n274 ,n29[17] ,n30[17]);
    dff g514(.RN(n1), .SN(1'b1), .CK(n0), .D(n1290), .Q(n32[6]));
    nand g515(n883 ,n31[1] ,n352);
    nand g516(n1760 ,n981 ,n1725);
    nand g517(n1676 ,n657 ,n935);
    dff g518(.RN(n1), .SN(1'b1), .CK(n0), .D(n1339), .Q(n13[1]));
    nand g519(n1840 ,n1152 ,n1835);
    nand g520(n1115 ,n33[20] ,n355);
    nand g521(n983 ,n13[22] ,n49);
    nand g522(n1670 ,n1237 ,n919);
    nand g523(n677 ,n11[30] ,n50);
    nand g524(n232 ,n28[22] ,n32[22]);
    nand g525(n1122 ,n28[18] ,n46);
    nand g526(n1654 ,n910 ,n663);
    nand g527(n894 ,n4[12] ,n349);
    nand g528(n750 ,n26[5] ,n354);
    nand g529(n1628 ,n646 ,n884);
    nand g530(n1800 ,n783 ,n1513);
    dff g531(.RN(n1), .SN(1'b1), .CK(n0), .D(n1602), .Q(n33[29]));
    nand g532(n1689 ,n1249 ,n944);
    nand g533(n1275 ,n35[15] ,n44);
    nor g534(n448 ,n122 ,n353);
    nor g535(n87 ,n26[25] ,n33[21]);
    xnor g536(n253 ,n31[3] ,n34[3]);
    nand g537(n831 ,n34[20] ,n352);
    nand g538(n1163 ,n30[23] ,n54);
    nand g539(n1871 ,n24[18] ,n1864);
    dff g540(.RN(n1), .SN(1'b1), .CK(n0), .D(n1683), .Q(n24[17]));
    nor g541(n456 ,n118 ,n356);
    nand g542(n651 ,n21[10] ,n348);
    nand g543(n646 ,n21[15] ,n347);
    nand g544(n869 ,n31[0] ,n41);
    dff g545(.RN(n1), .SN(1'b1), .CK(n0), .D(n1437), .Q(n11[1]));
    dff g546(.RN(n1), .SN(1'b1), .CK(n0), .D(n1475), .Q(n28[23]));
    nand g547(n1786 ,n809 ,n1531);
    dff g548(.RN(n1), .SN(1'b1), .CK(n0), .D(n1304), .Q(n35[23]));
    dff g549(.RN(n1), .SN(1'b1), .CK(n0), .D(n1679), .Q(n21[4]));
    dff g550(.RN(n1), .SN(1'b1), .CK(n0), .D(n1833), .Q(n13[0]));
    nand g551(n236 ,n31[16] ,n34[16]);
    dff g552(.RN(n1), .SN(1'b1), .CK(n0), .D(n1294), .Q(n32[1]));
    nor g553(n454 ,n91 ,n48);
    buf g554(n16[8], n15[4]);
    dff g555(.RN(n1), .SN(1'b1), .CK(n0), .D(n1476), .Q(n28[22]));
    nand g556(n1252 ,n24[11] ,n347);
    dff g557(.RN(n1), .SN(1'b1), .CK(n0), .D(n1560), .Q(n30[26]));
    nand g558(n624 ,n30[2] ,n47);
    nand g559(n1104 ,n32[10] ,n350);
    nand g560(n1537 ,n871 ,n1155);
    nand g561(n1242 ,n24[28] ,n347);
    nand g562(n1707 ,n1263 ,n954);
    xnor g563(n359 ,n7[2] ,n27[2]);
    dff g564(.RN(n1), .SN(1'b1), .CK(n0), .D(n1569), .Q(n30[24]));
    dff g565(.RN(n1), .SN(1'b1), .CK(n0), .D(n1438), .Q(n26[29]));
    xnor g566(n261 ,n28[24] ,n32[24]);
    nand g567(n627 ,n36[3] ,n346);
    nand g568(n1911 ,n1880 ,n1886);
    nand g569(n1572 ,n1181 ,n841);
    nand g570(n155 ,n27[1] ,n27[2]);
    nand g571(n1773 ,n613 ,n1649);
    nand g572(n1371 ,n1079 ,n382);
    nand g573(n655 ,n21[4] ,n51);
    nand g574(n1048 ,n26[11] ,n45);
    nand g575(n976 ,n13[27] ,n345);
    nand g576(n876 ,n4[16] ,n43);
    xnor g577(n271 ,n31[8] ,n34[8]);
    nand g578(n586 ,n21[30] ,n52);
    nand g579(n764 ,n26[14] ,n354);
    nand g580(n847 ,n5[3] ,n43);
    nand g581(n569 ,n22[7] ,n355);
    nand g582(n1369 ,n1075 ,n379);
    nand g583(n1749 ,n1017 ,n1743);
    nand g584(n683 ,n11[26] ,n50);
    nand g585(n1562 ,n818 ,n1172);
    nand g586(n1781 ,n747 ,n1588);
    nand g587(n1105 ,n35[31] ,n44);
    nand g588(n1464 ,n1103 ,n587);
    dff g589(.RN(n1), .SN(1'b1), .CK(n0), .D(n1495), .Q(n28[14]));
    nand g590(n1907 ,n1889 ,n1888);
    nand g591(n747 ,n34[3] ,n353);
    or g592(n417 ,n251 ,n352);
    dff g593(.RN(n1), .SN(1'b1), .CK(n0), .D(n1809), .Q(n32[0]));
    nor g594(n1876 ,n24[31] ,n24[30]);
    buf g595(n12[26], n11[26]);
    dff g596(.RN(n1), .SN(1'b1), .CK(n0), .D(n1463), .Q(n28[28]));
    nor g597(n507 ,n100 ,n50);
    nand g598(n1509 ,n228 ,n437);
    nor g599(n1516 ,n350 ,n549);
    nand g600(n566 ,n22[5] ,n347);
    not g601(n61 ,n27[2]);
    dff g602(.RN(n1), .SN(1'b1), .CK(n0), .D(n1402), .Q(n11[28]));
    dff g603(.RN(n1), .SN(1'b1), .CK(n0), .D(n1470), .Q(n28[26]));
    nor g604(n363 ,n96 ,n49);
    or g605(n370 ,n339 ,n351);
    dff g606(.RN(n1), .SN(1'b1), .CK(n0), .D(n1828), .Q(n29[8]));
    nand g607(n213 ,n22[2] ,n35[2]);
    nand g608(n181 ,n28[0] ,n32[0]);
    nand g609(n605 ,n21[11] ,n52);
    dff g610(.RN(n1), .SN(1'b1), .CK(n0), .D(n1757), .Q(n29[22]));
    nand g611(n815 ,n35[2] ,n356);
    nand g612(n1049 ,n29[9] ,n351);
    dff g613(.RN(n1), .SN(1'b1), .CK(n0), .D(n1731), .Q(n15[10]));
    nand g614(n737 ,n26[22] ,n354);
    nand g615(n979 ,n13[25] ,n50);
    dff g616(.RN(n1), .SN(1'b1), .CK(n0), .D(n1534), .Q(n26[9]));
    nand g617(n1170 ,n30[28] ,n48);
    dff g618(.RN(n1), .SN(1'b1), .CK(n0), .D(n1451), .Q(n26[26]));
    dff g619(.RN(n1), .SN(1'b1), .CK(n0), .D(n1328), .Q(n31[16]));
    nand g620(n1538 ,n631 ,n819);
    dff g621(.RN(n1), .SN(1'b1), .CK(n0), .D(n1292), .Q(n32[3]));
    nand g622(n1565 ,n1174 ,n837);
    dff g623(.RN(n1), .SN(1'b1), .CK(n0), .D(n1352), .Q(n13[17]));
    dff g624(.RN(n1), .SN(1'b1), .CK(n0), .D(n1675), .Q(n24[21]));
    nand g625(n1801 ,n843 ,n1514);
    xnor g626(n273 ,n31[2] ,n34[2]);
    nand g627(n1240 ,n24[21] ,n347);
    dff g628(.RN(n1), .SN(1'b1), .CK(n0), .D(n1423), .Q(n11[13]));
    nand g629(n938 ,n5[17] ,n349);
    nand g630(n1668 ,n566 ,n921);
    or g631(n427 ,n257 ,n41);
    dff g632(.RN(n1), .SN(1'b1), .CK(n0), .D(n1623), .Q(n21[16]));
    buf g633(n14[30], n12[30]);
    dff g634(.RN(n1), .SN(1'b1), .CK(n0), .D(n1332), .Q(n31[7]));
    nand g635(n794 ,n35[18] ,n356);
    buf g636(n15[15], 1'b0);
    nand g637(n1041 ,n33[31] ,n355);
    nand g638(n1675 ,n1240 ,n931);
    nand g639(n1652 ,n653 ,n909);
    nand g640(n1281 ,n28[2] ,n350);
    or g641(n480 ,n326 ,n47);
    buf g642(n12[21], n11[21]);
    nand g643(n989 ,n13[19] ,n49);
    nand g644(n618 ,n32[4] ,n350);
    dff g645(.RN(n1), .SN(1'b1), .CK(n0), .D(n1652), .Q(n21[8]));
    nand g646(n204 ,n28[26] ,n32[26]);
    dff g647(.RN(n1), .SN(1'b1), .CK(n0), .D(n1289), .Q(n32[7]));
    nand g648(n988 ,n13[20] ,n50);
    nor g649(n380 ,n151 ,n46);
    nand g650(n1407 ,n686 ,n1031);
    dff g651(.RN(n1), .SN(1'b1), .CK(n0), .D(n1427), .Q(n11[9]));
    buf g652(n12[17], n11[17]);
    nor g653(n138 ,n28[11] ,n32[11]);
    buf g654(n16[3], n15[11]);
    nor g655(n462 ,n115 ,n42);
    nand g656(n1761 ,n979 ,n1724);
    nand g657(n1042 ,n26[16] ,n45);
    dff g658(.RN(n1), .SN(1'b1), .CK(n0), .D(n1346), .Q(n13[27]));
    xnor g659(n269 ,n29[11] ,n30[11]);
    nand g660(n897 ,n33[7] ,n345);
    nand g661(n1271 ,n25[29] ,n51);
    dff g662(.RN(n1), .SN(1'b1), .CK(n0), .D(n1428), .Q(n11[8]));
    nand g663(n719 ,n26[29] ,n354);
    nand g664(n1165 ,n30[21] ,n54);
    nand g665(n1439 ,n722 ,n1064);
    nor g666(n1916 ,n1896 ,n1875);
    nand g667(n1892 ,n21[27] ,n1856);
    dff g668(.RN(n1), .SN(1'b1), .CK(n0), .D(n1642), .Q(n21[12]));
    nand g669(n1586 ,n851 ,n1190);
    nand g670(n1479 ,n576 ,n744);
    dff g671(.RN(n1), .SN(1'b1), .CK(n0), .D(n1325), .Q(n31[20]));
    nand g672(n1492 ,n1125 ,n600);
    or g673(n544 ,n281 ,n47);
    nand g674(n1126 ,n28[15] ,n350);
    dff g675(.RN(n1), .SN(1'b1), .CK(n0), .D(n1771), .Q(n26[0]));
    nand g676(n1544 ,n825 ,n1161);
    or g677(n408 ,n304 ,n350);
    nor g678(n77 ,n21[20] ,n24[20]);
    nor g679(n64 ,n26[16] ,n33[12]);
    nand g680(n825 ,n34[26] ,n353);
    nand g681(n1702 ,n1145 ,n611);
    nand g682(n1720 ,n1270 ,n965);
    nand g683(n1035 ,n26[21] ,n45);
    nand g684(n1706 ,n1261 ,n847);
    nand g685(n1598 ,n644 ,n858);
    nand g686(n1843 ,n1150 ,n1836);
    or g687(n432 ,n274 ,n353);
    buf g688(n12[0], n11[28]);
    nand g689(n1082 ,n32[22] ,n46);
    nand g690(n1386 ,n1279 ,n521);
    nand g691(n592 ,n21[24] ,n52);
    not g692(n355 ,n354);
    nand g693(n1409 ,n689 ,n1034);
    nand g694(n1592 ,n1192 ,n853);
    nand g695(n901 ,n5[12] ,n349);
    nand g696(n1178 ,n30[22] ,n54);
    nand g697(n1555 ,n831 ,n1166);
    nand g698(n1008 ,n13[8] ,n49);
    nand g699(n1290 ,n616 ,n406);
    nand g700(n918 ,n5[20] ,n43);
    nand g701(n1450 ,n190 ,n387);
    dff g702(.RN(n1), .SN(1'b1), .CK(n0), .D(n1499), .Q(n28[11]));
    nand g703(n1325 ,n769 ,n428);
    or g704(n465 ,n253 ,n356);
    nand g705(n1335 ,n813 ,n464);
    nor g706(n430 ,n97 ,n352);
    nand g707(n1341 ,n903 ,n375);
    nor g708(n1894 ,n1860 ,n24[8]);
    dff g709(.RN(n1), .SN(1'b1), .CK(n0), .D(n1302), .Q(n35[27]));
    nand g710(n1012 ,n15[5] ,n354);
    nand g711(n1768 ,n1262 ,n1703);
    nand g712(n1541 ,n468 ,n1199);
    nand g713(n1294 ,n621 ,n412);
    dff g714(.RN(n1), .SN(1'b1), .CK(n0), .D(n1653), .Q(n10[3]));
    nand g715(n668 ,n15[4] ,n354);
    dff g716(.RN(n1), .SN(1'b1), .CK(n0), .D(n1795), .Q(n31[9]));
    nand g717(n1420 ,n699 ,n1044);
    xnor g718(n326 ,n22[4] ,n32[4]);
    nand g719(n695 ,n32[11] ,n53);
    nand g720(n1388 ,n1284 ,n536);
    nand g721(n1499 ,n1133 ,n605);
    nand g722(n570 ,n22[6] ,n355);
    nor g723(n154 ,n60 ,n58);
    nand g724(n880 ,n35[1] ,n356);
    dff g725(.RN(n1), .SN(1'b1), .CK(n0), .D(n1639), .Q(n21[13]));
    nand g726(n622 ,n32[0] ,n350);
    dff g727(.RN(n1), .SN(1'b1), .CK(n0), .D(n1622), .Q(n30[9]));
    nand g728(n1298 ,n625 ,n489);
    nand g729(n1053 ,n26[8] ,n346);
    or g730(n442 ,n266 ,n356);
    nand g731(n875 ,n32[10] ,n53);
    nand g732(n1570 ,n840 ,n1179);
    dff g733(.RN(n1), .SN(1'b1), .CK(n0), .D(n1344), .Q(n13[30]));
    nand g734(n1723 ,n1271 ,n970);
    nand g735(n684 ,n33[21] ,n344);
    nand g736(n860 ,n32[16] ,n53);
    nand g737(n1674 ,n557 ,n927);
    nand g738(n803 ,n34[22] ,n352);
    dff g739(.RN(n1), .SN(1'b1), .CK(n0), .D(n1487), .Q(n26[18]));
    xnor g740(n323 ,n32[1] ,n28[1]);
    nand g741(n863 ,n32[15] ,n53);
    nor g742(n517 ,n87 ,n50);
    nand g743(n1258 ,n24[6] ,n51);
    nand g744(n814 ,n32[24] ,n53);
    nand g745(n652 ,n21[9] ,n51);
    dff g746(.RN(n1), .SN(1'b1), .CK(n0), .D(n1367), .Q(n29[6]));
    nand g747(n1926 ,n1913 ,n1910);
    nand g748(n744 ,n6[2] ,n349);
    nand g749(n1729 ,n169 ,n523);
    nand g750(n858 ,n4[20] ,n349);
    nand g751(n1534 ,n879 ,n1151);
    nand g752(n705 ,n11[11] ,n49);
    dff g753(.RN(n1), .SN(1'b1), .CK(n0), .D(n1711), .Q(n24[0]));
    dff g754(.RN(n1), .SN(1'b1), .CK(n0), .D(n1306), .Q(n35[18]));
    xor g755(n334 ,n7[1] ,n27[1]);
    or g756(n548 ,n341 ,n351);
    nor g757(n137 ,n21[0] ,n24[0]);
    not g758(n47 ,n53);
    nand g759(n1798 ,n734 ,n1288);
    nand g760(n1631 ,n202 ,n447);
    dff g761(.RN(n1), .SN(1'b1), .CK(n0), .D(n1760), .Q(n13[24]));
    nand g762(n1381 ,n1281 ,n449);
    dff g763(.RN(n1), .SN(1'b1), .CK(n0), .D(n1515), .Q(n34[10]));
    dff g764(.RN(n1), .SN(1'b1), .CK(n0), .D(n1707), .Q(n25[31]));
    nor g765(n458 ,n111 ,n353);
    nand g766(n662 ,n36[0] ,n355);
    nor g767(n540 ,n121 ,n344);
    nor g768(n528 ,n143 ,n352);
    nand g769(n1587 ,n750 ,n1144);
    nor g770(n1877 ,n24[11] ,n24[10]);
    nand g771(n703 ,n11[12] ,n49);
    nand g772(n1591 ,n160 ,n470);
    buf g773(n14[17], n11[17]);
    nand g774(n1914 ,n1874 ,n1873);
    nand g775(n977 ,n13[26] ,n344);
    dff g776(.RN(n1), .SN(1'b1), .CK(n0), .D(n1693), .Q(n24[11]));
    nand g777(n1046 ,n26[13] ,n45);
    nand g778(n895 ,n33[8] ,n49);
    nor g779(n545 ,n138 ,n351);
    nor g780(n403 ,n62 ,n350);
    dff g781(.RN(n1), .SN(1'b1), .CK(n0), .D(n1818), .Q(n32[19]));
    nor g782(n133 ,n29[4] ,n30[4]);
    nand g783(n941 ,n5[29] ,n349);
    nand g784(n1769 ,n1256 ,n1697);
    nand g785(n930 ,n9[2] ,n349);
    nand g786(n1161 ,n30[26] ,n54);
    nand g787(n1732 ,n224 ,n526);
    nand g788(n1152 ,n28[0] ,n46);
    nand g789(n1313 ,n815 ,n475);
    nand g790(n1594 ,n1194 ,n857);
    xnor g791(n36[2] ,n1933 ,n25[30]);
    nand g792(n1807 ,n756 ,n1491);
    nand g793(n1810 ,n617 ,n1471);
    nand g794(n1025 ,n26[28] ,n45);
    nand g795(n734 ,n31[10] ,n353);
    nand g796(n682 ,n33[20] ,n345);
    nand g797(n975 ,n13[28] ,n49);
    nand g798(n40 ,n27[2] ,n2);
    nand g799(n193 ,n26[26] ,n33[22]);
    dff g800(.RN(n1), .SN(1'b1), .CK(n0), .D(n1396), .Q(n12[28]));
    nand g801(n165 ,n26[14] ,n33[10]);
    nor g802(n505 ,n107 ,n351);
    nand g803(n568 ,n22[4] ,n55);
    nand g804(n1613 ,n1207 ,n704);
    nand g805(n1093 ,n32[15] ,n350);
    nand g806(n1793 ,n994 ,n1523);
    xnor g807(n319 ,n30[1] ,n23[1]);
    dff g808(.RN(n1), .SN(1'b1), .CK(n0), .D(n1772), .Q(n33[0]));
    or g809(n504 ,n312 ,n50);
    nand g810(n1626 ,n1218 ,n882);
    dff g811(.RN(n1), .SN(1'b1), .CK(n0), .D(n1629), .Q(n26[3]));
    dff g812(.RN(n1), .SN(1'b1), .CK(n0), .D(n1498), .Q(n28[12]));
    nand g813(n1784 ,n812 ,n1533);
    dff g814(.RN(n1), .SN(1'b1), .CK(n0), .D(n1358), .Q(n13[9]));
    nand g815(n752 ,n31[30] ,n353);
    dff g816(.RN(n1), .SN(1'b1), .CK(n0), .D(n1511), .Q(n28[4]));
    dff g817(.RN(n1), .SN(1'b1), .CK(n0), .D(n1360), .Q(n13[5]));
    nand g818(n1456 ,n183 ,n398);
    nand g819(n628 ,n36[1] ,n44);
    dff g820(.RN(n1), .SN(1'b1), .CK(n0), .D(n1786), .Q(n35[6]));
    dff g821(.RN(n1), .SN(1'b1), .CK(n0), .D(n1710), .Q(n24[1]));
    nand g822(n687 ,n15[1] ,n354);
    not g823(n1856 ,n21[26]);
    nand g824(n1590 ,n642 ,n768);
    dff g825(.RN(n1), .SN(1'b1), .CK(n0), .D(n1442), .Q(n26[28]));
    dff g826(.RN(n1), .SN(1'b1), .CK(n0), .D(n1404), .Q(n15[2]));
    nand g827(n1135 ,n28[10] ,n46);
    nand g828(n1200 ,n35[29] ,n44);
    dff g829(.RN(n1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n13[11]));
    nand g830(n862 ,n5[7] ,n349);
    nand g831(n1116 ,n28[22] ,n350);
    nand g832(n597 ,n21[19] ,n52);
    nor g833(n73 ,n21[19] ,n24[19]);
    nand g834(n1091 ,n32[16] ,n350);
    nand g835(n998 ,n13[13] ,n49);
    nand g836(n1775 ,n900 ,n1644);
    xnor g837(n250 ,n29[31] ,n30[31]);
    nand g838(n1376 ,n1090 ,n392);
    nand g839(n732 ,n4[19] ,n43);
    dff g840(.RN(n1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n13[20]));
    nand g841(n1508 ,n778 ,n1138);
    nand g842(n1457 ,n731 ,n1092);
    nand g843(n709 ,n33[25] ,n345);
    nand g844(n824 ,n29[16] ,n351);
    nor g845(n493 ,n74 ,n354);
    nand g846(n799 ,n35[13] ,n356);
    nand g847(n1127 ,n28[14] ,n350);
    dff g848(.RN(n1), .SN(1'b1), .CK(n0), .D(n1778), .Q(n30[6]));
    nor g849(n94 ,n26[28] ,n33[24]);
    nor g850(n463 ,n131 ,n42);
    nand g851(n712 ,n11[7] ,n345);
    nor g852(n483 ,n133 ,n352);
    nand g853(n1792 ,n999 ,n1524);
    nand g854(n1354 ,n995 ,n524);
    nand g855(n1421 ,n690 ,n563);
    nand g856(n1336 ,n883 ,n492);
    nand g857(n1215 ,n33[4] ,n55);
    nand g858(n1112 ,n28[25] ,n46);
    dff g859(.RN(n1), .SN(1'b1), .CK(n0), .D(n1503), .Q(n26[16]));
    xnor g860(n1850 ,n21[1] ,n22[1]);
    nand g861(n620 ,n32[2] ,n46);
    dff g862(.RN(n1), .SN(1'b1), .CK(n0), .D(n1576), .Q(n34[9]));
    dff g863(.RN(n1), .SN(1'b1), .CK(n0), .D(n1661), .Q(n24[29]));
    nand g864(n1577 ,n1183 ,n791);
    dff g865(.RN(n1), .SN(1'b1), .CK(n0), .D(n1353), .Q(n13[16]));
    nor g866(n479 ,n68 ,n49);
    nand g867(n926 ,n5[23] ,n43);
    nand g868(n1110 ,n28[27] ,n46);
    xnor g869(n256 ,n29[22] ,n30[22]);
    nand g870(n782 ,n26[12] ,n354);
    nand g871(n1593 ,n720 ,n1215);
    nand g872(n1182 ,n30[10] ,n54);
    nand g873(n690 ,n15[0] ,n354);
    nand g874(n762 ,n31[24] ,n352);
    or g875(n440 ,n246 ,n356);
    nand g876(n608 ,n21[8] ,n52);
    nand g877(n1368 ,n1068 ,n371);
    dff g878(.RN(n1), .SN(1'b1), .CK(n0), .D(n1480), .Q(n28[21]));
    nand g879(n1267 ,n24[0] ,n51);
    nand g880(n1699 ,n1257 ,n862);
    nand g881(n1488 ,n241 ,n420);
    nand g882(n845 ,n34[8] ,n353);
    or g883(n449 ,n321 ,n350);
    nand g884(n1205 ,n35[25] ,n45);
    nand g885(n1445 ,n174 ,n380);
    nand g886(n1433 ,n714 ,n1058);
    or g887(n435 ,n279 ,n356);
    nand g888(n1611 ,n701 ,n1206);
    nand g889(n1476 ,n1116 ,n594);
    buf g890(n14[21], n11[21]);
    nand g891(n1367 ,n1066 ,n370);
    nand g892(n1295 ,n623 ,n481);
    or g893(n419 ,n252 ,n353);
    nand g894(n219 ,n31[4] ,n34[4]);
    nand g895(n1305 ,n789 ,n414);
    xnor g896(n292 ,n26[20] ,n33[16]);
    nand g897(n784 ,n35[24] ,n356);
    nor g898(n93 ,n29[27] ,n30[27]);
    nand g899(n1728 ,n232 ,n519);
    dff g900(.RN(n1), .SN(1'b1), .CK(n0), .D(n1330), .Q(n31[14]));
    dff g901(.RN(n1), .SN(1'b1), .CK(n0), .D(n1430), .Q(n11[7]));
    nand g902(n864 ,n5[8] ,n43);
    nand g903(n1132 ,n28[12] ,n46);
    nand g904(n1440 ,n171 ,n372);
    nand g905(n1567 ,n838 ,n1198);
    dff g906(.RN(n1), .SN(1'b1), .CK(n0), .D(n1584), .Q(n34[5]));
    dff g907(.RN(n1), .SN(1'b1), .CK(n0), .D(n1296), .Q(n30[2]));
    buf g908(n16[1], n15[9]);
    dff g909(.RN(n1), .SN(1'b1), .CK(n0), .D(n1566), .Q(n34[14]));
    nand g910(n1206 ,n35[24] ,n45);
    nand g911(n1667 ,n1235 ,n922);
    buf g912(n17[6], 1'b0);
    nand g913(n743 ,n6[3] ,n43);
    nand g914(n813 ,n31[2] ,n352);
    dff g915(.RN(n1), .SN(1'b1), .CK(n0), .D(n1324), .Q(n31[21]));
    or g916(n404 ,n302 ,n46);
    dff g917(.RN(n1), .SN(1'b1), .CK(n0), .D(n1388), .Q(n29[17]));
    dff g918(.RN(n1), .SN(1'b1), .CK(n0), .D(n1486), .Q(n28[18]));
    or g919(n530 ,n242 ,n50);
    nand g920(n1484 ,n1119 ,n596);
    not g921(n1862 ,n21[29]);
    nand g922(n1238 ,n24[23] ,n348);
    nand g923(n1579 ,n845 ,n1184);
    xnor g924(n310 ,n30[2] ,n29[2]);
    nand g925(n1179 ,n30[12] ,n54);
    nand g926(n216 ,n31[6] ,n34[6]);
    not g927(n49 ,n45);
    nand g928(n1210 ,n30[11] ,n47);
    dff g929(.RN(n1), .SN(1'b1), .CK(n0), .D(n1459), .Q(n28[31]));
    nand g930(n1465 ,n189 ,n403);
    nand g931(n1493 ,n772 ,n1131);
    nor g932(n529 ,n134 ,n344);
    dff g933(.RN(n1), .SN(1'b1), .CK(n0), .D(n1336), .Q(n31[1]));
    nand g934(n1247 ,n24[15] ,n348);
    nand g935(n39 ,n27[1] ,n60);
    nand g936(n1282 ,n29[19] ,n48);
    nand g937(n636 ,n21[28] ,n51);
    nand g938(n1716 ,n968 ,n554);
    nand g939(n1117 ,n33[19] ,n355);
    nand g940(n994 ,n35[16] ,n356);
    nand g941(n842 ,n34[23] ,n352);
    nand g942(n903 ,n33[4] ,n345);
    nand g943(n1254 ,n24[9] ,n348);
    nand g944(n696 ,n11[17] ,n49);
    or g945(n455 ,n248 ,n352);
    nand g946(n935 ,n4[5] ,n43);
    dff g947(.RN(n1), .SN(1'b1), .CK(n0), .D(n1568), .Q(n34[13]));
    nand g948(n1134 ,n30[6] ,n54);
    buf g949(n12[19], n11[19]);
    not g950(n1854 ,n21[17]);
    dff g951(.RN(n1), .SN(1'b1), .CK(n0), .D(n1779), .Q(n30[7]));
    or g952(n375 ,n325 ,n345);
    nand g953(n196 ,n29[23] ,n30[23]);
    nand g954(n1321 ,n761 ,n423);
    nand g955(n1460 ,n185 ,n400);
    xnor g956(n303 ,n21[7] ,n24[7]);
    or g957(n453 ,n298 ,n356);
    or g958(n542 ,n268 ,n356);
    nand g959(n1698 ,n1255 ,n864);
    nand g960(n1218 ,n30[8] ,n47);
    nand g961(n1767 ,n2 ,n1709);
    dff g962(.RN(n1), .SN(1'b1), .CK(n0), .D(n1483), .Q(n23[0]));
    nand g963(n593 ,n21[23] ,n52);
    nand g964(n1007 ,n15[3] ,n354);
    nand g965(n1686 ,n1247 ,n885);
    dff g966(.RN(n1), .SN(1'b1), .CK(n0), .D(n1537), .Q(n34[31]));
    dff g967(.RN(n1), .SN(1'b1), .CK(n0), .D(n1695), .Q(n24[10]));
    nand g968(n1331 ,n787 ,n441);
    buf g969(n16[12], 1'b0);
    nand g970(n1096 ,n32[14] ,n46);
    nor g971(n110 ,n31[13] ,n34[13]);
    dff g972(.RN(n1), .SN(1'b1), .CK(n0), .D(n1688), .Q(n24[14]));
    nand g973(n900 ,n33[5] ,n345);
    nor g974(n74 ,n18[0] ,n33[0]);
    nor g975(n1902 ,n1869 ,n24[29]);
    dff g976(.RN(n1), .SN(1'b1), .CK(n0), .D(n1654), .Q(n10[2]));
    dff g977(.RN(n1), .SN(1'b1), .CK(n0), .D(n1317), .Q(n31[31]));
    dff g978(.RN(n1), .SN(1'b1), .CK(n0), .D(n1673), .Q(n24[22]));
    dff g979(.RN(n1), .SN(1'b1), .CK(n0), .D(n1563), .Q(n21[26]));
    nand g980(n1622 ,n1033 ,n674);
    nand g981(n1214 ,n35[19] ,n346);
    xnor g982(n278 ,n31[9] ,n34[9]);
    nand g983(n1033 ,n30[9] ,n48);
    dff g984(.RN(n1), .SN(1'b1), .CK(n0), .D(n1359), .Q(n13[7]));
    dff g985(.RN(n1), .SN(1'b1), .CK(n0), .D(n1845), .Q(n27[2]));
    nand g986(n1583 ,n774 ,n1134);
    nand g987(n1782 ,n869 ,n1536);
    nand g988(n1901 ,n21[23] ,n21[22]);
    nand g989(n1157 ,n30[30] ,n54);
    nand g990(n1580 ,n1186 ,n846);
    buf g991(n14[14], n11[14]);
    nand g992(n1542 ,n854 ,n1193);
    nand g993(n870 ,n32[13] ,n53);
    dff g994(.RN(n1), .SN(1'b1), .CK(n0), .D(n1606), .Q(n30[14]));
    nand g995(n1737 ,n231 ,n533);
    nand g996(n1018 ,n31[14] ,n41);
    nand g997(n1055 ,n29[8] ,n351);
    xnor g998(n291 ,n29[7] ,n30[7]);
    nor g999(n513 ,n94 ,n345);
    nand g1000(n713 ,n33[26] ,n345);
    nand g1001(n1278 ,n29[22] ,n351);
    nand g1002(n1359 ,n1010 ,n534);
    nand g1003(n879 ,n26[9] ,n354);
    nand g1004(n872 ,n4[1] ,n43);
    nand g1005(n816 ,n26[8] ,n354);
    nand g1006(n623 ,n30[3] ,n47);
    nand g1007(n1812 ,n1102 ,n1462);
    nand g1008(n1398 ,n677 ,n630);
    dff g1009(.RN(n1), .SN(1'b1), .CK(n0), .D(n1583), .Q(n34[6]));
    nand g1010(n1411 ,n223 ,n545);
    nand g1011(n748 ,n6[0] ,n43);
    nand g1012(n797 ,n33[9] ,n345);
    dff g1013(.RN(n1), .SN(1'b1), .CK(n0), .D(n1651), .Q(n21[9]));
    nand g1014(n962 ,n10[3] ,n356);
    nand g1015(n163 ,n7[1] ,n59);
    dff g1016(.RN(n1), .SN(1'b1), .CK(n0), .D(n1295), .Q(n30[3]));
    xor g1017(n361 ,n21[1] ,n23[1]);
    nand g1018(n1190 ,n30[4] ,n54);
    nand g1019(n658 ,n21[17] ,n348);
    dff g1020(.RN(n1), .SN(1'b1), .CK(n0), .D(n1434), .Q(n11[4]));
    nand g1021(n757 ,n26[17] ,n354);
    dff g1022(.RN(n1), .SN(1'b1), .CK(n0), .D(n1702), .Q(n28[5]));
    nand g1023(n1642 ,n649 ,n894);
    nand g1024(n208 ,n28[30] ,n32[30]);
    nand g1025(n973 ,n13[30] ,n345);
    nand g1026(n572 ,n27[0] ,n359);
    nor g1027(n72 ,n28[0] ,n32[0]);
    nor g1028(n80 ,n21[13] ,n24[13]);
    or g1029(n1846 ,n1837 ,n1842);
    nand g1030(n1733 ,n165 ,n415);
    dff g1031(.RN(n1), .SN(1'b1), .CK(n0), .D(n1573), .Q(n21[25]));
    or g1032(n1920 ,n1911 ,n1906);
    dff g1033(.RN(n1), .SN(1'b1), .CK(n0), .D(n1723), .Q(n25[29]));
    nand g1034(n925 ,n9[4] ,n349);
    nand g1035(n1467 ,n737 ,n1101);
    nand g1036(n1621 ,n669 ,n1216);
    dff g1037(.RN(n1), .SN(1'b1), .CK(n0), .D(n1784), .Q(n35[4]));
    dff g1038(.RN(n1), .SN(1'b1), .CK(n0), .D(n1481), .Q(n26[19]));
    dff g1039(.RN(n1), .SN(1'b1), .CK(n0), .D(n1750), .Q(n13[4]));
    nand g1040(n1084 ,n29[2] ,n47);
    nand g1041(n723 ,n4[18] ,n349);
    nand g1042(n969 ,n14[1] ,n50);
    nor g1043(n502 ,n112 ,n351);
    xnor g1044(n340 ,n32[7] ,n28[7]);
    or g1045(n1872 ,n20[1] ,n20[0]);
    nand g1046(n993 ,n13[16] ,n49);
    xnor g1047(n284 ,n26[11] ,n33[7]);
    xnor g1048(n246 ,n31[25] ,n34[25]);
    nand g1049(n555 ,n22[1] ,n45);
    dff g1050(.RN(n1), .SN(1'b1), .CK(n0), .D(n1414), .Q(n26[31]));
    nor g1051(n78 ,n21[15] ,n24[15]);
    dff g1052(.RN(n1), .SN(1'b1), .CK(n0), .D(n1410), .Q(n11[21]));
    nand g1053(n1230 ,n35[12] ,n346);
    nand g1054(n1306 ,n794 ,n542);
    nand g1055(n1102 ,n32[11] ,n46);
    nand g1056(n1884 ,n24[16] ,n1870);
    nand g1057(n905 ,n33[3] ,n344);
    nand g1058(n1256 ,n29[30] ,n351);
    nor g1059(n65 ,n26[29] ,n33[25]);
    xnor g1060(n301 ,n21[10] ,n24[10]);
    not g1061(n1860 ,n24[9]);
    dff g1062(.RN(n1), .SN(1'b1), .CK(n0), .D(n1574), .Q(n21[24]));
    nand g1063(n694 ,n11[18] ,n344);
    nand g1064(n1310 ,n928 ,n491);
    nand g1065(n1569 ,n1176 ,n814);
    nand g1066(n671 ,n12[31] ,n345);
    nor g1067(n66 ,n22[6] ,n35[6]);
    nand g1068(n1346 ,n976 ,n508);
    xnor g1069(n1851 ,n21[0] ,n22[0]);
    dff g1070(.RN(n1), .SN(1'b1), .CK(n0), .D(n1788), .Q(n31[5]));
    nand g1071(n585 ,n21[31] ,n52);
    nand g1072(n1638 ,n797 ,n1226);
    or g1073(n509 ,n283 ,n47);
    nand g1074(n574 ,n18[0] ,n358);
    nand g1075(n896 ,n35[3] ,n42);
    dff g1076(.RN(n1), .SN(1'b1), .CK(n0), .D(n1521), .Q(n26[11]));
    nand g1077(n995 ,n13[15] ,n344);
    dff g1078(.RN(n1), .SN(1'b1), .CK(n0), .D(n1810), .Q(n32[5]));
    nand g1079(n1721 ,n204 ,n505);
    or g1080(n436 ,n276 ,n353);
    nor g1081(n1879 ,n1867 ,n24[15]);
    not g1082(n1866 ,n24[12]);
    xnor g1083(n268 ,n31[18] ,n34[18]);
    nand g1084(n1372 ,n1080 ,n384);
    or g1085(n416 ,n250 ,n352);
    nand g1086(n1692 ,n580 ,n872);
    xnor g1087(n19[1] ,n1850 ,n18[1]);
    nand g1088(n170 ,n28[5] ,n32[5]);
    nand g1089(n715 ,n11[4] ,n50);
    nand g1090(n1754 ,n1004 ,n1733);
    nand g1091(n617 ,n32[5] ,n350);
    nand g1092(n787 ,n31[11] ,n352);
    nand g1093(n1418 ,n217 ,n497);
    nand g1094(n1358 ,n1006 ,n532);
    nand g1095(n1000 ,n13[12] ,n49);
    dff g1096(.RN(n1), .SN(1'b1), .CK(n0), .D(n1492), .Q(n28[16]));
    xnor g1097(n248 ,n29[6] ,n30[6]);
    dff g1098(.RN(n1), .SN(1'b1), .CK(n0), .D(n1320), .Q(n31[26]));
    nand g1099(n1068 ,n32[30] ,n350);
    nand g1100(n1332 ,n796 ,n451);
    dff g1101(.RN(n1), .SN(1'b1), .CK(n0), .D(n1595), .Q(n21[21]));
    xnor g1102(n244 ,n26[9] ,n33[5]);
    nand g1103(n917 ,n31[3] ,n352);
    nor g1104(n111 ,n29[5] ,n30[5]);
    nand g1105(n645 ,n21[18] ,n347);
    nor g1106(n125 ,n22[7] ,n32[7]);
    nand g1107(n1304 ,n788 ,n442);
    buf g1108(n17[7], 1'b0);
    dff g1109(.RN(n1), .SN(1'b1), .CK(n0), .D(n1579), .Q(n34[8]));
    nand g1110(n670 ,n13[0] ,n345);
    or g1111(n490 ,n17[0] ,n357);
    dff g1112(.RN(n1), .SN(1'b1), .CK(n0), .D(n1762), .Q(n13[28]));
    nand g1113(n166 ,n28[13] ,n32[13]);
    or g1114(n524 ,n293 ,n50);
    nand g1115(n1551 ,n636 ,n852);
    dff g1116(.RN(n1), .SN(1'b1), .CK(n0), .D(n1787), .Q(n31[4]));
    nand g1117(n558 ,n22[2] ,n51);
    or g1118(n369 ,n340 ,n48);
    nor g1119(n372 ,n106 ,n46);
    nand g1120(n1378 ,n1104 ,n402);
    dff g1121(.RN(n1), .SN(1'b1), .CK(n0), .D(n1735), .Q(n15[9]));
    dff g1122(.RN(n1), .SN(1'b1), .CK(n0), .D(n1802), .Q(n31[13]));
    nand g1123(n916 ,n11[13] ,n50);
    nand g1124(n1087 ,n32[19] ,n350);
    nand g1125(n1417 ,n696 ,n1040);
    nand g1126(n1337 ,n738 ,n471);
    nand g1127(n1414 ,n702 ,n1041);
    nand g1128(n203 ,n29[10] ,n30[10]);
    nand g1129(n1436 ,n717 ,n1061);
    dff g1130(.RN(n1), .SN(1'b1), .CK(n0), .D(n1758), .Q(n13[21]));
    dff g1131(.RN(n1), .SN(1'b1), .CK(n0), .D(n1378), .Q(n32[10]));
    nand g1132(n802 ,n35[12] ,n356);
    or g1133(n482 ,n330 ,n344);
    dff g1134(.RN(n1), .SN(1'b1), .CK(n0), .D(n1744), .Q(n15[6]));
    nand g1135(n1383 ,n1274 ,n509);
    dff g1136(.RN(n1), .SN(1'b1), .CK(n0), .D(n1624), .Q(n33[17]));
    nand g1137(n1270 ,n25[30] ,n348);
    nand g1138(n1588 ,n159 ,n418);
    dff g1139(.RN(n1), .SN(1'b1), .CK(n0), .D(n1682), .Q(n22[1]));
    nand g1140(n933 ,n5[19] ,n349);
    or g1141(n487 ,n17[2] ,n357);
    nand g1142(n226 ,n31[28] ,n34[28]);
    xnor g1143(n264 ,n31[30] ,n34[30]);
    nand g1144(n552 ,n22[0] ,n45);
    dff g1145(.RN(n1), .SN(1'b1), .CK(n0), .D(n1351), .Q(n13[18]));
    nor g1146(n1918 ,n1901 ,n1900);
    nand g1147(n1581 ,n848 ,n1185);
    buf g1148(n12[25], n11[25]);
    nand g1149(n1426 ,n707 ,n1050);
    nand g1150(n1783 ,n880 ,n1535);
    dff g1151(.RN(n1), .SN(1'b1), .CK(n0), .D(n488), .Q(n17[1]));
    nand g1152(n1387 ,n1282 ,n366);
    nand g1153(n69 ,n60 ,n58);
    xnor g1154(n254 ,n29[26] ,n30[26]);
    dff g1155(.RN(n1), .SN(1'b1), .CK(n0), .D(n1756), .Q(n29[20]));
    nand g1156(n1750 ,n1015 ,n1741);
    dff g1157(.RN(n1), .SN(1'b1), .CK(n0), .D(n1612), .Q(n33[23]));
    nand g1158(n1111 ,n28[26] ,n350);
    nand g1159(n907 ,n33[2] ,n49);
    nand g1160(n557 ,n22[3] ,n348);
    nand g1161(n972 ,n13[31] ,n50);
    nand g1162(n821 ,n4[26] ,n43);
    xor g1163(n19[3] ,n21[3] ,n22[3]);
    nand g1164(n1655 ,n912 ,n664);
    not g1165(n41 ,n54);
    dff g1166(.RN(n1), .SN(1'b1), .CK(n0), .D(n1409), .Q(n11[22]));
    xnor g1167(n19[0] ,n1851 ,n18[0]);
    nor g1168(n1878 ,n1866 ,n24[13]);
    dff g1169(.RN(n1), .SN(1'b1), .CK(n0), .D(n1806), .Q(n31[23]));
    dff g1170(.RN(n1), .SN(1'b1), .CK(n0), .D(n1565), .Q(n30[25]));
    nand g1171(n809 ,n35[6] ,n356);
    dff g1172(.RN(n1), .SN(1'b1), .CK(n0), .D(n1315), .Q(n35[10]));
    nand g1173(n1207 ,n30[12] ,n48);
    nand g1174(n664 ,n36[1] ,n56);
    or g1175(n377 ,n258 ,n356);
    nand g1176(n1649 ,n214 ,n484);
    nand g1177(n1385 ,n1277 ,n516);
    dff g1178(.RN(n1), .SN(1'b1), .CK(n0), .D(n1364), .Q(n29[9]));
    nand g1179(n1600 ,n733 ,n1197);
    nand g1180(n672 ,n12[30] ,n50);
    nand g1181(n1529 ,n801 ,n1149);
    nor g1182(n415 ,n140 ,n344);
    nand g1183(n1257 ,n24[7] ,n51);
    dff g1184(.RN(n1), .SN(1'b1), .CK(n0), .D(n1793), .Q(n35[16]));
    nand g1185(n162 ,n7[0] ,n59);
    nand g1186(n963 ,n8[1] ,n43);
    or g1187(n492 ,n307 ,n353);
    xnor g1188(n36[1] ,n1933 ,n25[29]);
    nand g1189(n1416 ,n694 ,n1039);
    nand g1190(n1724 ,n194 ,n511);
    nand g1191(n1262 ,n29[29] ,n351);
    buf g1192(n16[15], 1'b0);
    buf g1193(n16[11], n15[7]);
    buf g1194(n14[11], n11[11]);
    nand g1195(n982 ,n13[23] ,n345);
    nand g1196(n1168 ,n30[18] ,n54);
    nor g1197(n409 ,n71 ,n356);
    nand g1198(n1648 ,n893 ,n1273);
    dff g1199(.RN(n1), .SN(1'b1), .CK(n0), .D(n1547), .Q(n26[8]));
    xnor g1200(n331 ,n22[1] ,n32[1]);
    or g1201(n356 ,n40 ,n69);
    nor g1202(n135 ,n28[10] ,n32[10]);
    nand g1203(n1138 ,n33[13] ,n55);
    nand g1204(n554 ,n22[2] ,n45);
    nand g1205(n1478 ,n575 ,n743);
    nand g1206(n1458 ,n184 ,n399);
    buf g1207(n14[4], n11[28]);
    nor g1208(n134 ,n22[0] ,n35[0]);
    dff g1209(.RN(n1), .SN(1'b1), .CK(n0), .D(n1812), .Q(n32[11]));
    dff g1210(.RN(n1), .SN(1'b1), .CK(n0), .D(n1831), .Q(n29[13]));
    or g1211(n429 ,n324 ,n354);
    nand g1212(n1751 ,n1011 ,n1738);
    nand g1213(n51 ,n148 ,n99);
    dff g1214(.RN(n1), .SN(1'b1), .CK(n0), .D(n1403), .Q(n11[27]));
    nand g1215(n1607 ,n713 ,n1203);
    nand g1216(n1054 ,n26[7] ,n45);
    dff g1217(.RN(n1), .SN(1'b1), .CK(n0), .D(n1627), .Q(n33[15]));
    nand g1218(n912 ,n10[1] ,n42);
    nand g1219(n1834 ,n7[0] ,n1517);
    dff g1220(.RN(n1), .SN(1'b1), .CK(n0), .D(n1436), .Q(n11[2]));
    nand g1221(n805 ,n35[9] ,n356);
    nand g1222(n1708 ,n1264 ,n958);
    nand g1223(n1364 ,n1049 ,n476);
    nor g1224(n85 ,n21[22] ,n24[22]);
    nand g1225(n1370 ,n1078 ,n381);
    nand g1226(n1243 ,n24[19] ,n348);
    nand g1227(n892 ,n33[10] ,n49);
    nand g1228(n562 ,n22[1] ,n355);
    buf g1229(n16[4], n15[0]);
    nand g1230(n1599 ,n867 ,n1158);
    nand g1231(n1787 ,n807 ,n1530);
    nand g1232(n1921 ,n1905 ,n1917);
    nand g1233(n1605 ,n721 ,n1202);
    xnor g1234(n337 ,n21[30] ,n24[30]);
    nand g1235(n1771 ,n953 ,n1662);
    dff g1236(.RN(n1), .SN(1'b1), .CK(n0), .D(n1347), .Q(n13[26]));
    dff g1237(.RN(n1), .SN(1'b1), .CK(n0), .D(n1775), .Q(n33[5]));
    nand g1238(n1755 ,n1000 ,n1732);
    nand g1239(n1602 ,n865 ,n1200);
    nand g1240(n1900 ,n21[21] ,n21[20]);
    dff g1241(.RN(n1), .SN(1'b1), .CK(n0), .D(n1805), .Q(n31[19]));
    nand g1242(n1443 ,n172 ,n376);
    or g1243(n485 ,n332 ,n48);
    nand g1244(n1092 ,n33[24] ,n355);
    nand g1245(n1788 ,n804 ,n1528);
    xnor g1246(n279 ,n31[31] ,n34[31]);
    dff g1247(.RN(n1), .SN(1'b1), .CK(n0), .D(n1613), .Q(n30[12]));
    nor g1248(n500 ,n125 ,n351);
    dff g1249(.RN(n1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n29[12]));
    nand g1250(n1297 ,n626 ,n469);
    or g1251(n390 ,n323 ,n351);
    nor g1252(n1915 ,n1887 ,n1885);
    nand g1253(n1226 ,n35[9] ,n45);
    nand g1254(n661 ,n36[1] ,n355);
    or g1255(n518 ,n288 ,n50);
    nand g1256(n1816 ,n1095 ,n1454);
    buf g1257(n12[1], n11[29]);
    nand g1258(n1061 ,n26[2] ,n346);
    nor g1259(n143 ,n29[13] ,n30[13]);
    nand g1260(n1563 ,n639 ,n821);
    dff g1261(.RN(n1), .SN(1'b1), .CK(n0), .D(n1781), .Q(n34[3]));
    nand g1262(n625 ,n30[1] ,n351);
    nand g1263(n191 ,n31[26] ,n34[26]);
    dff g1264(.RN(n1), .SN(1'b1), .CK(n0), .D(n1314), .Q(n35[0]));
    xnor g1265(n314 ,n21[6] ,n24[6]);
    buf g1266(n14[26], n11[26]);
    or g1267(n508 ,n265 ,n50);
    dff g1268(.RN(n1), .SN(1'b1), .CK(n0), .D(n1656), .Q(n10[0]));
    nand g1269(n1548 ,n826 ,n1141);
    nand g1270(n1615 ,n874 ,n1209);
    dff g1271(.RN(n1), .SN(1'b1), .CK(n0), .D(n1338), .Q(n34[0]));
    nand g1272(n1553 ,n836 ,n1165);
    nand g1273(n808 ,n35[7] ,n42);
    nand g1274(n1756 ,n1280 ,n1729);
    nor g1275(n457 ,n146 ,n356);
    nand g1276(n221 ,n31[12] ,n34[12]);
    nand g1277(n807 ,n31[4] ,n352);
    nand g1278(n1362 ,n1020 ,n548);
    dff g1279(.RN(n1), .SN(1'b1), .CK(n0), .D(n1408), .Q(n11[23]));
    nand g1280(n819 ,n4[31] ,n43);
    nand g1281(n1657 ,n654 ,n913);
    dff g1282(.RN(n1), .SN(1'b1), .CK(n0), .D(n1803), .Q(n35[28]));
    nand g1283(n1389 ,n1012 ,n571);
    buf g1284(n12[10], n11[10]);
    nand g1285(n1076 ,n32[26] ,n46);
    nand g1286(n881 ,n26[3] ,n354);
    nand g1287(n1289 ,n615 ,n405);
    nand g1288(n1481 ,n745 ,n1117);
    xnor g1289(n338 ,n21[31] ,n24[31]);
    nor g1290(n84 ,n21[5] ,n24[5]);
    nand g1291(n1402 ,n680 ,n629);
    not g1292(n1855 ,n21[19]);
    nand g1293(n37 ,n2 ,n61);
    buf g1294(n17[3], 1'b0);
    nand g1295(n1080 ,n32[23] ,n350);
    nand g1296(n1014 ,n13[5] ,n49);
    dff g1297(.RN(n1), .SN(1'b1), .CK(n0), .D(n1478), .Q(n23[3]));
    nand g1298(n948 ,n5[10] ,n349);
    xnor g1299(n251 ,n29[30] ,n30[30]);
    nand g1300(n1260 ,n24[4] ,n51);
    nor g1301(n519 ,n75 ,n47);
    or g1302(n397 ,n249 ,n50);
    nand g1303(n1013 ,n15[6] ,n354);
    nand g1304(n1539 ,n873 ,n1157);
    nand g1305(n882 ,n32[8] ,n53);
    nor g1306(n79 ,n21[14] ,n24[14]);
    xor g1307(n19[2] ,n21[2] ,n22[2]);
    nand g1308(n38 ,n27[0] ,n58);
    nand g1309(n1739 ,n1005 ,n662);
    nand g1310(n774 ,n34[6] ,n41);
    nand g1311(n833 ,n4[27] ,n43);
    nand g1312(n1532 ,n222 ,n462);
    nand g1313(n1379 ,n1109 ,n404);
    nand g1314(n635 ,n21[23] ,n348);
    nand g1315(n919 ,n5[24] ,n349);
    nand g1316(n1274 ,n29[25] ,n351);
    nand g1317(n835 ,n34[18] ,n353);
    nor g1318(n515 ,n89 ,n345);
    nand g1319(n1494 ,n1126 ,n601);
    dff g1320(.RN(n1), .SN(1'b1), .CK(n0), .D(n1592), .Q(n30[18]));
    nand g1321(n1779 ,n1221 ,n1632);
    dff g1322(.RN(n1), .SN(1'b1), .CK(n0), .D(n1714), .Q(n18[0]));
    nand g1323(n736 ,n26[23] ,n354);
    nor g1324(n388 ,n77 ,n350);
    nand g1325(n1543 ,n1160 ,n740);
    dff g1326(.RN(n1), .SN(1'b1), .CK(n0), .D(n1585), .Q(n30[20]));
    dff g1327(.RN(n1), .SN(1'b1), .CK(n0), .D(n1391), .Q(n12[31]));
    nand g1328(n1232 ,n24[30] ,n51);
    nand g1329(n1757 ,n1278 ,n1728);
    nand g1330(n1352 ,n991 ,n374);
    nand g1331(n943 ,n5[14] ,n43);
    nand g1332(n1334 ,n917 ,n495);
    nand g1333(n846 ,n32[21] ,n53);
    nand g1334(n1066 ,n29[6] ,n48);
    nor g1335(n393 ,n72 ,n48);
    dff g1336(.RN(n1), .SN(1'b1), .CK(n0), .D(n1291), .Q(n32[4]));
    nand g1337(n698 ,n11[16] ,n50);
    nand g1338(n890 ,n33[11] ,n50);
    dff g1339(.RN(n1), .SN(1'b1), .CK(n0), .D(n1383), .Q(n29[25]));
    dff g1340(.RN(n1), .SN(1'b1), .CK(n0), .D(n1406), .Q(n11[25]));
    nand g1341(n1736 ,n1265 ,n984);
    nand g1342(n1703 ,n220 ,n498);
    dff g1343(.RN(n1), .SN(1'b1), .CK(n0), .D(n1467), .Q(n26[22]));
    buf g1344(n12[3], n11[31]);
    nand g1345(n1145 ,n28[5] ,n350);
    nand g1346(n960 ,n5[1] ,n349);
    nor g1347(n447 ,n103 ,n42);
    nand g1348(n885 ,n5[15] ,n349);
    nand g1349(n174 ,n21[26] ,n24[26]);
    nand g1350(n631 ,n21[31] ,n51);
    xor g1351(n19[7] ,n21[7] ,n22[7]);
    nand g1352(n583 ,n21[0] ,n347);
    nand g1353(n171 ,n21[29] ,n24[29]);
    nand g1354(n767 ,n31[21] ,n352);
    buf g1355(n16[7], n15[3]);
    nand g1356(n721 ,n33[27] ,n49);
    nand g1357(n1547 ,n816 ,n1156);
    nand g1358(n192 ,n21[0] ,n24[0]);
    nand g1359(n959 ,n31[13] ,n41);
    nand g1360(n653 ,n21[8] ,n51);
    dff g1361(.RN(n1), .SN(1'b1), .CK(n0), .D(n1706), .Q(n24[3]));
    nand g1362(n1645 ,n650 ,n898);
    nand g1363(n179 ,n29[9] ,n30[9]);
    xnor g1364(n257 ,n29[21] ,n30[21]);
    nor g1365(n407 ,n84 ,n46);
    nand g1366(n1229 ,n30[4] ,n48);
    nand g1367(n1017 ,n13[3] ,n50);
    dff g1368(.RN(n1), .SN(1'b1), .CK(n0), .D(n1586), .Q(n34[4]));
    nand g1369(n1459 ,n1097 ,n585);
    nand g1370(n188 ,n22[5] ,n35[5]);
    nand g1371(n996 ,n15[10] ,n354);
    dff g1372(.RN(n1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n13[2]));
    nand g1373(n837 ,n32[25] ,n53);
    nand g1374(n1083 ,n32[21] ,n46);
    nand g1375(n575 ,n23[3] ,n347);
    nand g1376(n629 ,n36[0] ,n45);
    dff g1377(.RN(n1), .SN(1'b1), .CK(n0), .D(n1600), .Q(n33[30]));
    nand g1378(n710 ,n11[8] ,n344);
    nand g1379(n1651 ,n652 ,n906);
    nand g1380(n725 ,n26[28] ,n354);
    nand g1381(n699 ,n11[15] ,n49);
    nand g1382(n1216 ,n35[18] ,n45);
    nand g1383(n921 ,n9[5] ,n43);
    nand g1384(n584 ,n18[1] ,n347);
    dff g1385(.RN(n1), .SN(1'b1), .CK(n0), .D(n1657), .Q(n21[7]));
    nor g1386(n89 ,n26[26] ,n33[22]);
    nand g1387(n1839 ,n2 ,n1764);
    nand g1388(n1109 ,n32[8] ,n350);
    xnor g1389(n1852 ,n23[0] ,n24[0]);
    nand g1390(n1139 ,n28[8] ,n46);
    buf g1391(n12[23], n11[23]);
    nand g1392(n1089 ,n29[1] ,n48);
    nand g1393(n817 ,n4[25] ,n43);
    nand g1394(n1635 ,n890 ,n1223);
    nand g1395(n1500 ,n199 ,n430);
    not g1396(n1858 ,n24[4]);
    nand g1397(n1823 ,n1076 ,n1445);
    nand g1398(n1373 ,n1081 ,n383);
    nand g1399(n718 ,n11[1] ,n49);
    nand g1400(n1043 ,n29[10] ,n47);
    nand g1401(n818 ,n34[16] ,n352);
    dff g1402(.RN(n1), .SN(1'b1), .CK(n0), .D(n1783), .Q(n35[1]));
    nand g1403(n1312 ,n896 ,n465);
    dff g1404(.RN(n1), .SN(1'b1), .CK(n0), .D(n1840), .Q(n28[0]));
    nand g1405(n865 ,n33[29] ,n345);
    nand g1406(n1520 ,n195 ,n362);
    dff g1407(.RN(n1), .SN(1'b1), .CK(n0), .D(n1684), .Q(n24[16]));
    dff g1408(.RN(n1), .SN(1'b1), .CK(n0), .D(n1619), .Q(n30[10]));
    nand g1409(n1062 ,n29[7] ,n351);
    nand g1410(n1345 ,n974 ,n452);
    nand g1411(n1603 ,n724 ,n1201);
    xnor g1412(n339 ,n32[6] ,n28[6]);
    nand g1413(n1887 ,n21[13] ,n21[12]);
    nor g1414(n1748 ,n27[1] ,n1518);
    nor g1415(n122 ,n29[8] ,n30[8]);
    nor g1416(n145 ,n26[10] ,n33[6]);
    nand g1417(n1647 ,n213 ,n540);
    dff g1418(.RN(n1), .SN(1'b1), .CK(n0), .D(n1333), .Q(n31[6]));
    xnor g1419(n272 ,n31[7] ,n34[7]);
    nand g1420(n1423 ,n916 ,n1046);
    nand g1421(n675 ,n12[28] ,n345);
    nand g1422(n1744 ,n1013 ,n570);
    xnor g1423(n288 ,n26[24] ,n33[20]);
    dff g1424(.RN(n1), .SN(1'b1), .CK(n0), .D(n1299), .Q(n35[31]));
    dff g1425(.RN(n1), .SN(1'b1), .CK(n0), .D(n1413), .Q(n11[20]));
    nand g1426(n720 ,n26[4] ,n354);
    nand g1427(n783 ,n31[12] ,n352);
    nand g1428(n949 ,n5[9] ,n43);
    nand g1429(n1601 ,n1136 ,n863);
    dff g1430(.RN(n1), .SN(1'b1), .CK(n0), .D(n1327), .Q(n31[17]));
    nand g1431(n1485 ,n1121 ,n597);
    nand g1432(n1393 ,n672 ,n1022);
    nand g1433(n1660 ,n567 ,n915);
    nand g1434(n1432 ,n868 ,n1056);
    nor g1435(n396 ,n78 ,n350);
    or g1436(n481 ,n329 ,n48);
    nand g1437(n1709 ,n7[2] ,n823);
    nand g1438(n827 ,n32[26] ,n53);
    nand g1439(n234 ,n21[5] ,n24[5]);
    nand g1440(n904 ,n33[12] ,n49);
    not g1441(n43 ,n51);
    nor g1442(n1928 ,n1922 ,n1924);
    nand g1443(n1431 ,n706 ,n1052);
    nand g1444(n1107 ,n28[28] ,n46);
    dff g1445(.RN(n1), .SN(1'b1), .CK(n0), .D(n1578), .Q(n26[6]));
    nand g1446(n1029 ,n26[25] ,n44);
    dff g1447(.RN(n1), .SN(1'b1), .CK(n0), .D(n1625), .Q(n33[16]));
    nand g1448(n1530 ,n212 ,n483);
    dff g1449(.RN(n1), .SN(1'b1), .CK(n0), .D(n1420), .Q(n11[15]));
    nand g1450(n1395 ,n668 ,n568);
    buf g1451(n12[16], n11[16]);
    dff g1452(.RN(n1), .SN(1'b1), .CK(n0), .D(n1342), .Q(n33[3]));
    nand g1453(n746 ,n6[1] ,n43);
    xnor g1454(n295 ,n28[19] ,n32[19]);
    nand g1455(n215 ,n22[0] ,n35[0]);
    nand g1456(n1051 ,n26[9] ,n45);
    nand g1457(n567 ,n22[7] ,n348);
    nand g1458(n691 ,n11[21] ,n49);
    nand g1459(n1404 ,n678 ,n561);
    nand g1460(n1363 ,n1030 ,n544);
    dff g1461(.RN(n1), .SN(1'b1), .CK(n0), .D(n1830), .Q(n29[11]));
    nand g1462(n159 ,n30[3] ,n23[3]);
    dff g1463(.RN(n1), .SN(1'b1), .CK(n0), .D(n1590), .Q(n21[22]));
    nand g1464(n1009 ,n15[7] ,n354);
    nand g1465(n168 ,n28[8] ,n32[8]);
    dff g1466(.RN(n1), .SN(1'b1), .CK(n0), .D(n1558), .Q(n34[18]));
    xnor g1467(n297 ,n31[17] ,n34[17]);
    nor g1468(n418 ,n139 ,n352);
    nor g1469(n141 ,n26[12] ,n33[8]);
    nand g1470(n686 ,n11[24] ,n344);
    dff g1471(.RN(n1), .SN(1'b1), .CK(n0), .D(n1431), .Q(n26[30]));
    nand g1472(n1785 ,n811 ,n1532);
    nand g1473(n648 ,n21[13] ,n51);
    nand g1474(n968 ,n14[2] ,n50);
    nor g1475(n121 ,n22[2] ,n35[2]);
    nand g1476(n1726 ,n193 ,n515);
    or g1477(n499 ,n275 ,n42);
    nand g1478(n908 ,n4[3] ,n43);
    xnor g1479(n315 ,n30[0] ,n23[0]);
    nand g1480(n212 ,n29[4] ,n30[4]);
    or g1481(n371 ,n337 ,n350);
    buf g1482(n14[31], n12[31]);
    nand g1483(n1350 ,n989 ,n397);
    dff g1484(.RN(n1), .SN(1'b1), .CK(n0), .D(n1821), .Q(n32[21]));
    dff g1485(.RN(n1), .SN(1'b1), .CK(n0), .D(n1316), .Q(n26[1]));
    nand g1486(n1419 ,n698 ,n1042);
    dff g1487(.RN(n1), .SN(1'b1), .CK(n0), .D(n1599), .Q(n34[29]));
    nand g1488(n958 ,n5[2] ,n43);
    nand g1489(n855 ,n4[29] ,n349);
    nor g1490(n76 ,n28[2] ,n32[2]);
    nand g1491(n1120 ,n33[18] ,n55);
    nand g1492(n1099 ,n32[12] ,n350);
    nand g1493(n891 ,n5[16] ,n349);
    nand g1494(n707 ,n11[10] ,n50);
    nor g1495(n362 ,n67 ,n356);
    dff g1496(.RN(n1), .SN(1'b1), .CK(n0), .D(n1502), .Q(n28[9]));
    nand g1497(n1303 ,n785 ,n440);
    dff g1498(.RN(n1), .SN(1'b1), .CK(n0), .D(n1374), .Q(n32[18]));
    or g1499(n366 ,n295 ,n351);
    dff g1500(.RN(n1), .SN(1'b1), .CK(n0), .D(n1634), .Q(n33[12]));
    nand g1501(n1349 ,n988 ,n518);
    dff g1502(.RN(n1), .SN(1'b1), .CK(n0), .D(n1379), .Q(n32[8]));
    nor g1503(n116 ,n29[12] ,n30[12]);
    nand g1504(n945 ,n5[30] ,n43);
    or g1505(n471 ,n319 ,n41);
    nand g1506(n730 ,n26[25] ,n354);
    dff g1507(.RN(n1), .SN(1'b1), .CK(n0), .D(n1761), .Q(n13[25]));
    nand g1508(n828 ,n34[15] ,n353);
    nor g1509(n1908 ,n1892 ,n1891);
    dff g1510(.RN(n1), .SN(1'b1), .CK(n0), .D(n1765), .Q(n29[27]));
    nor g1511(n100 ,n33[28] ,n36[0]);
    nor g1512(n364 ,n98 ,n351);
    nand g1513(n1119 ,n28[20] ,n46);
    xnor g1514(n299 ,n21[17] ,n24[17]);
    nand g1515(n1738 ,n238 ,n537);
    xnor g1516(n36[0] ,n1933 ,n25[28]);
    nand g1517(n1564 ,n828 ,n1154);
    nand g1518(n796 ,n31[7] ,n352);
    nand g1519(n1627 ,n980 ,n1275);
    nand g1520(n198 ,n22[6] ,n35[6]);
    nand g1521(n1797 ,n726 ,n1631);
    nand g1522(n1561 ,n640 ,n833);
    dff g1523(.RN(n1), .SN(1'b1), .CK(n0), .D(n1546), .Q(n21[29]));
    dff g1524(.RN(n1), .SN(1'b1), .CK(n0), .D(n1545), .Q(n30[30]));
    dff g1525(.RN(n1), .SN(1'b1), .CK(n0), .D(n1542), .Q(n34[27]));
    nand g1526(n1453 ,n180 ,n389);
    dff g1527(.RN(n1), .SN(1'b1), .CK(n0), .D(n1820), .Q(n29[2]));
    nand g1528(n1392 ,n164 ,n364);
    nand g1529(n1199 ,n30[28] ,n54);
    buf g1530(n14[13], n11[13]);
    dff g1531(.RN(n1), .SN(1'b1), .CK(n0), .D(n1814), .Q(n32[13]));
    or g1532(n467 ,n338 ,n350);
    xnor g1533(n277 ,n29[25] ,n30[25]);
    dff g1534(.RN(n1), .SN(1'b1), .CK(n0), .D(n1596), .Q(n30[16]));
    dff g1535(.RN(n1), .SN(1'b1), .CK(n0), .D(n1813), .Q(n32[12]));
    nand g1536(n1772 ,n614 ,n1650);
    nand g1537(n1159 ,n30[26] ,n351);
    nand g1538(n1071 ,n32[28] ,n46);
    dff g1539(.RN(n1), .SN(1'b1), .CK(n0), .D(n1674), .Q(n22[3]));
    buf g1540(n16[2], n15[10]);
    nand g1541(n1497 ,n1129 ,n603);
    nand g1542(n1357 ,n1002 ,n530);
    nand g1543(n237 ,n28[18] ,n32[18]);
    nand g1544(n1246 ,n24[16] ,n348);
    nand g1545(n753 ,n31[29] ,n41);
    nand g1546(n728 ,n26[27] ,n354);
    nand g1547(n1121 ,n28[19] ,n350);
    nand g1548(n561 ,n22[2] ,n355);
    nand g1549(n598 ,n21[18] ,n52);
    nand g1550(n760 ,n34[5] ,n353);
    nand g1551(n735 ,n33[31] ,n50);
    xor g1552(n19[5] ,n21[5] ,n22[5]);
    or g1553(n452 ,n309 ,n50);
    nand g1554(n211 ,n29[27] ,n30[27]);
    xor g1555(n20[2] ,n23[2] ,n24[2]);
    nand g1556(n1463 ,n1107 ,n588);
    nand g1557(n834 ,n26[6] ,n354);
    nand g1558(n1489 ,n757 ,n1123);
    dff g1559(.RN(n1), .SN(1'b1), .CK(n0), .D(n1618), .Q(n33[20]));
    nand g1560(n1882 ,n19[5] ,n1865);
    nand g1561(n667 ,n13[1] ,n345);
    nand g1562(n604 ,n21[12] ,n52);
    nand g1563(n1031 ,n26[24] ,n45);
    nand g1564(n927 ,n9[3] ,n349);
    nand g1565(n1629 ,n881 ,n1195);
    dff g1566(.RN(n1), .SN(1'b1), .CK(n0), .D(n1838), .Q(n29[16]));
    nor g1567(n531 ,n144 ,n351);
    nand g1568(n811 ,n35[5] ,n356);
    dff g1569(.RN(n1), .SN(1'b1), .CK(n0), .D(n1601), .Q(n30[15]));
    nand g1570(n1505 ,n764 ,n1130);
    nand g1571(n999 ,n35[15] ,n356);
    nor g1572(n823 ,n163 ,n342);
    nand g1573(n1695 ,n1253 ,n948);
    nor g1574(n550 ,n18[0] ,n358);
    nand g1575(n868 ,n11[6] ,n49);
    nand g1576(n1316 ,n911 ,n429);
    nand g1577(n1831 ,n1026 ,n1399);
    nand g1578(n829 ,n34[19] ,n41);
    nand g1579(n1001 ,n15[9] ,n354);
    nand g1580(n1556 ,n829 ,n1173);
    nand g1581(n644 ,n21[20] ,n347);
    nand g1582(n596 ,n21[20] ,n52);
    nand g1583(n1202 ,n35[27] ,n44);
    nand g1584(n1397 ,n676 ,n627);
    dff g1585(.RN(n1), .SN(1'b1), .CK(n0), .D(n1829), .Q(n29[10]));
    or g1586(n379 ,n306 ,n351);
    nand g1587(n1811 ,n1106 ,n1465);
    nand g1588(n1796 ,n793 ,n1520);
    nor g1589(n82 ,n21[11] ,n24[11]);
    nand g1590(n1490 ,n1124 ,n599);
    or g1591(n473 ,n315 ,n353);
    nand g1592(n228 ,n31[29] ,n34[29]);
    or g1593(n477 ,n327 ,n49);
    nand g1594(n594 ,n21[22] ,n52);
    or g1595(n551 ,n7[3] ,n360);
    xor g1596(n20[3] ,n23[3] ,n24[3]);
    dff g1597(.RN(n1), .SN(1'b1), .CK(n0), .D(n1798), .Q(n31[10]));
    nand g1598(n1630 ,n886 ,n1220);
    nand g1599(n152 ,n27[0] ,n2);
    nand g1600(n1188 ,n30[20] ,n351);
    nand g1601(n217 ,n28[10] ,n32[10]);
    nand g1602(n1656 ,n951 ,n665);
    nand g1603(n1052 ,n33[30] ,n355);
    nand g1604(n1264 ,n24[2] ,n51);
    nor g1605(n523 ,n119 ,n351);
    dff g1606(.RN(n1), .SN(1'b1), .CK(n0), .D(n1301), .Q(n35[24]));
    nand g1607(n1710 ,n1266 ,n960);
    nand g1608(n1340 ,n897 ,n477);
    dff g1609(.RN(n1), .SN(1'b1), .CK(n0), .D(n1337), .Q(n34[1]));
    nor g1610(n1910 ,n1871 ,n1884);
    buf g1611(n16[6], n15[2]);
    xnor g1612(n311 ,n30[3] ,n29[3]);
    nand g1613(n946 ,n4[6] ,n349);
    nand g1614(n910 ,n10[2] ,n356);
    nand g1615(n1661 ,n1233 ,n941);
    nand g1616(n1070 ,n29[5] ,n351);
    nand g1617(n920 ,n5[27] ,n349);
    xnor g1618(n307 ,n30[1] ,n29[1]);
    dff g1619(.RN(n1), .SN(1'b1), .CK(n0), .D(n1350), .Q(n13[19]));
    or g1620(n464 ,n310 ,n41);
    nand g1621(n619 ,n32[3] ,n350);
    nand g1622(n1704 ,n1260 ,n957);
    nand g1623(n1641 ,n158 ,n454);
    nand g1624(n1338 ,n861 ,n473);
    nand g1625(n676 ,n11[31] ,n50);
    or g1626(n382 ,n305 ,n46);
    nand g1627(n1072 ,n30[14] ,n47);
    nand g1628(n626 ,n30[0] ,n351);
    or g1629(n441 ,n269 ,n353);
    dff g1630(.RN(n1), .SN(1'b1), .CK(n0), .D(n1719), .Q(n14[0]));
    buf g1631(n12[6], n11[6]);
    nand g1632(n888 ,n4[14] ,n349);
    dff g1633(.RN(n1), .SN(1'b1), .CK(n0), .D(n1668), .Q(n22[5]));
    not g1634(n353 ,n54);
    dff g1635(.RN(n1), .SN(1'b1), .CK(n0), .D(n1701), .Q(n24[5]));
    nand g1636(n776 ,n31[16] ,n353);
    dff g1637(.RN(n1), .SN(1'b1), .CK(n0), .D(n1539), .Q(n34[30]));
    nand g1638(n1173 ,n30[19] ,n54);
    nand g1639(n850 ,n32[19] ,n53);
    xnor g1640(n333 ,n21[23] ,n24[23]);
    xnor g1641(n293 ,n26[19] ,n33[15]);
    nand g1642(n955 ,n5[6] ,n349);
    nand g1643(n1778 ,n1224 ,n1637);
    nand g1644(n1522 ,n167 ,n448);
    nand g1645(n1646 ,n651 ,n902);
    nor g1646(n114 ,n28[28] ,n32[28]);
    dff g1647(.RN(n1), .SN(1'b1), .CK(n0), .D(n1681), .Q(n24[18]));
    nand g1648(n1311 ,n808 ,n460);
    nand g1649(n239 ,n29[13] ,n30[13]);
    nand g1650(n1610 ,n645 ,n723);
    nand g1651(n602 ,n21[14] ,n52);
    dff g1652(.RN(n1), .SN(1'b1), .CK(n0), .D(n1493), .Q(n26[15]));
    dff g1653(.RN(n1), .SN(1'b1), .CK(n0), .D(n1776), .Q(n33[6]));
    dff g1654(.RN(n1), .SN(1'b1), .CK(n0), .D(n1538), .Q(n21[31]));
    or g1655(n412 ,n318 ,n46);
    dff g1656(.RN(n1), .SN(1'b1), .CK(n0), .D(n1505), .Q(n26[14]));
    nand g1657(n929 ,n5[22] ,n43);
    dff g1658(.RN(n1), .SN(1'b1), .CK(n0), .D(n1655), .Q(n10[1]));
    nand g1659(n934 ,n9[1] ,n43);
    nand g1660(n600 ,n21[16] ,n52);
    buf g1661(n16[14], 1'b0);
    nand g1662(n1406 ,n685 ,n1029);
    nand g1663(n1758 ,n986 ,n1727);
    nor g1664(n106 ,n21[29] ,n24[29]);
    dff g1665(.RN(n1), .SN(1'b1), .CK(n0), .D(n1848), .Q(n27[0]));
    dff g1666(.RN(n1), .SN(1'b1), .CK(n0), .D(n1457), .Q(n26[24]));
    not g1667(n60 ,n27[0]);
    or g1668(n1875 ,n21[9] ,n21[8]);
    or g1669(n410 ,n316 ,n350);
    nand g1670(n1799 ,n771 ,n1746);
    dff g1671(.RN(n1), .SN(1'b1), .CK(n0), .D(n1312), .Q(n35[3]));
    nand g1672(n1268 ,n29[28] ,n351);
    nand g1673(n1669 ,n1236 ,n923);
    dff g1674(.RN(n1), .SN(1'b1), .CK(n0), .D(n1665), .Q(n21[6]));
    xnor g1675(n335 ,n32[3] ,n28[3]);
    nor g1676(n389 ,n73 ,n350);
    dff g1677(.RN(n1), .SN(1'b1), .CK(n0), .D(n1827), .Q(n32[29]));
    dff g1678(.RN(n1), .SN(1'b1), .CK(n0), .D(n1362), .Q(n29[15]));
    nor g1679(n123 ,n28[8] ,n32[8]);
    nor g1680(n1880 ,n1862 ,n21[28]);
    dff g1681(.RN(n1), .SN(1'b1), .CK(n0), .D(n1380), .Q(n28[3]));
    nand g1682(n1320 ,n758 ,n422);
    nor g1683(n67 ,n31[19] ,n34[19]);
    buf g1684(n12[2], n11[30]);
    nand g1685(n1186 ,n30[21] ,n351);
    nand g1686(n1241 ,n24[20] ,n347);
    or g1687(n510 ,n285 ,n49);
    nor g1688(n420 ,n92 ,n353);
    nand g1689(n1365 ,n1062 ,n369);
    dff g1690(.RN(n1), .SN(1'b1), .CK(n0), .D(n1416), .Q(n11[18]));
    not g1691(n1867 ,n24[14]);
    dff g1692(.RN(n1), .SN(1'b1), .CK(n0), .D(n1736), .Q(n25[28]));
    nand g1693(n965 ,n3[30] ,n349);
    nor g1694(n445 ,n70 ,n356);
    nand g1695(n1249 ,n24[13] ,n348);
    dff g1696(.RN(n1), .SN(1'b1), .CK(n0), .D(n1610), .Q(n21[18]));
    nand g1697(n1410 ,n691 ,n1035);
    nand g1698(n804 ,n31[5] ,n353);
    nand g1699(n1010 ,n13[7] ,n50);
    nand g1700(n1342 ,n905 ,n482);
    nand g1701(n1137 ,n28[9] ,n350);
    dff g1702(.RN(n1), .SN(1'b1), .CK(n0), .D(n1419), .Q(n11[16]));
    nor g1703(n128 ,n31[16] ,n34[16]);
    nand g1704(n810 ,n4[24] ,n43);
    xnor g1705(n287 ,n28[23] ,n32[23]);
    nand g1706(n1671 ,n564 ,n925);
    nand g1707(n1471 ,n234 ,n407);
    nand g1708(n992 ,n15[11] ,n354);
    dff g1709(.RN(n1), .SN(1'b1), .CK(n0), .D(n1422), .Q(n11[14]));
    or g1710(n411 ,n317 ,n46);
    nand g1711(n1003 ,n33[16] ,n344);
    dff g1712(.RN(n1), .SN(1'b1), .CK(n0), .D(n1646), .Q(n21[10]));
    buf g1713(n12[12], n11[12]);
    dff g1714(.RN(n1), .SN(1'b1), .CK(n0), .D(n1587), .Q(n26[5]));
    xor g1715(n358 ,n21[0] ,n23[0]);
    dff g1716(.RN(n1), .SN(1'b1), .CK(n0), .D(n1608), .Q(n30[13]));
    nand g1717(n1819 ,n1086 ,n1452);
    xnor g1718(n302 ,n21[8] ,n24[8]);
    nand g1719(n666 ,n36[3] ,n56);
    dff g1720(.RN(n1), .SN(1'b1), .CK(n0), .D(n1826), .Q(n32[28]));
    nand g1721(n931 ,n5[21] ,n43);
    nand g1722(n1403 ,n681 ,n1027);
    nand g1723(n856 ,n4[21] ,n43);
    nand g1724(n1219 ,n35[16] ,n346);
    nand g1725(n1663 ,n565 ,n942);
    nand g1726(n210 ,n28[31] ,n32[31]);
    nor g1727(n97 ,n29[19] ,n30[19]);
    nand g1728(n1881 ,n24[5] ,n1858);
    dff g1729(.RN(n1), .SN(1'b1), .CK(n0), .D(n1664), .Q(n24[28]));
    nand g1730(n738 ,n34[1] ,n352);
    nand g1731(n587 ,n21[29] ,n52);
    nand g1732(n1184 ,n30[8] ,n54);
    dff g1733(.RN(n1), .SN(1'b1), .CK(n0), .D(n1763), .Q(n29[26]));
    nand g1734(n1075 ,n29[4] ,n47);
    dff g1735(.RN(n1), .SN(1'b1), .CK(n0), .D(n1581), .Q(n34[7]));
    xnor g1736(n316 ,n21[3] ,n24[3]);
    nand g1737(n986 ,n13[21] ,n50);
    nand g1738(n1540 ,n638 ,n877);
    nand g1739(n1195 ,n33[3] ,n355);
    dff g1740(.RN(n1), .SN(1'b1), .CK(n0), .D(n1800), .Q(n31[12]));
    nand g1741(n1212 ,n35[20] ,n45);
    nor g1742(n439 ,n116 ,n352);
    nand g1743(n889 ,n4[13] ,n349);
    dff g1744(.RN(n1), .SN(1'b1), .CK(n0), .D(n1699), .Q(n24[7]));
    nand g1745(n1430 ,n712 ,n1054);
    dff g1746(.RN(n1), .SN(1'b1), .CK(n0), .D(n1796), .Q(n35[19]));
    nand g1747(n1069 ,n32[29] ,n350);
    nand g1748(n1727 ,n230 ,n517);
    nand g1749(n1835 ,n574 ,n1287);
    nand g1750(n1838 ,n824 ,n1742);
    nand g1751(n1113 ,n28[24] ,n46);
    dff g1752(.RN(n1), .SN(1'b1), .CK(n0), .D(n1386), .Q(n29[21]));
    buf g1753(n14[20], n11[20]);
    nand g1754(n786 ,n34[11] ,n353);
    nand g1755(n1279 ,n29[21] ,n48);
    dff g1756(.RN(n1), .SN(1'b1), .CK(n0), .D(n1417), .Q(n11[17]));
    nand g1757(n1237 ,n24[24] ,n51);
    nand g1758(n1550 ,n842 ,n1163);
    nor g1759(n1518 ,n162 ,n572);
    nand g1760(n1209 ,n35[22] ,n45);
    nand g1761(n1019 ,n13[2] ,n49);
    nor g1762(n1929 ,n1926 ,n1920);
    dff g1763(.RN(n1), .SN(1'b1), .CK(n0), .D(n1319), .Q(n31[29]));
    nor g1764(n1913 ,n1899 ,n1890);
    dff g1765(.RN(n1), .SN(1'b1), .CK(n0), .D(n1614), .Q(n21[17]));
    nand g1766(n1384 ,n1276 ,n512);
    nand g1767(n1609 ,n709 ,n1205);
    nand g1768(n1568 ,n806 ,n1177);
    nand g1769(n820 ,n35[0] ,n356);
    nand g1770(n1065 ,n32[31] ,n46);
    nand g1771(n739 ,n26[21] ,n354);
    nand g1772(n1427 ,n708 ,n1051);
    or g1773(n522 ,n292 ,n50);
    dff g1774(.RN(n1), .SN(1'b1), .CK(n0), .D(n1435), .Q(n11[3]));
    nand g1775(n693 ,n11[19] ,n49);
    xnor g1776(n332 ,n22[2] ,n32[2]);
    dff g1777(.RN(n1), .SN(1'b1), .CK(n0), .D(n1667), .Q(n24[26]));
    not g1778(n349 ,n51);
    nand g1779(n1527 ,n207 ,n457);
    xnor g1780(n266 ,n31[23] ,n34[23]);
    not g1781(n1859 ,n21[24]);
    dff g1782(.RN(n1), .SN(1'b1), .CK(n0), .D(n1474), .Q(n28[24]));
    xnor g1783(n321 ,n21[2] ,n23[2]);
    nand g1784(n595 ,n21[21] ,n52);
    nand g1785(n1285 ,n34[17] ,n353);
    not g1786(n1864 ,n24[19]);
    nand g1787(n565 ,n22[6] ,n51);
    buf g1788(n16[13], 1'b0);
    xnor g1789(n305 ,n21[24] ,n24[24]);
    nand g1790(n1058 ,n26[5] ,n44);
    nand g1791(n1130 ,n33[14] ,n55);
    or g1792(n384 ,n333 ,n350);
    dff g1793(.RN(n1), .SN(1'b1), .CK(n0), .D(n1561), .Q(n21[27]));
    nand g1794(n1519 ,n179 ,n446);
    or g1795(n444 ,n320 ,n46);
    dff g1796(.RN(n1), .SN(1'b1), .CK(n0), .D(n1407), .Q(n11[24]));
    nand g1797(n1677 ,n558 ,n930);
    dff g1798(.RN(n1), .SN(1'b1), .CK(n0), .D(n1617), .Q(n33[21]));
    dff g1799(.RN(n1), .SN(1'b1), .CK(n0), .D(n1506), .Q(n28[7]));
    nor g1800(n511 ,n65 ,n50);
    dff g1801(.RN(n1), .SN(1'b1), .CK(n0), .D(n1658), .Q(n24[31]));
    nand g1802(n830 ,n32[28] ,n53);
    nand g1803(n1077 ,n33[26] ,n355);
    nand g1804(n656 ,n21[6] ,n51);
    dff g1805(.RN(n1), .SN(1'b1), .CK(n0), .D(n1819), .Q(n32[20]));
    dff g1806(.RN(n1), .SN(1'b1), .CK(n0), .D(n1382), .Q(n30[4]));
    nand g1807(n659 ,n36[3] ,n355);
    nand g1808(n731 ,n26[24] ,n354);
    nand g1809(n1922 ,n1915 ,n1903);
    nor g1810(n55 ,n40 ,n39);
    xnor g1811(n36[3] ,n1933 ,n25[31]);
    nand g1812(n1794 ,n795 ,n1522);
    dff g1813(.RN(n1), .SN(1'b1), .CK(n0), .D(n1730), .Q(n15[11]));
    dff g1814(.RN(n1), .SN(1'b1), .CK(n0), .D(n1432), .Q(n11[6]));
    nand g1815(n1045 ,n26[14] ,n44);
    nand g1816(n798 ,n35[14] ,n356);
    nand g1817(n701 ,n33[24] ,n49);
    nand g1818(n1524 ,n233 ,n409);
    nand g1819(n197 ,n26[28] ,n33[24]);
    dff g1820(.RN(n1), .SN(1'b1), .CK(n0), .D(n1769), .Q(n29[30]));
    nand g1821(n1680 ,n1243 ,n933);
    nand g1822(n1319 ,n753 ,n419);
    nand g1823(n1666 ,n1234 ,n920);
    dff g1824(.RN(n1), .SN(1'b1), .CK(n0), .D(n1797), .Q(n35[20]));
    dff g1825(.RN(n1), .SN(1'b1), .CK(n0), .D(n1552), .Q(n34[22]));
    dff g1826(.RN(n1), .SN(1'b1), .CK(n0), .D(n1780), .Q(n34[2]));
    xnor g1827(n294 ,n26[18] ,n33[14]);
    nand g1828(n1413 ,n692 ,n1036);
    dff g1829(.RN(n1), .SN(1'b1), .CK(n0), .D(n1548), .Q(n34[24]));
    dff g1830(.RN(n1), .SN(1'b1), .CK(n0), .D(n1334), .Q(n31[3]));
    nand g1831(n1284 ,n29[17] ,n47);
    nand g1832(n1815 ,n1096 ,n1456);
    nand g1833(n157 ,n22[6] ,n32[6]);
    nand g1834(n853 ,n32[18] ,n53);
    nand g1835(n1461 ,n1100 ,n586);
    dff g1836(.RN(n1), .SN(1'b1), .CK(n0), .D(n1549), .Q(n30[29]));
    xnor g1837(n20[0] ,n1852 ,n18[0]);
    nand g1838(n1451 ,n729 ,n1077);
    not g1839(n56 ,n356);
    nand g1840(n1351 ,n990 ,n520);
    nor g1841(n474 ,n124 ,n351);
    nand g1842(n871 ,n34[31] ,n353);
    nand g1843(n1725 ,n197 ,n513);
    xnor g1844(n265 ,n26[31] ,n33[27]);
    nand g1845(n922 ,n5[26] ,n43);
    or g1846(n434 ,n263 ,n352);
    or g1847(n405 ,n303 ,n46);
    or g1848(n494 ,n280 ,n42);
    nor g1849(n129 ,n22[6] ,n32[6]);
    nand g1850(n790 ,n4[23] ,n349);
    dff g1851(.RN(n1), .SN(1'b1), .CK(n0), .D(n1421), .Q(n15[0]));
    nand g1852(n1742 ,n235 ,n539);
    nand g1853(n1208 ,n35[23] ,n346);
    nand g1854(n1830 ,n1037 ,n1411);
    nand g1855(n223 ,n28[11] ,n32[11]);
    nand g1856(n678 ,n15[2] ,n354);
    buf g1857(n17[4], 1'b0);
    dff g1858(.RN(n1), .SN(1'b1), .CK(n0), .D(n1323), .Q(n31[22]));
    nand g1859(n1486 ,n1122 ,n598);
    nand g1860(n1824 ,n1073 ,n1444);
    nand g1861(n836 ,n34[21] ,n352);
    nand g1862(n1575 ,n777 ,n1162);
    nand g1863(n1026 ,n29[13] ,n351);
    nand g1864(n643 ,n21[29] ,n51);
    dff g1865(.RN(n1), .SN(1'b1), .CK(n0), .D(n1799), .Q(n35[21]));
    nand g1866(n1156 ,n33[8] ,n55);
    xnor g1867(n281 ,n28[12] ,n32[12]);
    nand g1868(n706 ,n26[30] ,n354);
    nand g1869(n1634 ,n904 ,n1230);
    nand g1870(n716 ,n11[3] ,n50);
    or g1871(n367 ,n294 ,n49);
    nand g1872(n1595 ,n634 ,n856);
    or g1873(n391 ,n322 ,n350);
    nand g1874(n940 ,n35[10] ,n356);
    nor g1875(n376 ,n108 ,n350);
    nand g1876(n899 ,n33[6] ,n49);
    xnor g1877(n283 ,n28[25] ,n32[25]);
    nand g1878(n1734 ,n237 ,n531);
    buf g1879(n14[6], n11[30]);
    dff g1880(.RN(n1), .SN(1'b1), .CK(n0), .D(n1540), .Q(n21[30]));
    nand g1881(n771 ,n35[21] ,n356);
    nor g1882(n413 ,n137 ,n350);
    nand g1883(n1498 ,n1132 ,n604);
    or g1884(n392 ,n299 ,n46);
    buf g1885(n14[7], n11[31]);
    nand g1886(n206 ,n28[28] ,n32[28]);
    nor g1887(n378 ,n104 ,n46);
    nand g1888(n884 ,n4[15] ,n349);
    xnor g1889(n325 ,n22[4] ,n35[4]);
    or g1890(n489 ,n331 ,n47);
    nand g1891(n886 ,n33[14] ,n50);
    nand g1892(n1259 ,n24[5] ,n51);
    xnor g1893(n260 ,n29[18] ,n30[18]);
    nor g1894(n146 ,n31[11] ,n34[11]);
    nand g1895(n1473 ,n1112 ,n591);
    nor g1896(n1905 ,n1883 ,n1881);
    dff g1897(.RN(n1), .SN(1'b1), .CK(n0), .D(n1616), .Q(n30[11]));
    nand g1898(n238 ,n26[10] ,n33[6]);
    nand g1899(n1608 ,n1204 ,n870);
    buf g1900(n12[7], n11[7]);
    nand g1901(n763 ,n31[23] ,n352);
    nand g1902(n1315 ,n940 ,n494);
    nor g1903(n53 ,n39 ,n37);
    nand g1904(n1714 ,n579 ,n964);
    nand g1905(n180 ,n21[19] ,n24[19]);
    nand g1906(n1236 ,n24[25] ,n51);
    or g1907(n395 ,n300 ,n350);
    nand g1908(n227 ,n33[28] ,n36[0]);
    buf g1909(n14[19], n11[19]);
    not g1910(n1865 ,n19[4]);
    nand g1911(n1523 ,n236 ,n450);
    nand g1912(n1356 ,n998 ,n525);
    nand g1913(n1644 ,n188 ,n479);
    nand g1914(n1625 ,n1003 ,n1219);
    nand g1915(n1225 ,n35[10] ,n44);
    nand g1916(n1836 ,n573 ,n1516);
    nand g1917(n1454 ,n181 ,n393);
    xnor g1918(n328 ,n22[0] ,n32[0]);
    nand g1919(n1712 ,n584 ,n963);
    buf g1920(n14[10], n11[10]);
    dff g1921(.RN(n1), .SN(1'b1), .CK(n0), .D(n1405), .Q(n11[26]));
    or g1922(n495 ,n311 ,n352);
    nand g1923(n1028 ,n26[26] ,n45);
    nand g1924(n1442 ,n725 ,n1067);
    nand g1925(n1322 ,n762 ,n424);
    xnor g1926(n296 ,n31[27] ,n34[27]);
    nand g1927(n1480 ,n1118 ,n595);
    or g1928(n538 ,n244 ,n49);
    xnor g1929(n249 ,n26[23] ,n33[19]);
    or g1930(n535 ,n297 ,n42);
    or g1931(n525 ,n282 ,n345);
    nand g1932(n840 ,n34[12] ,n41);
    nand g1933(n581 ,n21[2] ,n348);
    or g1934(n534 ,n284 ,n50);
    dff g1935(.RN(n1), .SN(1'b1), .CK(n0), .D(n1341), .Q(n33[4]));
    nor g1936(n1286 ,n27[2] ,n823);
    xnor g1937(n312 ,n36[3] ,n33[31]);
    dff g1938(.RN(n1), .SN(1'b1), .CK(n0), .D(n1393), .Q(n12[30]));
    nand g1939(n755 ,n33[17] ,n49);
    nand g1940(n1441 ,n170 ,n373);
    nand g1941(n1394 ,n673 ,n1024);
    nand g1942(n1596 ,n1196 ,n860);
    nand g1943(n1526 ,n221 ,n456);
    dff g1944(.RN(n1), .SN(1'b1), .CK(n0), .D(n1645), .Q(n21[11]));
    nand g1945(n1074 ,n33[27] ,n355);
    or g1946(n424 ,n255 ,n353);
    nand g1947(n1283 ,n29[18] ,n48);
    nand g1948(n1124 ,n28[17] ,n46);
    dff g1949(.RN(n1), .SN(1'b1), .CK(n0), .D(n1687), .Q(n21[3]));
    nand g1950(n1842 ,n2 ,n1834);
    nand g1951(n201 ,n26[4] ,n33[0]);
    dff g1952(.RN(n1), .SN(1'b1), .CK(n0), .D(n1704), .Q(n24[4]));
    nand g1953(n639 ,n21[26] ,n348);
    nor g1954(n398 ,n79 ,n46);
    nand g1955(n1795 ,n792 ,n1519);
    nand g1956(n1637 ,n157 ,n486);
    dff g1957(.RN(n1), .SN(1'b1), .CK(n0), .D(n1577), .Q(n30[22]));
    dff g1958(.RN(n1), .SN(1'b1), .CK(n0), .D(n1698), .Q(n24[8]));
    or g1959(n428 ,n259 ,n352);
    nand g1960(n634 ,n21[21] ,n348);
    buf g1961(n12[8], n11[8]);
    nand g1962(n936 ,n5[18] ,n349);
    nor g1963(n373 ,n113 ,n351);
    or g1964(n512 ,n261 ,n48);
    nand g1965(n874 ,n33[22] ,n50);
    buf g1966(n14[16], n11[16]);
    nand g1967(n1536 ,n209 ,n546);
    dff g1968(.RN(n1), .SN(1'b1), .CK(n0), .D(n1807), .Q(n31[27]));
    dff g1969(.RN(n1), .SN(1'b1), .CK(n0), .D(n1298), .Q(n30[1]));
    or g1970(n451 ,n291 ,n41);
    or g1971(n521 ,n290 ,n47);
    nand g1972(n1679 ,n655 ,n924);
    nand g1973(n1158 ,n30[29] ,n54);
    nor g1974(n109 ,n31[28] ,n34[28]);
    nand g1975(n1474 ,n1113 ,n592);
    nand g1976(n1280 ,n29[20] ,n47);
    dff g1977(.RN(n1), .SN(1'b1), .CK(n0), .D(n1598), .Q(n21[20]));
    nand g1978(n1103 ,n28[29] ,n46);
    nand g1979(n1057 ,n33[29] ,n355);
    nand g1980(n161 ,n18[0] ,n33[0]);
    nand g1981(n1185 ,n30[7] ,n54);
    nand g1982(n1348 ,n982 ,n514);
    nand g1983(n1192 ,n30[18] ,n47);
    nand g1984(n1377 ,n1091 ,n395);
    dff g1985(.RN(n1), .SN(1'b1), .CK(n0), .D(n1745), .Q(n26[12]));
    nand g1986(n1020 ,n29[15] ,n351);
    nand g1987(n1250 ,n24[12] ,n347);
    nand g1988(n1513 ,n200 ,n439);
    dff g1989(.RN(n1), .SN(1'b1), .CK(n0), .D(n1811), .Q(n32[9]));
    nand g1990(n1817 ,n1093 ,n1455);
    nand g1991(n795 ,n31[8] ,n353);
    dff g1992(.RN(n1), .SN(1'b1), .CK(n0), .D(n1400), .Q(n11[29]));
    nand g1993(n663 ,n36[2] ,n56);
    nand g1994(n638 ,n21[30] ,n348);
    dff g1995(.RN(n1), .SN(1'b1), .CK(n0), .D(n1832), .Q(n29[14]));
    nand g1996(n1024 ,n26[29] ,n44);
    nand g1997(n231 ,n26[12] ,n33[8]);
    nand g1998(n654 ,n21[7] ,n51);
    dff g1999(.RN(n1), .SN(1'b1), .CK(n0), .D(n1469), .Q(n26[20]));
    dff g2000(.RN(n1), .SN(1'b1), .CK(n0), .D(n1791), .Q(n35[13]));
    nand g2001(n1829 ,n1043 ,n1418);
    buf g2002(n12[22], n11[22]);
    dff g2003(.RN(n1), .SN(1'b1), .CK(n0), .D(n1343), .Q(n13[31]));
    dff g2004(.RN(n1), .SN(1'b1), .CK(n0), .D(n1824), .Q(n32[27]));
    nand g2005(n641 ,n21[25] ,n347);
    nand g2006(n589 ,n21[27] ,n52);
    nand g2007(n1422 ,n700 ,n1045);
    nand g2008(n1004 ,n13[10] ,n345);
    nor g2009(n103 ,n31[20] ,n34[20]);
    nand g2010(n1774 ,n907 ,n1647);
    nand g2011(n650 ,n21[11] ,n51);
    xnor g2012(n290 ,n28[21] ,n32[21]);
    nand g2013(n1141 ,n30[24] ,n54);
    dff g2014(.RN(n1), .SN(1'b1), .CK(n0), .D(n1326), .Q(n31[18]));
    nand g2015(n560 ,n22[3] ,n355);
    dff g2016(.RN(n1), .SN(1'b1), .CK(n0), .D(n1504), .Q(n28[8]));
    dff g2017(.RN(n1), .SN(1'b1), .CK(n0), .D(n1508), .Q(n26[13]));
    or g2018(n438 ,n296 ,n356);
    nand g2019(n1503 ,n759 ,n1128);
    dff g2020(.RN(n1), .SN(1'b1), .CK(n0), .D(n1490), .Q(n28[17]));
    nand g2021(n1160 ,n30[31] ,n351);
    nand g2022(n1741 ,n240 ,n541);
    nand g2023(n1452 ,n178 ,n388);
    dff g2024(.RN(n1), .SN(1'b1), .CK(n0), .D(n1717), .Q(n14[1]));
    nor g2025(n52 ,n38 ,n37);
    dff g2026(.RN(n1), .SN(1'b1), .CK(n0), .D(n1580), .Q(n30[21]));
    dff g2027(.RN(n1), .SN(1'b1), .CK(n0), .D(n1387), .Q(n29[19]));
    nand g2028(n1265 ,n25[28] ,n348);
    nand g2029(n571 ,n22[5] ,n355);
    nand g2030(n759 ,n26[16] ,n354);
    nand g2031(n1390 ,n201 ,n363);
    nand g2032(n717 ,n11[2] ,n344);
    nand g2033(n967 ,n35[27] ,n356);
    nand g2034(n1694 ,n581 ,n939);
    or g2035(n149 ,n60 ,n2);
    not g2036(n1861 ,n24[6]);
    nand g2037(n1759 ,n983 ,n1726);
    or g2038(n422 ,n254 ,n352);
    nand g2039(n660 ,n36[2] ,n355);
    nand g2040(n582 ,n21[3] ,n347);
    nand g2041(n205 ,n31[13] ,n34[13]);
    nand g2042(n689 ,n11[22] ,n50);
    nand g2043(n1180 ,n30[11] ,n54);
    or g2044(n431 ,n260 ,n353);
    nand g2045(n1203 ,n35[26] ,n45);
    or g2046(n475 ,n273 ,n356);
    or g2047(n1844 ,n1748 ,n1839);
    nand g2048(n909 ,n4[8] ,n43);
    dff g2049(.RN(n1), .SN(1'b1), .CK(n0), .D(n1621), .Q(n33[18]));
    or g2050(n459 ,n278 ,n356);
    nor g2051(n386 ,n76 ,n351);
    nor g2052(n399 ,n80 ,n46);
    nor g2053(n119 ,n28[20] ,n32[20]);
    xnor g2054(n329 ,n22[3] ,n32[3]);
    nor g2055(n461 ,n130 ,n356);
    xnor g2056(n245 ,n28[9] ,n32[9]);
    dff g2057(.RN(n1), .SN(1'b1), .CK(n0), .D(n1603), .Q(n33[28]));
    nand g2058(n1106 ,n32[9] ,n46);
    nand g2059(n913 ,n4[7] ,n349);
    dff g2060(.RN(n1), .SN(1'b1), .CK(n0), .D(n1313), .Q(n35[2]));
    nand g2061(n775 ,n31[17] ,n41);
    nand g2062(n1239 ,n24[22] ,n347);
    nand g2063(n780 ,n34[9] ,n352);
    nand g2064(n1789 ,n950 ,n1527);
    nor g2065(n151 ,n21[26] ,n24[26]);
    dff g2066(.RN(n1), .SN(1'b1), .CK(n0), .D(n1466), .Q(n26[23]));
    nand g2067(n724 ,n33[28] ,n49);
    nand g2068(n1640 ,n895 ,n1227);
    dff g2069(.RN(n1), .SN(1'b1), .CK(n0), .D(n1433), .Q(n11[5]));
    nor g2070(n549 ,n18[1] ,n361);
    nand g2071(n1153 ,n28[4] ,n46);
    nand g2072(n1883 ,n24[7] ,n1861);
    nand g2073(n1114 ,n28[23] ,n350);
    dff g2074(.RN(n1), .SN(1'b1), .CK(n0), .D(n1774), .Q(n33[2]));
    dff g2075(.RN(n1), .SN(1'b1), .CK(n0), .D(n1303), .Q(n35[25]));
    nand g2076(n1552 ,n803 ,n1178);
    nand g2077(n1039 ,n26[18] ,n45);
    nand g2078(n841 ,n32[23] ,n53);
    nand g2079(n1136 ,n30[15] ,n351);
    nand g2080(n939 ,n4[2] ,n43);
    or g2081(n491 ,n271 ,n356);
    dff g2082(.RN(n1), .SN(1'b1), .CK(n0), .D(n1335), .Q(n31[2]));
    buf g2083(n12[15], n11[15]);
    dff g2084(.RN(n1), .SN(1'b1), .CK(n0), .D(n1395), .Q(n15[4]));
    dff g2085(.RN(n1), .SN(1'b1), .CK(n0), .D(n1384), .Q(n29[24]));
    nand g2086(n727 ,n26[11] ,n354);
    dff g2087(.RN(n1), .SN(1'b1), .CK(n0), .D(n1446), .Q(n26[27]));
    nor g2088(n503 ,n109 ,n42);
    buf g2089(n12[11], n11[11]);
    nand g2090(n1375 ,n1089 ,n390);
    nand g2091(n997 ,n13[14] ,n50);
    nand g2092(n1079 ,n32[24] ,n350);
    dff g2093(.RN(n1), .SN(1'b1), .CK(n0), .D(n1543), .Q(n30[31]));
    nand g2094(n1606 ,n1072 ,n866);
    dff g2095(.RN(n1), .SN(1'b1), .CK(n0), .D(n1397), .Q(n11[31]));
    nor g2096(n1517 ,n334 ,n551);
    dff g2097(.RN(n1), .SN(1'b1), .CK(n0), .D(n1630), .Q(n33[14]));
    dff g2098(.RN(n1), .SN(1'b1), .CK(n0), .D(n1594), .Q(n30[17]));
    nand g2099(n1329 ,n779 ,n434);
    not g2100(n46 ,n52);
    nor g2101(n104 ,n21[27] ,n24[27]);
    not g2102(n45 ,n50);
    not g2103(n348 ,n43);
    nand g2104(n749 ,n31[31] ,n353);
    nor g2105(n533 ,n141 ,n344);
    nand g2106(n950 ,n35[11] ,n356);
    dff g2107(.RN(n1), .SN(1'b1), .CK(n0), .D(n1331), .Q(n31[11]));
    nor g2108(n1874 ,n19[3] ,n19[2]);
    nor g2109(n400 ,n81 ,n46);
    nand g2110(n187 ,n31[21] ,n34[21]);
    nand g2111(n468 ,n34[28] ,n353);
    nor g2112(n102 ,n22[1] ,n35[1]);
    nor g2113(n496 ,n120 ,n351);
    nand g2114(n1032 ,n26[23] ,n346);
    nand g2115(n1510 ,n239 ,n528);
    nand g2116(n1477 ,n192 ,n413);
    nand g2117(n175 ,n31[1] ,n34[1]);
    nor g2118(n425 ,n95 ,n353);
    dff g2119(.RN(n1), .SN(1'b1), .CK(n0), .D(n1389), .Q(n15[5]));
    nand g2120(n1899 ,n24[27] ,n24[26]);
    dff g2121(.RN(n1), .SN(1'b1), .CK(n0), .D(n1715), .Q(n14[3]));
    nand g2122(n1659 ,n1232 ,n945);
    nand g2123(n1064 ,n26[0] ,n45);
    nand g2124(n954 ,n3[31] ,n349);
    dff g2125(.RN(n1), .SN(1'b1), .CK(n0), .D(n1372), .Q(n32[23]));
    nand g2126(n937 ,n9[0] ,n349);
    nand g2127(n851 ,n34[4] ,n353);
    nand g2128(n178 ,n21[20] ,n24[20]);
    nand g2129(n1011 ,n13[6] ,n49);
    nand g2130(n773 ,n31[18] ,n352);
    xor g2131(n19[4] ,n21[4] ,n22[4]);
    nand g2132(n806 ,n34[13] ,n353);
    nand g2133(n229 ,n26[7] ,n33[3]);
    buf g2134(n15[13], 1'b0);
    nand g2135(n1633 ,n647 ,n888);
    nand g2136(n758 ,n31[26] ,n41);
    dff g2137(.RN(n1), .SN(1'b1), .CK(n0), .D(n490), .Q(n17[0]));
    nand g2138(n1172 ,n30[16] ,n54);
    nand g2139(n1101 ,n33[22] ,n355);
    nand g2140(n792 ,n31[9] ,n352);
    nand g2141(n906 ,n4[9] ,n43);
    nor g2142(n136 ,n29[9] ,n30[9]);
    xnor g2143(n267 ,n31[22] ,n34[22]);
    nand g2144(n150 ,n27[2] ,n57);
    nand g2145(n729 ,n26[26] ,n354);
    or g2146(n426 ,n256 ,n353);
    nand g2147(n1233 ,n24[29] ,n347);
    nand g2148(n235 ,n28[16] ,n32[16]);
    dff g2149(.RN(n1), .SN(1'b1), .CK(n0), .D(n1740), .Q(n15[7]));
    nor g2150(n81 ,n21[12] ,n24[12]);
    buf g2151(n14[9], n11[9]);
    dff g2152(.RN(n1), .SN(1'b1), .CK(n0), .D(n1669), .Q(n24[25]));
    xnor g2153(n255 ,n29[24] ,n30[24]);
    nand g2154(n852 ,n4[28] ,n349);
    nand g2155(n1277 ,n29[23] ,n48);
    nand g2156(n588 ,n21[28] ,n52);
    nand g2157(n1825 ,n1070 ,n1441);
    nor g2158(n117 ,n28[29] ,n32[29]);
    or g2159(n406 ,n314 ,n350);
    nand g2160(n1222 ,n35[13] ,n346);
    nand g2161(n1715 ,n966 ,n553);
    nand g2162(n1261 ,n24[3] ,n51);
    nand g2163(n777 ,n34[25] ,n352);
    dff g2164(.RN(n1), .SN(1'b1), .CK(n0), .D(n1308), .Q(n35[14]));
    nor g2165(n1917 ,n1897 ,n1872);
    nand g2166(n189 ,n21[9] ,n24[9]);
    nor g2167(n1873 ,n19[1] ,n19[0]);
    buf g2168(n16[10], n15[6]);
    buf g2169(n14[12], n11[12]);
    nand g2170(n1743 ,n229 ,n543);
    or g2171(n147 ,n58 ,n2);
    dff g2172(.RN(n1), .SN(1'b1), .CK(n0), .D(n1635), .Q(n33[11]));
    nand g2173(n1662 ,n161 ,n493);
    nand g2174(n1415 ,n693 ,n1038);
    nand g2175(n1221 ,n30[7] ,n48);
    nand g2176(n756 ,n31[27] ,n353);
    buf g2177(n14[5], n11[29]);
    nand g2178(n1612 ,n697 ,n1208);
    nand g2179(n1022 ,n26[30] ,n45);
    nor g2180(n506 ,n105 ,n356);
    nand g2181(n1067 ,n33[28] ,n355);
    buf g2182(n14[27], n11[27]);
    nand g2183(n740 ,n32[31] ,n53);
    nand g2184(n1034 ,n26[22] ,n44);
    xnor g2185(n1849 ,n23[1] ,n24[1]);
    nor g2186(n1888 ,n1854 ,n21[16]);
    dff g2187(.RN(n1), .SN(1'b1), .CK(n0), .D(n1615), .Q(n33[22]));
    or g2188(n1923 ,n1907 ,n1914);
    nand g2189(n1131 ,n33[15] ,n55);
    nand g2190(n578 ,n23[0] ,n51);
    dff g2191(.RN(n1), .SN(1'b1), .CK(n0), .D(n1381), .Q(n28[2]));
    nor g2192(n443 ,n83 ,n353);
    nand g2193(n932 ,n5[28] ,n43);
    nand g2194(n1088 ,n32[18] ,n46);
    nand g2195(n1361 ,n1019 ,n547);
    nand g2196(n1273 ,n33[2] ,n355);
    dff g2197(.RN(n1), .SN(1'b1), .CK(n0), .D(n1425), .Q(n11[11]));
    buf g2198(n12[9], n11[9]);
    xnor g2199(n242 ,n26[15] ,n33[11]);
    nand g2200(n1063 ,n26[1] ,n44);
    nand g2201(n1895 ,n24[22] ,n1853);
    nand g2202(n1401 ,n1007 ,n560);
    dff g2203(.RN(n1), .SN(1'b1), .CK(n0), .D(n1479), .Q(n23[2]));
    nand g2204(n766 ,n32[30] ,n53);
    nor g2205(n1287 ,n350 ,n550);
    nand g2206(n789 ,n35[22] ,n356);
    nand g2207(n714 ,n11[5] ,n345);
    nand g2208(n1300 ,n781 ,n527);
    xnor g2209(n20[1] ,n1849 ,n18[1]);
    nand g2210(n832 ,n32[27] ,n53);
    nand g2211(n1650 ,n215 ,n529);
    nand g2212(n1037 ,n29[11] ,n351);
    nand g2213(n768 ,n4[22] ,n43);
    nand g2214(n559 ,n22[0] ,n348);
    nand g2215(n1620 ,n878 ,n1214);
    nor g2216(n148 ,n57 ,n27[2]);
    dff g2217(.RN(n1), .SN(1'b1), .CK(n0), .D(n1785), .Q(n35[5]));
    nand g2218(n202 ,n31[20] ,n34[20]);
    buf g2219(n12[13], n11[13]);
    nand g2220(n579 ,n18[0] ,n348);
    nand g2221(n224 ,n26[16] ,n33[12]);
    nand g2222(n220 ,n28[29] ,n32[29]);
    nand g2223(n1123 ,n33[17] ,n55);
    nand g2224(n1317 ,n749 ,n416);
    nand g2225(n1462 ,n186 ,n401);
    or g2226(n423 ,n277 ,n352);
    nand g2227(n1006 ,n13[9] ,n49);
    nand g2228(n1162 ,n30[25] ,n54);
    nor g2229(n113 ,n28[5] ,n32[5]);
    xnor g2230(n258 ,n31[24] ,n34[24]);
    buf g2231(n12[14], n11[14]);
    nand g2232(n674 ,n32[9] ,n53);
    nand g2233(n1448 ,n176 ,n385);
    nand g2234(n1197 ,n35[30] ,n45);
    nand g2235(n1030 ,n29[12] ,n47);
    dff g2236(.RN(n1), .SN(1'b1), .CK(n0), .D(n1847), .Q(n27[1]));
    nand g2237(n961 ,n5[0] ,n43);
    nand g2238(n1050 ,n26[10] ,n44);
    nand g2239(n1235 ,n24[26] ,n348);
    nor g2240(n497 ,n135 ,n47);
    dff g2241(.RN(n1), .SN(1'b1), .CK(n0), .D(n1753), .Q(n29[18]));
    nand g2242(n1618 ,n682 ,n1212);
    not g2243(n57 ,n2);
    dff g2244(.RN(n1), .SN(1'b1), .CK(n0), .D(n1464), .Q(n28[29]));
    nand g2245(n1449 ,n177 ,n386);
    nand g2246(n944 ,n5[13] ,n349);
    dff g2247(.RN(n1), .SN(1'b1), .CK(n0), .D(n1659), .Q(n24[30]));
    nand g2248(n207 ,n31[11] ,n34[11]);
    nand g2249(n849 ,n32[20] ,n53);
    or g2250(n547 ,n343 ,n49);
    nand g2251(n878 ,n33[19] ,n345);
    nand g2252(n1446 ,n728 ,n1074);
    nand g2253(n1764 ,n7[1] ,n1518);
    dff g2254(.RN(n1), .SN(1'b1), .CK(n0), .D(n1752), .Q(n13[8]));
    nand g2255(n1405 ,n683 ,n1028);
    dff g2256(.RN(n1), .SN(1'b1), .CK(n0), .D(n1792), .Q(n35[15]));
    nand g2257(n877 ,n4[30] ,n349);
    or g2258(n472 ,n313 ,n50);
    nand g2259(n1525 ,n205 ,n394);
    nand g2260(n1833 ,n670 ,n1390);
    nand g2261(n613 ,n33[1] ,n50);
    nand g2262(n838 ,n26[7] ,n354);
    nor g2263(n83 ,n29[10] ,n30[10]);
    nor g2264(n470 ,n132 ,n41);
    nand g2265(n1685 ,n559 ,n937);
    dff g2266(.RN(n1), .SN(1'b1), .CK(n0), .D(n1708), .Q(n24[2]));
    dff g2267(.RN(n1), .SN(1'b1), .CK(n0), .D(n1696), .Q(n24[9]));
    nand g2268(n770 ,n31[19] ,n352);
    not g2269(n351 ,n53);
    nand g2270(n1730 ,n992 ,n659);
    nand g2271(n1396 ,n675 ,n1025);
    dff g2272(.RN(n1), .SN(1'b1), .CK(n0), .D(n1777), .Q(n30[5]));
    nand g2273(n1713 ,n206 ,n501);
    dff g2274(.RN(n1), .SN(1'b1), .CK(n0), .D(n1678), .Q(n24[20]));
    dff g2275(.RN(n1), .SN(1'b1), .CK(n0), .D(n1461), .Q(n28[30]));
    nand g2276(n1665 ,n656 ,n946);
    nand g2277(n1434 ,n715 ,n1059);
    nand g2278(n1740 ,n1009 ,n569);
    nand g2279(n1511 ,n1153 ,n612);
    nand g2280(n1187 ,n30[30] ,n351);
    nand g2281(n924 ,n4[4] ,n43);
    nor g2282(n1886 ,n21[31] ,n21[30]);
    not g2283(n42 ,n56);
    nand g2284(n923 ,n5[25] ,n349);
    nand g2285(n1314 ,n820 ,n499);
    nand g2286(n1078 ,n32[25] ,n46);
    nand g2287(n1752 ,n1008 ,n1737);
    nand g2288(n1094 ,n33[23] ,n355);
    nand g2289(n1171 ,n30[17] ,n54);
    nor g2290(n63 ,n21[21] ,n24[21]);
    nand g2291(n164 ,n28[14] ,n32[14]);
    nand g2292(n1673 ,n1239 ,n929);
    dff g2293(.RN(n1), .SN(1'b1), .CK(n0), .D(n1794), .Q(n31[8]));
    dff g2294(.RN(n1), .SN(1'b1), .CK(n0), .D(n1751), .Q(n13[6]));
    nand g2295(n1047 ,n26[12] ,n44);
    dff g2296(.RN(n1), .SN(1'b1), .CK(n0), .D(n1482), .Q(n23[1]));
    or g2297(n516 ,n287 ,n351);
    nand g2298(n637 ,n21[24] ,n347);
    dff g2299(.RN(n1), .SN(1'b1), .CK(n0), .D(n1628), .Q(n21[15]));
    nand g2300(n688 ,n11[23] ,n50);
    dff g2301(.RN(n1), .SN(1'b1), .CK(n0), .D(n1371), .Q(n32[24]));
    nand g2302(n970 ,n3[29] ,n349);
    nand g2303(n1360 ,n1014 ,n538);
    not g2304(n344 ,n346);
    dff g2305(.RN(n1), .SN(1'b1), .CK(n0), .D(n1700), .Q(n24[6]));
    nand g2306(n1576 ,n780 ,n1143);
    xnor g2307(n327 ,n22[7] ,n35[7]);
    dff g2308(.RN(n1), .SN(1'b1), .CK(n0), .D(n1375), .Q(n29[1]));
    nand g2309(n1574 ,n637 ,n810);
    nand g2310(n1166 ,n30[20] ,n54);
    nand g2311(n1925 ,n1918 ,n1908);
    nand g2312(n177 ,n28[2] ,n32[2]);
    nand g2313(n914 ,n5[31] ,n43);
    buf g2314(n16[9], n15[5]);
    nand g2315(n1554 ,n1170 ,n830);
    dff g2316(.RN(n1), .SN(1'b1), .CK(n0), .D(n1501), .Q(n28[10]));
    nor g2317(n107 ,n28[26] ,n32[26]);
    nand g2318(n1507 ,n1142 ,n610);
    dff g2319(.RN(n1), .SN(1'b1), .CK(n0), .D(n1559), .Q(n34[17]));
    nand g2320(n1636 ,n892 ,n1225);
    nand g2321(n1578 ,n834 ,n1169);
    nand g2322(n1597 ,n735 ,n1105);
    xnor g2323(n304 ,n21[4] ,n24[4]);
    nand g2324(n599 ,n21[17] ,n52);
    nand g2325(n742 ,n34[2] ,n352);
    nor g2326(n71 ,n31[15] ,n34[15]);
    nand g2327(n1487 ,n751 ,n1120);
    nand g2328(n1766 ,n1268 ,n1713);
    dff g2329(.RN(n1), .SN(1'b1), .CK(n0), .D(n1373), .Q(n29[3]));
    nand g2330(n1813 ,n1099 ,n1460);
    dff g2331(.RN(n1), .SN(1'b1), .CK(n0), .D(n1366), .Q(n32[31]));
    nand g2332(n185 ,n21[12] ,n24[12]);
    nand g2333(n848 ,n34[7] ,n352);
    nand g2334(n1309 ,n805 ,n459);
    nand g2335(n1546 ,n643 ,n855);
    buf g2336(n12[18], n11[18]);
    nand g2337(n1251 ,n29[31] ,n48);
    nand g2338(n800 ,n31[6] ,n352);
    nand g2339(n1898 ,n19[7] ,n19[6]);
    xnor g2340(n330 ,n22[3] ,n35[3]);
    dff g2341(.RN(n1), .SN(1'b1), .CK(n0), .D(n1770), .Q(n29[31]));
    nand g2342(n610 ,n21[6] ,n52);
    nand g2343(n1005 ,n15[8] ,n354);
    nor g2344(n115 ,n31[5] ,n34[5]);
    nand g2345(n1696 ,n1254 ,n949);
    dff g2346(.RN(n1), .SN(1'b1), .CK(n0), .D(n1789), .Q(n35[11]));
    nor g2347(n1903 ,n1895 ,n1893);
    nand g2348(n1194 ,n30[17] ,n351);
    nand g2349(n200 ,n29[12] ,n30[12]);
    nand g2350(n1780 ,n742 ,n1591);
    nand g2351(n182 ,n21[15] ,n24[15]);
    nand g2352(n1177 ,n30[13] ,n54);
    nand g2353(n1848 ,n149 ,n1846);
    nand g2354(n218 ,n29[5] ,n30[5]);
    nor g2355(n357 ,n155 ,n152);
    nand g2356(n1731 ,n996 ,n660);
    nand g2357(n1763 ,n1272 ,n1721);
    dff g2358(.RN(n1), .SN(1'b1), .CK(n0), .D(n1660), .Q(n22[7]));
    nand g2359(n902 ,n4[10] ,n43);
    dff g2360(.RN(n1), .SN(1'b1), .CK(n0), .D(n1825), .Q(n29[5]));
    nand g2361(n1412 ,n687 ,n562);
    nand g2362(n647 ,n21[14] ,n348);
    dff g2363(.RN(n1), .SN(1'b1), .CK(n0), .D(n1300), .Q(n35[30]));
    nand g2364(n1890 ,n24[25] ,n1863);
    nand g2365(n1227 ,n35[8] ,n45);
    nand g2366(n1244 ,n24[18] ,n348);
    nand g2367(n1470 ,n1111 ,n590);
    nand g2368(n1090 ,n32[17] ,n350);
    nand g2369(n928 ,n35[8] ,n356);
    dff g2370(.RN(n1), .SN(1'b1), .CK(n0), .D(n1570), .Q(n34[12]));
    dff g2371(.RN(n1), .SN(1'b1), .CK(n0), .D(n1377), .Q(n32[16]));
    nand g2372(n1806 ,n763 ,n1496);
    dff g2373(.RN(n1), .SN(1'b1), .CK(n0), .D(n1773), .Q(n33[1]));
    nand g2374(n1521 ,n727 ,n1147);
    nor g2375(n501 ,n114 ,n351);
    dff g2376(.RN(n1), .SN(1'b1), .CK(n0), .D(n1611), .Q(n33[24]));
    nand g2377(n1038 ,n26[19] ,n346);
    nand g2378(n1147 ,n33[11] ,n55);
    nand g2379(n556 ,n22[1] ,n348);
    dff g2380(.RN(n1), .SN(1'b1), .CK(n0), .D(n1321), .Q(n31[25]));
    nand g2381(n1198 ,n33[7] ,n55);
    or g2382(n383 ,n335 ,n48);
    nand g2383(n183 ,n21[14] ,n24[14]);
    nand g2384(n788 ,n35[23] ,n356);
    dff g2385(.RN(n1), .SN(1'b1), .CK(n0), .D(n1305), .Q(n35[22]));
    dff g2386(.RN(n1), .SN(1'b1), .CK(n0), .D(n1663), .Q(n22[6]));
    dff g2387(.RN(n1), .SN(1'b1), .CK(n0), .D(n1322), .Q(n31[24]));
    nor g2388(n1930 ,n1925 ,n1923);
    nand g2389(n1056 ,n26[6] ,n346);
    xnor g2390(n343 ,n26[6] ,n33[2]);
    nor g2391(n112 ,n28[27] ,n32[27]);
    nand g2392(n708 ,n11[9] ,n345);
    nand g2393(n665 ,n36[0] ,n56);
    nand g2394(n1263 ,n25[31] ,n51);
    nand g2395(n1293 ,n620 ,n411);
    nand g2396(n978 ,n35[29] ,n42);
    nand g2397(n1790 ,n802 ,n1526);
    nand g2398(n1803 ,n985 ,n1512);
    dff g2399(.RN(n1), .SN(1'b1), .CK(n0), .D(n1572), .Q(n30[23]));
    nand g2400(n1148 ,n28[3] ,n46);
    nand g2401(n1495 ,n1127 ,n602);
    nand g2402(n167 ,n29[8] ,n30[8]);
    nor g2403(n124 ,n28[31] ,n32[31]);
    dff g2404(.RN(n1), .SN(1'b1), .CK(n0), .D(n1648), .Q(n26[2]));
    nand g2405(n607 ,n21[9] ,n52);
    nor g2406(n96 ,n26[4] ,n33[0]);
    nand g2407(n971 ,n14[0] ,n50);
    nand g2408(n1582 ,n635 ,n790);
    dff g2409(.RN(n1), .SN(1'b1), .CK(n0), .D(n1365), .Q(n29[7]));
    nor g2410(n541 ,n142 ,n49);
    dff g2411(.RN(n1), .SN(1'b1), .CK(n0), .D(n1554), .Q(n30[28]));
    nand g2412(n772 ,n26[15] ,n354);
    nand g2413(n1036 ,n26[20] ,n45);
    or g2414(n527 ,n264 ,n356);
    nand g2415(n603 ,n21[13] ,n52);
    nand g2416(n741 ,n26[20] ,n354);
    nand g2417(n1095 ,n29[0] ,n47);
    nand g2418(n857 ,n32[17] ,n53);
    nor g2419(n450 ,n128 ,n42);
    nor g2420(n537 ,n145 ,n49);
    dff g2421(.RN(n1), .SN(1'b1), .CK(n0), .D(n1670), .Q(n24[24]));
    nand g2422(n1455 ,n182 ,n396);
    or g2423(n1841 ,n1286 ,n1767);
    nor g2424(n126 ,n31[1] ,n34[1]);
    nand g2425(n1175 ,n30[14] ,n54);
    nand g2426(n1201 ,n35[28] ,n45);
    nand g2427(n1682 ,n556 ,n934);
    nand g2428(n1255 ,n24[8] ,n51);
    dff g2429(.RN(n1), .SN(1'b1), .CK(n0), .D(n1293), .Q(n32[2]));
    dff g2430(.RN(n1), .SN(1'b1), .CK(n0), .D(n1311), .Q(n35[7]));
    nand g2431(n692 ,n11[20] ,n49);
    nand g2432(n614 ,n33[0] ,n49);
    nor g2433(n98 ,n28[14] ,n32[14]);
    nand g2434(n1482 ,n577 ,n746);
    nand g2435(n1425 ,n705 ,n1048);
    nand g2436(n1891 ,n21[25] ,n1859);
    nand g2437(n184 ,n21[13] ,n24[13]);
    nand g2438(n826 ,n34[24] ,n41);
    nand g2439(n1573 ,n641 ,n817);
    nand g2440(n1827 ,n1069 ,n1440);
    nand g2441(n577 ,n23[1] ,n348);
    dff g2442(.RN(n1), .SN(1'b1), .CK(n0), .D(n1550), .Q(n34[23]));
    buf g2443(n12[4], n11[4]);
    nand g2444(n1085 ,n33[25] ,n355);
    nand g2445(n633 ,n21[19] ,n348);
    nor g2446(n1889 ,n1855 ,n21[18]);
    nand g2447(n186 ,n21[11] ,n24[11]);
    nand g2448(n893 ,n26[2] ,n354);
    nand g2449(n953 ,n26[0] ,n354);
    nand g2450(n616 ,n32[6] ,n350);
    dff g2451(.RN(n1), .SN(1'b1), .CK(n0), .D(n1739), .Q(n15[8]));
    dff g2452(.RN(n1), .SN(1'b1), .CK(n0), .D(n1816), .Q(n29[0]));
    dff g2453(.RN(n1), .SN(1'b1), .CK(n0), .D(n1562), .Q(n34[16]));
    nor g2454(n92 ,n29[28] ,n30[28]);
    nand g2455(n1015 ,n13[4] ,n49);
    nand g2456(n612 ,n21[4] ,n52);
    dff g2457(.RN(n1), .SN(1'b1), .CK(n0), .D(n1415), .Q(n11[19]));
endmodule
