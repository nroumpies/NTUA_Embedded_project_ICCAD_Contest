module top (n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [2:0] n6;
    wire [15:0] n7;
    wire [7:0] n8;
    wire n9, n10, n11, n12, n13, n14, n15, n16;
    wire n17, n18, n19, n20, n21, n22, n23, n24;
    wire n25, n26, n27, n28, n29, n30, n31, n32;
    wire n33, n34, n35, n36, n37, n38, n39, n40;
    wire n41, n42, n43, n44, n45, n46, n47, n48;
    wire n49, n50, n51, n52, n53, n54, n55, n56;
    wire n57, n58, n59, n60, n61, n62, n63, n64;
    wire n65, n66, n67, n68, n69, n70, n71, n72;
    wire n73, n74, n75, n76, n77, n78, n79, n80;
    wire n81, n82, n83, n84, n85, n86, n87, n88;
    wire n89, n90, n91, n92, n93, n94, n95, n96;
    wire n97, n98, n99, n100, n101, n102, n103, n104;
    wire n105, n106, n107, n108, n109, n110, n111, n112;
    wire n113, n114, n115, n116, n117, n118, n119, n120;
    wire n121, n122, n123, n124, n125, n126, n127, n128;
    wire n129, n130, n131, n132, n133, n134, n135, n136;
    wire n137, n138, n139, n140, n141, n142, n143, n144;
    wire n145, n146, n147, n148, n149, n150, n151, n152;
    wire n153, n154, n155, n156, n157, n158, n159, n160;
    wire n161, n162, n163, n164, n165, n166, n167, n168;
    wire n169, n170, n171, n172, n173, n174, n175, n176;
    wire n177, n178, n179, n180, n181, n182, n183, n184;
    wire n185, n186, n187, n188, n189, n190, n191, n192;
    wire n193, n194, n195, n196, n197, n198, n199, n200;
    wire n201, n202, n203, n204, n205, n206, n207, n208;
    wire n209, n210, n211, n212, n213, n214, n215, n216;
    wire n217, n218, n219, n220, n221, n222, n223, n224;
    wire n225, n226, n227, n228, n229, n230, n231, n232;
    wire n233, n234, n235, n236, n237, n238, n239, n240;
    wire n241, n242, n243, n244, n245, n246, n247, n248;
    wire n249, n250, n251, n252, n253, n254, n255, n256;
    wire n257, n258, n259, n260, n261, n262, n263, n264;
    wire n265, n266, n267, n268, n269, n270, n271, n272;
    wire n273, n274, n275, n276, n277, n278, n279, n280;
    wire n281, n282, n283, n284, n285, n286, n287, n288;
    wire n289, n290, n291, n292, n293, n294, n295, n296;
    wire n297, n298, n299, n300, n301, n302, n303, n304;
    wire n305, n306, n307, n308, n309, n310, n311, n312;
    wire n313, n314, n315, n316, n317, n318, n319, n320;
    wire n321, n322, n323, n324, n325, n326, n327, n328;
    wire n329, n330, n331, n332, n333, n334, n335, n336;
    wire n337, n338, n339, n340, n341, n342, n343, n344;
    wire n345, n346, n347, n348, n349, n350, n351, n352;
    wire n353, n354, n355, n356, n357, n358, n359, n360;
    wire n361, n362, n363, n364, n365, n366, n367, n368;
    wire n369, n370, n371, n372, n373, n374, n375, n376;
    wire n377, n378, n379, n380, n381, n382, n383, n384;
    wire n385, n386, n387, n388, n389, n390, n391, n392;
    wire n393, n394, n395, n396, n397, n398, n399, n400;
    wire n401, n402, n403, n404, n405, n406, n407, n408;
    wire n409, n410, n411, n412, n413, n414, n415, n416;
    wire n417, n418, n419, n420, n421, n422, n423, n424;
    wire n425, n426, n427, n428, n429, n430, n431, n432;
    wire n433, n434, n435, n436, n437, n438, n439, n440;
    wire n441, n442, n443, n444, n445, n446, n447, n448;
    wire n449, n450, n451, n452, n453, n454, n455, n456;
    wire n457, n458, n459, n460, n461, n462, n463, n464;
    wire n465, n466, n467, n468, n469, n470, n471, n472;
    wire n473, n474, n475, n476, n477, n478, n479, n480;
    wire n481, n482, n483, n484, n485, n486, n487, n488;
    wire n489, n490, n491, n492, n493, n494, n495, n496;
    wire n497, n498, n499, n500, n501, n502, n503, n504;
    wire n505, n506, n507, n508, n509, n510, n511, n512;
    wire n513, n514, n515, n516, n517, n518, n519, n520;
    wire n521, n522, n523, n524, n525, n526, n527, n528;
    wire n529, n530, n531, n532, n533, n534, n535, n536;
    wire n537, n538, n539, n540, n541, n542, n543, n544;
    wire n545, n546, n547, n548, n549, n550, n551, n552;
    wire n553, n554, n555, n556, n557, n558, n559, n560;
    wire n561, n562, n563, n564, n565, n566, n567, n568;
    wire n569, n570, n571, n572, n573, n574, n575, n576;
    wire n577, n578, n579, n580, n581, n582, n583, n584;
    wire n585, n586, n587, n588, n589, n590, n591, n592;
    wire n593, n594, n595, n596, n597, n598, n599, n600;
    wire n601, n602, n603, n604, n605, n606, n607, n608;
    wire n609, n610, n611, n612, n613, n614, n615, n616;
    wire n617, n618, n619, n620, n621, n622, n623, n624;
    wire n625, n626, n627, n628, n629, n630, n631, n632;
    wire n633, n634, n635, n636, n637, n638, n639, n640;
    wire n641, n642, n643, n644, n645, n646, n647, n648;
    wire n649, n650, n651, n652, n653, n654, n655, n656;
    wire n657, n658, n659, n660, n661, n662, n663, n664;
    wire n665, n666, n667, n668, n669, n670, n671, n672;
    wire n673, n674, n675, n676, n677, n678, n679, n680;
    wire n681, n682, n683, n684, n685, n686, n687, n688;
    wire n689, n690, n691, n692, n693, n694, n695, n696;
    wire n697, n698, n699, n700, n701, n702, n703, n704;
    wire n705, n706, n707, n708, n709, n710, n711, n712;
    wire n713, n714, n715, n716, n717, n718, n719, n720;
    wire n721, n722, n723, n724, n725, n726, n727, n728;
    wire n729, n730, n731, n732, n733, n734, n735, n736;
    wire n737, n738, n739, n740, n741, n742, n743, n744;
    wire n745, n746, n747, n748, n749, n750, n751, n752;
    wire n753, n754, n755, n756, n757, n758, n759, n760;
    wire n761, n762, n763, n764, n765, n766, n767, n768;
    wire n769, n770, n771, n772, n773, n774, n775, n776;
    wire n777, n778, n779, n780, n781, n782, n783, n784;
    wire n785, n786, n787, n788, n789, n790, n791, n792;
    wire n793, n794, n795, n796, n797, n798, n799, n800;
    wire n801, n802, n803, n804, n805, n806, n807, n808;
    wire n809, n810, n811, n812, n813, n814, n815, n816;
    wire n817, n818, n819, n820, n821, n822, n823, n824;
    wire n825, n826, n827, n828, n829, n830, n831, n832;
    wire n833, n834, n835, n836, n837, n838, n839, n840;
    wire n841, n842, n843, n844, n845, n846, n847, n848;
    wire n849, n850, n851, n852, n853, n854, n855, n856;
    wire n857, n858, n859, n860, n861, n862, n863, n864;
    wire n865, n866, n867, n868, n869, n870, n871, n872;
    wire n873, n874, n875, n876, n877, n878, n879, n880;
    wire n881, n882, n883, n884, n885, n886, n887, n888;
    wire n889, n890, n891, n892, n893, n894, n895, n896;
    wire n897, n898, n899, n900, n901, n902, n903, n904;
    wire n905, n906, n907, n908, n909, n910, n911, n912;
    wire n913, n914, n915, n916, n917, n918, n919, n920;
    wire n921, n922, n923, n924, n925, n926, n927, n928;
    wire n929, n930, n931, n932, n933, n934, n935, n936;
    wire n937, n938, n939, n940, n941, n942, n943, n944;
    wire n945, n946, n947, n948, n949, n950, n951, n952;
    wire n953, n954, n955, n956, n957, n958, n959, n960;
    wire n961, n962, n963, n964, n965, n966, n967, n968;
    wire n969, n970, n971, n972, n973, n974, n975, n976;
    wire n977, n978, n979, n980, n981, n982, n983, n984;
    wire n985, n986, n987, n988, n989, n990, n991, n992;
    wire n993, n994, n995, n996, n997, n998, n999, n1000;
    wire n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008;
    wire n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016;
    wire n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
    wire n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
    wire n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040;
    wire n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
    wire n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056;
    wire n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064;
    wire n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072;
    wire n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080;
    wire n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088;
    wire n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096;
    wire n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104;
    wire n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112;
    wire n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120;
    wire n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128;
    wire n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136;
    wire n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144;
    wire n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152;
    wire n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160;
    wire n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168;
    wire n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176;
    wire n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184;
    wire n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192;
    wire n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200;
    wire n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208;
    wire n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216;
    wire n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224;
    wire n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232;
    wire n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240;
    wire n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248;
    wire n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256;
    wire n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264;
    wire n1265, n1266, n1267, n1268;
    nand g0(n368 ,n6[1] ,n362);
    dff g1(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n999), .Q(n3[6]));
    xnor g2(n1265 ,n8[4] ,n1199);
    dff g3(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n930), .Q(n4[51]));
    nand g4(n606 ,n3[19] ,n353);
    nor g5(n480 ,n1 ,n354);
    nand g6(n1223 ,n1 ,n2[15]);
    xnor g7(n1150 ,n3[49] ,n153);
    nand g8(n811 ,n7[15] ,n648);
    nand g9(n97 ,n3[16] ,n95);
    nand g10(n835 ,n3[11] ,n639);
    nand g11(n993 ,n791 ,n945);
    nand g12(n733 ,n491 ,n669);
    nand g13(n526 ,n1136 ,n378);
    not g14(n950 ,n904);
    nand g15(n787 ,n7[4] ,n621);
    nand g16(n700 ,n583 ,n518);
    nand g17(n1236 ,n1 ,n2[1]);
    nand g18(n207 ,n7[6] ,n182);
    not g19(n943 ,n897);
    nand g20(n201 ,n7[15] ,n188);
    nand g21(n749 ,n4[41] ,n351);
    xnor g22(n221 ,n4[3] ,n7[3]);
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1003), .Q(n3[10]));
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n704), .Q(n3[39]));
    nand g25(n470 ,n1078 ,n379);
    dff g26(.RN(n1208), .SN(n1224), .CK(n0), .D(n1248), .Q(n7[14]));
    nand g27(n437 ,n1052 ,n379);
    nand g28(n885 ,n464 ,n777);
    nor g29(n806 ,n361 ,n641);
    xnor g30(n60 ,n7[10] ,n3[10]);
    nand g31(n1224 ,n1 ,n2[14]);
    xor g32(n1025 ,n617 ,n975);
    not g33(n1196 ,n1195);
    xor g34(n1022 ,n614 ,n978);
    or g35(n492 ,n7[5] ,n374);
    or g36(n1001 ,n778 ,n869);
    nand g37(n447 ,n1103 ,n355);
    buf g38(n5[61], 1'b0);
    or g39(n658 ,n476 ,n412);
    nand g40(n542 ,n1122 ,n379);
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n924), .Q(n4[56]));
    nor g42(n109 ,n17 ,n108);
    nand g43(n867 ,n555 ,n759);
    nand g44(n248 ,n197 ,n247);
    nand g45(n1010 ,n459 ,n855);
    nand g46(n558 ,n1091 ,n379);
    not g47(n105 ,n104);
    nand g48(n604 ,n3[21] ,n376);
    nand g49(n760 ,n4[33] ,n668);
    nand g50(n742 ,n486 ,n669);
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n937), .Q(n4[45]));
    nor g52(n151 ,n12 ,n150);
    nand g53(n681 ,n566 ,n498);
    nand g54(n234 ,n206 ,n233);
    xor g55(n1021 ,n615 ,n979);
    nand g56(n277 ,n4[26] ,n274);
    or g57(n21 ,n3[13] ,n7[13]);
    xnor g58(n1052 ,n215 ,n254);
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n715), .Q(n3[28]));
    xnor g60(n1045 ,n224 ,n240);
    nand g61(n1015 ,n533 ,n1014);
    dff g62(.RN(n1218), .SN(n1234), .CK(n0), .D(n1258), .Q(n7[4]));
    nand g63(n245 ,n213 ,n244);
    nand g64(n841 ,n7[0] ,n670);
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1035), .Q(n5[5]));
    nand g66(n679 ,n7[9] ,n478);
    xnor g67(n1254 ,n2[8] ,n1180);
    not g68(n478 ,n477);
    nand g69(n335 ,n4[55] ,n332);
    xnor g70(n59 ,n7[2] ,n3[2]);
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1006), .Q(n3[13]));
    nand g72(n78 ,n35 ,n77);
    nor g73(n391 ,n4[13] ,n374);
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1001), .Q(n3[8]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n705), .Q(n3[38]));
    not g76(n942 ,n896);
    nand g77(n977 ,n5[12] ,n890);
    not g78(n135 ,n134);
    buf g79(n5[35], 1'b0);
    nor g80(n397 ,n4[15] ,n374);
    or g81(n270 ,n4[23] ,n268);
    nand g82(n600 ,n3[25] ,n376);
    nand g83(n1187 ,n2[11] ,n1186);
    xnor g84(n1123 ,n3[22] ,n106);
    dff g85(.RN(n1219), .SN(n1235), .CK(n0), .D(n1259), .Q(n7[3]));
    nor g86(n406 ,n3[14] ,n374);
    nand g87(n1018 ,n841 ,n1013);
    dff g88(.RN(n1205), .SN(1'b1), .CK(n0), .D(n1263), .Q(n8[6]));
    nand g89(n1054 ,n259 ,n258);
    nand g90(n530 ,n1132 ,n379);
    nand g91(n775 ,n7[5] ,n662);
    nand g92(n736 ,n489 ,n669);
    or g93(n1209 ,n1205 ,n2[13]);
    buf g94(n5[53], 1'b0);
    nand g95(n279 ,n4[27] ,n276);
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1008), .Q(n3[12]));
    xnor g97(n1122 ,n3[21] ,n104);
    nand g98(n509 ,n1093 ,n379);
    or g99(n276 ,n4[26] ,n274);
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n939), .Q(n4[43]));
    nand g101(n1074 ,n299 ,n298);
    nand g102(n735 ,n487 ,n669);
    not g103(n369 ,n370);
    nand g104(n872 ,n417 ,n765);
    nand g105(n1063 ,n277 ,n276);
    nand g106(n90 ,n21 ,n89);
    or g107(n260 ,n4[18] ,n258);
    nand g108(n773 ,n4[23] ,n668);
    nand g109(n473 ,n1079 ,n354);
    nand g110(n305 ,n4[40] ,n302);
    or g111(n1210 ,n1205 ,n2[11]);
    nand g112(n256 ,n201 ,n255);
    nand g113(n753 ,n7[9] ,n638);
    xnor g114(n1112 ,n61 ,n85);
    not g115(n142 ,n141);
    nand g116(n724 ,n606 ,n544);
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n929), .Q(n4[52]));
    buf g118(n5[40], 1'b0);
    not g119(n358 ,n1);
    nor g120(n392 ,n4[1] ,n374);
    nand g121(n594 ,n3[31] ,n353);
    nand g122(n267 ,n4[21] ,n264);
    nand g123(n566 ,n3[62] ,n376);
    or g124(n1207 ,n1205 ,n2[12]);
    nand g125(n720 ,n602 ,n540);
    xor g126(n1020 ,n616 ,n965);
    nand g127(n1095 ,n341 ,n340);
    nand g128(n708 ,n590 ,n526);
    nand g129(n869 ,n552 ,n756);
    nand g130(n1243 ,n8[7] ,n1242);
    not g131(n107 ,n106);
    nand g132(n698 ,n565 ,n516);
    nand g133(n649 ,n485 ,n479);
    nor g134(n363 ,n6[0] ,n6[1]);
    nor g135(n1189 ,n2[13] ,n1188);
    or g136(n485 ,n7[15] ,n374);
    nor g137(n412 ,n3[10] ,n374);
    nand g138(n515 ,n1100 ,n355);
    nand g139(n868 ,n431 ,n760);
    nand g140(n427 ,n1149 ,n356);
    not g141(n13 ,n3[27]);
    nand g142(n809 ,n3[7] ,n665);
    xnor g143(n1126 ,n3[25] ,n111);
    nand g144(n582 ,n3[44] ,n353);
    nand g145(n647 ,n495 ,n479);
    nand g146(n865 ,n556 ,n757);
    nand g147(n675 ,n7[4] ,n478);
    xor g148(n1024 ,n618 ,n976);
    or g149(n1219 ,n1205 ,n2[3]);
    buf g150(n5[20], 1'b0);
    nand g151(n840 ,n3[10] ,n656);
    buf g152(n5[49], 1'b0);
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n725), .Q(n3[18]));
    nand g154(n42 ,n3[8] ,n7[8]);
    nand g155(n231 ,n221 ,n230);
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n994), .Q(n4[13]));
    nand g157(n233 ,n226 ,n232);
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1020), .Q(n5[15]));
    nor g159(n1175 ,n2[5] ,n1174);
    buf g160(n5[52], 1'b0);
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1000), .Q(n3[7]));
    nand g162(n469 ,n1038 ,n379);
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n983), .Q(n4[6]));
    nand g164(n518 ,n1144 ,n354);
    nand g165(n275 ,n4[25] ,n272);
    not g166(n352 ,n376);
    nand g167(n510 ,n1151 ,n355);
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1025), .Q(n5[10]));
    not g169(n895 ,n889);
    nand g170(n827 ,n4[53] ,n351);
    xnor g171(n1139 ,n3[38] ,n134);
    nor g172(n1200 ,n1193 ,n1199);
    nand g173(n293 ,n4[34] ,n290);
    nand g174(n726 ,n608 ,n546);
    nand g175(n1204 ,n8[6] ,n1203);
    nand g176(n499 ,n1162 ,n356);
    nand g177(n111 ,n3[24] ,n109);
    nor g178(n1182 ,n2[9] ,n1181);
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n996), .Q(n3[4]));
    nand g180(n911 ,n469 ,n808);
    nand g181(n932 ,n434 ,n831);
    nand g182(n164 ,n3[54] ,n163);
    nor g183(n381 ,n4[6] ,n374);
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n925), .Q(n4[55]));
    xor g185(n1102 ,n57 ,n50);
    nand g186(n1227 ,n1 ,n2[11]);
    nand g187(n730 ,n494 ,n669);
    nand g188(n434 ,n1086 ,n378);
    nand g189(n738 ,n492 ,n669);
    not g190(n1013 ,n1012);
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1027), .Q(n5[8]));
    nand g192(n761 ,n4[32] ,n351);
    nand g193(n986 ,n849 ,n951);
    nand g194(n101 ,n3[18] ,n100);
    nand g195(n972 ,n5[7] ,n890);
    nand g196(n725 ,n607 ,n545);
    nand g197(n93 ,n41 ,n92);
    nand g198(n938 ,n416 ,n838);
    nand g199(n1075 ,n301 ,n300);
    or g200(n1215 ,n1205 ,n2[6]);
    nand g201(n1060 ,n271 ,n270);
    nand g202(n870 ,n563 ,n761);
    or g203(n637 ,n380 ,n402);
    nand g204(n204 ,n7[2] ,n193);
    dff g205(.RN(n1222), .SN(n1237), .CK(n0), .D(n2[0]), .Q(n7[0]));
    not g206(n1193 ,n8[4]);
    nand g207(n301 ,n4[38] ,n298);
    nand g208(n804 ,n3[0] ,n636);
    nand g209(n750 ,n4[40] ,n668);
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n877), .Q(n4[26]));
    nand g211(n984 ,n853 ,n955);
    nand g212(n307 ,n4[41] ,n304);
    or g213(n619 ,n380 ,n397);
    nor g214(n1149 ,n152 ,n154);
    xnor g215(n64 ,n7[14] ,n3[14]);
    xnor g216(n1039 ,n220 ,n228);
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n721), .Q(n3[22]));
    dff g218(.RN(n1205), .SN(1'b1), .CK(n0), .D(n1262), .Q(n8[7]));
    nand g219(n919 ,n456 ,n818);
    xnor g220(n1048 ,n212 ,n246);
    or g221(n324 ,n4[50] ,n322);
    nand g222(n129 ,n3[34] ,n128);
    xnor g223(n1251 ,n2[11] ,n1185);
    nand g224(n246 ,n205 ,n245);
    nand g225(n1171 ,n2[2] ,n1170);
    nor g226(n376 ,n1 ,n363);
    buf g227(n5[54], 1'b0);
    nor g228(n1264 ,n1201 ,n1203);
    nand g229(n496 ,n359 ,n375);
    nand g230(n609 ,n3[16] ,n376);
    not g231(n954 ,n908);
    nand g232(n674 ,n7[5] ,n478);
    nand g233(n624 ,n496 ,n479);
    nand g234(n940 ,n832 ,n840);
    nand g235(n774 ,n3[6] ,n663);
    nand g236(n896 ,n437 ,n784);
    not g237(n187 ,n7[0]);
    xnor g238(n62 ,n7[12] ,n3[12]);
    not g239(n374 ,n375);
    nand g240(n1097 ,n345 ,n344);
    xnor g241(n1163 ,n3[62] ,n176);
    nand g242(n416 ,n1081 ,n356);
    nand g243(n47 ,n3[10] ,n7[10]);
    nand g244(n1086 ,n323 ,n322);
    nand g245(n684 ,n568 ,n501);
    nand g246(n487 ,n360 ,n375);
    not g247(n952 ,n906);
    dff g248(.RN(n1205), .SN(1'b1), .CK(n0), .D(n1267), .Q(n8[2]));
    nand g249(n327 ,n4[51] ,n324);
    nand g250(n441 ,n1104 ,n379);
    nand g251(n917 ,n475 ,n815);
    nor g252(n158 ,n19 ,n157);
    xnor g253(n1140 ,n3[39] ,n136);
    buf g254(n5[60], 1'b0);
    nand g255(n783 ,n4[16] ,n668);
    nor g256(n124 ,n3[32] ,n123);
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n698), .Q(n3[45]));
    nand g258(n562 ,n1049 ,n356);
    nand g259(n36 ,n3[7] ,n7[7]);
    nand g260(n906 ,n451 ,n798);
    or g261(n28 ,n3[5] ,n7[5]);
    nand g262(n169 ,n3[57] ,n168);
    nand g263(n540 ,n1124 ,n378);
    or g264(n640 ,n476 ,n396);
    nand g265(n1180 ,n2[7] ,n1179);
    or g266(n280 ,n4[28] ,n278);
    or g267(n25 ,n3[2] ,n7[2]);
    xor g268(n1099 ,n4[62] ,n346);
    or g269(n316 ,n4[46] ,n314);
    nand g270(n448 ,n1088 ,n379);
    buf g271(n5[38], 1'b0);
    xnor g272(n1113 ,n62 ,n87);
    or g273(n300 ,n4[38] ,n298);
    nand g274(n82 ,n29 ,n81);
    xor g275(n1027 ,n671 ,n973);
    nor g276(n131 ,n3[36] ,n130);
    nor g277(n166 ,n3[56] ,n165);
    nand g278(n757 ,n4[36] ,n668);
    dff g279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n926), .Q(n4[54]));
    nand g280(n623 ,n488 ,n479);
    nor g281(n410 ,n3[9] ,n374);
    nor g282(n1133 ,n124 ,n126);
    or g283(n1216 ,n1205 ,n2[7]);
    nand g284(n46 ,n3[9] ,n7[9]);
    nand g285(n712 ,n594 ,n530);
    nand g286(n727 ,n609 ,n548);
    nand g287(n1081 ,n313 ,n312);
    not g288(n182 ,n4[6]);
    nand g289(n423 ,n1068 ,n355);
    nand g290(n777 ,n4[20] ,n351);
    nand g291(n907 ,n453 ,n799);
    nand g292(n884 ,n432 ,n775);
    nand g293(n197 ,n7[11] ,n191);
    nand g294(n1077 ,n305 ,n304);
    nand g295(n978 ,n5[13] ,n890);
    or g296(n1217 ,n1205 ,n2[5]);
    xnor g297(n1115 ,n64 ,n91);
    nand g298(n980 ,n801 ,n950);
    or g299(n482 ,n7[9] ,n374);
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n695), .Q(n3[48]));
    nand g301(n1089 ,n329 ,n328);
    or g302(n1214 ,n1205 ,n2[15]);
    dff g303(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1024), .Q(n5[11]));
    nand g304(n731 ,n495 ,n669);
    nand g305(n581 ,n3[46] ,n353);
    nand g306(n139 ,n3[40] ,n137);
    nand g307(n321 ,n4[48] ,n318);
    not g308(n894 ,n884);
    xnor g309(n1124 ,n3[23] ,n108);
    buf g310(n5[57], 1'b0);
    buf g311(n5[29], 1'b0);
    xor g312(n1031 ,n678 ,n966);
    dff g313(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1028), .Q(n5[7]));
    xnor g314(n1136 ,n3[35] ,n129);
    nand g315(n825 ,n3[12] ,n647);
    nand g316(n560 ,n1113 ,n378);
    nand g317(n596 ,n3[29] ,n353);
    nand g318(n457 ,n1042 ,n356);
    xnor g319(n1040 ,n221 ,n230);
    xnor g320(n1044 ,n217 ,n238);
    dff g321(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n875), .Q(n4[28]));
    or g322(n322 ,n4[49] ,n320);
    nand g323(n923 ,n508 ,n822);
    xnor g324(n1043 ,n225 ,n236);
    dff g325(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n709), .Q(n3[34]));
    nand g326(n616 ,n7[15] ,n478);
    not g327(n140 ,n139);
    or g328(n629 ,n476 ,n400);
    dff g329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n870), .Q(n4[32]));
    xnor g330(n218 ,n4[13] ,n7[13]);
    nand g331(n677 ,n7[2] ,n478);
    nor g332(n401 ,n4[12] ,n374);
    nand g333(n43 ,n3[15] ,n7[15]);
    dff g334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n690), .Q(n3[53]));
    nand g335(n1084 ,n319 ,n318);
    dff g336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n989), .Q(n4[10]));
    nand g337(n873 ,n421 ,n763);
    nand g338(n452 ,n1092 ,n356);
    nand g339(n1008 ,n560 ,n962);
    dff g340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n713), .Q(n3[30]));
    nand g341(n740 ,n488 ,n669);
    dff g342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n993), .Q(n3[3]));
    nand g343(n789 ,n7[3] ,n653);
    nand g344(n585 ,n3[40] ,n353);
    nand g345(n859 ,n463 ,n753);
    nor g346(n373 ,n6[2] ,n371);
    dff g347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n991), .Q(n4[0]));
    not g348(n361 ,n7[3]);
    nand g349(n1169 ,n2[1] ,n1246);
    nand g350(n843 ,n4[15] ,n728);
    nand g351(n257 ,n185 ,n256);
    nand g352(n987 ,n795 ,n949);
    nand g353(n784 ,n7[15] ,n619);
    nand g354(n535 ,n1129 ,n354);
    nand g355(n769 ,n4[26] ,n351);
    nand g356(n593 ,n3[32] ,n376);
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n916), .Q(n4[63]));
    nand g358(n370 ,n6[0] ,n362);
    nand g359(n590 ,n3[35] ,n376);
    xnor g360(n1256 ,n2[6] ,n1176);
    nand g361(n595 ,n3[30] ,n353);
    nand g362(n235 ,n223 ,n234);
    nand g363(n836 ,n4[46] ,n668);
    nand g364(n813 ,n7[14] ,n650);
    nand g365(n575 ,n3[52] ,n353);
    nand g366(n822 ,n4[57] ,n351);
    buf g367(n5[32], 1'b0);
    or g368(n634 ,n476 ,n411);
    nand g369(n925 ,n452 ,n824);
    xnor g370(n1247 ,n2[15] ,n1192);
    buf g371(n5[30], 1'b0);
    nand g372(n810 ,n4[22] ,n668);
    nand g373(n1230 ,n1 ,n2[8]);
    not g374(n949 ,n903);
    nand g375(n1241 ,n8[6] ,n8[5]);
    nand g376(n979 ,n5[14] ,n890);
    nand g377(n743 ,n497 ,n669);
    nand g378(n1005 ,n826 ,n960);
    or g379(n272 ,n4[24] ,n270);
    not g380(n1179 ,n1178);
    nor g381(n1194 ,n8[1] ,n8[0]);
    nand g382(n992 ,n846 ,n946);
    buf g383(n5[16], 1'b0);
    or g384(n644 ,n380 ,n386);
    nand g385(n693 ,n577 ,n510);
    nand g386(n254 ,n202 ,n253);
    nand g387(n759 ,n4[34] ,n351);
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1021), .Q(n5[14]));
    xnor g389(n61 ,n7[11] ,n3[11]);
    xor g390(n1028 ,n672 ,n972);
    xnor g391(n212 ,n4[11] ,n7[11]);
    dff g392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n724), .Q(n3[19]));
    nand g393(n831 ,n4[49] ,n351);
    not g394(n133 ,n132);
    nand g395(n463 ,n1110 ,n378);
    nand g396(n337 ,n4[56] ,n334);
    nand g397(n578 ,n3[49] ,n353);
    dff g398(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n998), .Q(n3[5]));
    xnor g399(n1252 ,n2[10] ,n1183);
    not g400(n1172 ,n1171);
    nor g401(n349 ,n4[62] ,n347);
    nand g402(n440 ,n1064 ,n379);
    xnor g403(n1266 ,n8[3] ,n1197);
    nand g404(n808 ,n7[1] ,n643);
    not g405(n1165 ,n2[4]);
    nand g406(n89 ,n37 ,n88);
    nand g407(n883 ,n461 ,n776);
    nand g408(n73 ,n38 ,n72);
    nand g409(n281 ,n4[28] ,n278);
    dff g410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n997), .Q(n4[15]));
    xnor g411(n1144 ,n3[43] ,n143);
    nand g412(n531 ,n1062 ,n378);
    nand g413(n325 ,n4[50] ,n322);
    nand g414(n793 ,n7[2] ,n627);
    not g415(n963 ,n934);
    nand g416(n418 ,n1066 ,n355);
    nand g417(n936 ,n564 ,n836);
    nand g418(n249 ,n222 ,n248);
    nand g419(n886 ,n433 ,n779);
    not g420(n195 ,n4[10]);
    nand g421(n436 ,n1054 ,n379);
    nand g422(n617 ,n7[10] ,n478);
    nand g423(n814 ,n4[63] ,n351);
    or g424(n643 ,n380 ,n392);
    nand g425(n1185 ,n2[10] ,n1184);
    nand g426(n435 ,n1152 ,n356);
    nand g427(n532 ,n1131 ,n378);
    nand g428(n844 ,n4[14] ,n729);
    nand g429(n539 ,n1125 ,n378);
    xnor g430(n1134 ,n3[33] ,n125);
    nand g431(n456 ,n1097 ,n355);
    nand g432(n323 ,n4[49] ,n320);
    nand g433(n141 ,n3[41] ,n140);
    dff g434(.RN(n1205), .SN(1'b1), .CK(n0), .D(n1266), .Q(n8[3]));
    or g435(n336 ,n4[56] ,n334);
    or g436(n334 ,n4[55] ,n332);
    nand g437(n1072 ,n295 ,n294);
    not g438(n10 ,n3[59]);
    xnor g439(n1128 ,n3[27] ,n115);
    xnor g440(n1042 ,n223 ,n234);
    nand g441(n689 ,n573 ,n506);
    nand g442(n888 ,n436 ,n781);
    nand g443(n817 ,n7[13] ,n645);
    nand g444(n475 ,n1099 ,n355);
    buf g445(n5[28], 1'b0);
    not g446(n19 ,n3[51]);
    not g447(n119 ,n118);
    nand g448(n438 ,n1105 ,n378);
    xnor g449(n224 ,n4[8] ,n7[8]);
    dff g450(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n922), .Q(n4[58]));
    xnor g451(n1108 ,n56 ,n77);
    nand g452(n345 ,n4[60] ,n342);
    nand g453(n707 ,n589 ,n525);
    nand g454(n104 ,n3[20] ,n102);
    nand g455(n80 ,n34 ,n79);
    xor g456(n1030 ,n676 ,n968);
    nor g457(n173 ,n3[60] ,n172);
    not g458(n170 ,n169);
    xor g459(n1037 ,n7[0] ,n4[0]);
    xnor g460(n54 ,n7[5] ,n3[5]);
    nand g461(n250 ,n196 ,n249);
    or g462(n650 ,n476 ,n406);
    nand g463(n569 ,n3[58] ,n353);
    dff g464(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1031), .Q(n5[1]));
    not g465(n951 ,n905);
    xnor g466(n1107 ,n55 ,n75);
    nand g467(n751 ,n7[12] ,n657);
    nand g468(n148 ,n3[45] ,n147);
    nand g469(n1085 ,n321 ,n320);
    nand g470(n563 ,n1069 ,n379);
    nand g471(n1003 ,n474 ,n964);
    xnor g472(n1120 ,n3[19] ,n101);
    nand g473(n127 ,n3[33] ,n126);
    nand g474(n1233 ,n1 ,n2[5]);
    or g475(n497 ,n7[0] ,n374);
    nand g476(n755 ,n4[37] ,n351);
    nand g477(n211 ,n7[5] ,n180);
    nand g478(n460 ,n1077 ,n379);
    nand g479(n765 ,n7[7] ,n666);
    xnor g480(n1114 ,n63 ,n89);
    nand g481(n695 ,n579 ,n427);
    dff g482(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n866), .Q(n4[35]));
    nand g483(n415 ,n1065 ,n356);
    nor g484(n405 ,n3[7] ,n374);
    xor g485(n1033 ,n677 ,n967);
    not g486(n180 ,n4[5]);
    or g487(n34 ,n3[8] ,n7[8]);
    or g488(n310 ,n4[43] ,n308);
    nand g489(n1202 ,n8[5] ,n1200);
    nand g490(n752 ,n4[39] ,n668);
    dff g491(.RN(n1216), .SN(n1231), .CK(n0), .D(n1255), .Q(n7[7]));
    dff g492(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1016), .Q(n4[3]));
    not g493(n1206 ,n8[0]);
    not g494(n946 ,n900);
    nand g495(n613 ,n7[12] ,n478);
    dff g496(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n868), .Q(n4[33]));
    nand g497(n511 ,n1150 ,n356);
    dff g498(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n744), .Q(n6[0]));
    nand g499(n253 ,n216 ,n252);
    nand g500(n792 ,n7[11] ,n625);
    not g501(n163 ,n162);
    nand g502(n243 ,n214 ,n242);
    dff g503(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n702), .Q(n3[41]));
    nand g504(n255 ,n215 ,n254);
    nor g505(n144 ,n15 ,n143);
    nand g506(n1093 ,n337 ,n336);
    nand g507(n573 ,n3[54] ,n353);
    nand g508(n1082 ,n315 ,n314);
    nand g509(n796 ,n7[9] ,n628);
    dff g510(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n931), .Q(n4[50]));
    nand g511(n206 ,n7[4] ,n192);
    nand g512(n580 ,n3[47] ,n353);
    dff g513(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n719), .Q(n3[24]));
    not g514(n191 ,n4[11]);
    nand g515(n914 ,n549 ,n811);
    nand g516(n297 ,n4[36] ,n294);
    nand g517(n1228 ,n1 ,n2[10]);
    dff g518(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n874), .Q(n4[29]));
    nand g519(n599 ,n3[26] ,n376);
    nand g520(n786 ,n7[14] ,n620);
    nand g521(n968 ,n5[3] ,n890);
    nand g522(n564 ,n1083 ,n378);
    or g523(n491 ,n7[10] ,n374);
    nand g524(n471 ,n1037 ,n379);
    buf g525(n5[36], 1'b0);
    nand g526(n795 ,n3[2] ,n624);
    nand g527(n242 ,n210 ,n241);
    nand g528(n238 ,n207 ,n237);
    or g529(n318 ,n4[47] ,n316);
    nand g530(n864 ,n559 ,n755);
    or g531(n1222 ,n1205 ,n2[0]);
    nand g532(n903 ,n447 ,n793);
    nand g533(n505 ,n1156 ,n355);
    dff g534(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1015), .Q(n4[4]));
    nand g535(n782 ,n3[5] ,n661);
    xnor g536(n1051 ,n216 ,n252);
    dff g537(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1019), .Q(n4[2]));
    nand g538(n818 ,n4[60] ,n351);
    nand g539(n550 ,n1050 ,n354);
    or g540(n1019 ,n807 ,n1011);
    nand g541(n146 ,n3[44] ,n144);
    or g542(n484 ,n7[4] ,n374);
    dff g543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n688), .Q(n3[55]));
    nand g544(n1011 ,n465 ,n856);
    nand g545(n713 ,n595 ,n532);
    nand g546(n76 ,n24 ,n75);
    dff g547(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n863), .Q(n4[38]));
    nand g548(n283 ,n4[29] ,n280);
    nand g549(n878 ,n531 ,n771);
    nand g550(n857 ,n4[1] ,n742);
    or g551(n266 ,n4[21] ,n264);
    xnor g552(n217 ,n4[7] ,n7[7]);
    not g553(n14 ,n3[39]);
    not g554(n366 ,n365);
    nand g555(n157 ,n3[50] ,n156);
    dff g556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n919), .Q(n4[60]));
    xnor g557(n1109 ,n58 ,n79);
    nand g558(n38 ,n3[4] ,n7[4]);
    nand g559(n1092 ,n335 ,n334);
    dff g560(.RN(n1205), .SN(1'b1), .CK(n0), .D(n1268), .Q(n8[1]));
    nand g561(n319 ,n4[47] ,n316);
    nor g562(n1121 ,n103 ,n105);
    or g563(n320 ,n4[48] ,n318);
    nand g564(n799 ,n7[7] ,n632);
    nand g565(n875 ,n415 ,n766);
    nor g566(n399 ,n4[3] ,n374);
    nand g567(n788 ,n7[13] ,n652);
    dff g568(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1033), .Q(n5[2]));
    buf g569(n5[39], 1'b0);
    nand g570(n691 ,n575 ,n454);
    dff g571(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n871), .Q(n4[31]));
    nor g572(n1249 ,n1189 ,n1191);
    nand g573(n701 ,n584 ,n519);
    not g574(n128 ,n127);
    nand g575(n605 ,n3[20] ,n353);
    or g576(n630 ,n380 ,n385);
    dff g577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n687), .Q(n3[56]));
    nand g578(n454 ,n1153 ,n355);
    not g579(n11 ,n3[55]);
    nand g580(n850 ,n4[8] ,n735);
    nand g581(n997 ,n843 ,n942);
    nand g582(n49 ,n3[2] ,n7[2]);
    or g583(n486 ,n7[1] ,n374);
    or g584(n1208 ,n1205 ,n2[14]);
    dff g585(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n936), .Q(n4[46]));
    buf g586(n5[37], 1'b0);
    nand g587(n502 ,n1159 ,n355);
    or g588(n413 ,n377 ,n380);
    nand g589(n663 ,n493 ,n479);
    nand g590(n639 ,n490 ,n479);
    nand g591(n829 ,n4[51] ,n668);
    or g592(n490 ,n7[11] ,n374);
    nand g593(n706 ,n588 ,n524);
    nand g594(n443 ,n1048 ,n354);
    or g595(n1016 ,n806 ,n1010);
    dff g596(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1030), .Q(n5[3]));
    nand g597(n115 ,n3[26] ,n114);
    dff g598(.RN(n1214), .SN(n1223), .CK(n0), .D(n1247), .Q(n7[15]));
    nand g599(n134 ,n3[37] ,n133);
    buf g600(n5[59], 1'b0);
    nand g601(n1006 ,n768 ,n961);
    nor g602(n1268 ,n1196 ,n1194);
    nand g603(n524 ,n1138 ,n378);
    nand g604(n904 ,n426 ,n797);
    xnor g605(n1152 ,n3[51] ,n157);
    nand g606(n549 ,n1116 ,n379);
    nand g607(n1226 ,n1 ,n2[12]);
    not g608(n1191 ,n1190);
    nand g609(n1009 ,n805 ,n854);
    nand g610(n901 ,n443 ,n792);
    dff g611(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n691), .Q(n3[52]));
    nand g612(n1079 ,n309 ,n308);
    nor g613(n744 ,n367 ,n669);
    nand g614(n41 ,n3[14] ,n7[14]);
    nand g615(n125 ,n3[32] ,n123);
    nand g616(n1007 ,n835 ,n963);
    buf g617(n5[42], 1'b0);
    nand g618(n309 ,n4[42] ,n306);
    nor g619(n375 ,n370 ,n371);
    nand g620(n905 ,n449 ,n796);
    xnor g621(n1164 ,n3[63] ,n178);
    nand g622(n597 ,n3[28] ,n376);
    nand g623(n832 ,n7[10] ,n658);
    or g624(n312 ,n4[44] ,n310);
    not g625(n190 ,n4[3]);
    nand g626(n876 ,n440 ,n767);
    nor g627(n103 ,n3[20] ,n102);
    dff g628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n927), .Q(n4[53]));
    dff g629(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n876), .Q(n4[27]));
    nand g630(n821 ,n3[9] ,n654);
    nand g631(n113 ,n3[25] ,n112);
    xnor g632(n1263 ,n8[6] ,n1202);
    nor g633(n1242 ,n1240 ,n1239);
    nand g634(n1090 ,n331 ,n330);
    nand g635(n739 ,n484 ,n669);
    nand g636(n711 ,n593 ,n547);
    nand g637(n704 ,n586 ,n450);
    nand g638(n610 ,n3[63] ,n376);
    nor g639(n96 ,n3[16] ,n95);
    nand g640(n667 ,n487 ,n479);
    nand g641(n541 ,n1123 ,n356);
    nand g642(n244 ,n200 ,n243);
    nand g643(n838 ,n4[44] ,n668);
    nand g644(n973 ,n5[8] ,n890);
    nor g645(n1117 ,n98 ,n96);
    or g646(n29 ,n3[9] ,n7[9]);
    xnor g647(n226 ,n4[4] ,n7[4]);
    or g648(n340 ,n4[58] ,n338);
    nand g649(n196 ,n7[12] ,n183);
    nand g650(n603 ,n3[22] ,n376);
    nor g651(n388 ,n4[11] ,n374);
    nand g652(n612 ,n3[41] ,n376);
    nand g653(n259 ,n4[17] ,n257);
    xnor g654(n1050 ,n218 ,n250);
    nand g655(n236 ,n211 ,n235);
    nor g656(n390 ,n4[5] ,n374);
    or g657(n288 ,n4[32] ,n286);
    nand g658(n680 ,n610 ,n557);
    nand g659(n988 ,n857 ,n957);
    buf g660(n5[31], 1'b0);
    nand g661(n839 ,n4[43] ,n351);
    nand g662(n239 ,n217 ,n238);
    nand g663(n1231 ,n1 ,n2[7]);
    nand g664(n91 ,n39 ,n90);
    nand g665(n912 ,n471 ,n746);
    nand g666(n1229 ,n1 ,n2[9]);
    nand g667(n709 ,n591 ,n527);
    dff g668(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n995), .Q(n4[14]));
    nand g669(n417 ,n1108 ,n354);
    or g670(n278 ,n4[27] ,n276);
    not g671(n956 ,n910);
    or g672(n35 ,n3[7] ,n7[7]);
    nand g673(n210 ,n7[8] ,n186);
    nand g674(n522 ,n1098 ,n379);
    not g675(n359 ,n7[2]);
    nand g676(n672 ,n7[7] ,n478);
    or g677(n262 ,n4[19] ,n260);
    buf g678(n5[23], 1'b0);
    nand g679(n445 ,n1087 ,n356);
    nand g680(n176 ,n3[61] ,n175);
    nand g681(n534 ,n1130 ,n378);
    xnor g682(n56 ,n7[7] ,n3[7]);
    or g683(n290 ,n4[33] ,n288);
    nand g684(n519 ,n1143 ,n354);
    nor g685(n1253 ,n1182 ,n1184);
    nor g686(n1261 ,n1170 ,n1168);
    nand g687(n517 ,n1082 ,n355);
    not g688(n186 ,n4[8]);
    not g689(n183 ,n4[12]);
    nand g690(n682 ,n611 ,n499);
    dff g691(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n880), .Q(n4[24]));
    nand g692(n1059 ,n269 ,n268);
    nand g693(n1096 ,n343 ,n342);
    nand g694(n458 ,n1076 ,n378);
    not g695(n114 ,n113);
    nor g696(n123 ,n18 ,n122);
    nand g697(n488 ,n361 ,n375);
    not g698(n891 ,n859);
    not g699(n364 ,n363);
    xnor g700(n1159 ,n3[58] ,n169);
    nand g701(n654 ,n482 ,n479);
    nand g702(n160 ,n3[52] ,n158);
    nand g703(n198 ,n7[1] ,n184);
    buf g704(n5[19], 1'b0);
    nand g705(n845 ,n4[13] ,n730);
    nand g706(n685 ,n569 ,n502);
    buf g707(n5[25], 1'b0);
    nand g708(n715 ,n597 ,n535);
    not g709(n960 ,n915);
    not g710(n351 ,n350);
    dff g711(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n886), .Q(n4[19]));
    nand g712(n1004 ,n812 ,n959);
    nand g713(n861 ,n460 ,n750);
    dff g714(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n921), .Q(n4[59]));
    nor g715(n116 ,n13 ,n115);
    dff g716(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1036), .Q(n5[0]));
    xnor g717(n1105 ,n53 ,n71);
    nand g718(n816 ,n4[61] ,n668);
    nor g719(n159 ,n3[52] ,n158);
    nand g720(n937 ,n517 ,n837);
    not g721(n378 ,n357);
    buf g722(n5[41], 1'b0);
    or g723(n268 ,n4[22] ,n266);
    nor g724(n130 ,n16 ,n129);
    nand g725(n331 ,n4[53] ,n328);
    not g726(n1167 ,n2[12]);
    nand g727(n1098 ,n348 ,n347);
    nand g728(n929 ,n424 ,n828);
    buf g729(n5[26], 1'b0);
    not g730(n185 ,n4[16]);
    not g731(n189 ,n4[7]);
    nand g732(n803 ,n7[5] ,n635);
    nand g733(n74 ,n28 ,n73);
    or g734(n32 ,n3[15] ,n7[15]);
    not g735(n350 ,n668);
    or g736(n22 ,n3[3] ,n7[3]);
    nand g737(n99 ,n3[17] ,n98);
    not g738(n948 ,n902);
    nand g739(n421 ,n1067 ,n356);
    nand g740(n999 ,n774 ,n893);
    or g741(n664 ,n476 ,n404);
    nand g742(n866 ,n553 ,n758);
    nand g743(n1234 ,n1 ,n2[4]);
    nor g744(n384 ,n4[2] ,n374);
    nand g745(n533 ,n1041 ,n378);
    nand g746(n766 ,n4[28] ,n668);
    nor g747(n642 ,n380 ,n384);
    dff g748(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n923), .Q(n4[57]));
    nand g749(n202 ,n7[14] ,n179);
    nand g750(n537 ,n1127 ,n379);
    nand g751(n1071 ,n293 ,n292);
    not g752(n957 ,n911);
    nand g753(n631 ,n486 ,n479);
    not g754(n1198 ,n1197);
    not g755(n12 ,n3[47]);
    nand g756(n1069 ,n289 ,n288);
    nand g757(n717 ,n599 ,n537);
    nand g758(n453 ,n1044 ,n379);
    nand g759(n614 ,n7[13] ,n478);
    nand g760(n969 ,n5[4] ,n890);
    nand g761(n856 ,n4[2] ,n741);
    not g762(n16 ,n3[35]);
    not g763(n892 ,n872);
    nand g764(n538 ,n1126 ,n378);
    dff g765(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n686), .Q(n3[57]));
    nand g766(n431 ,n1070 ,n379);
    nand g767(n120 ,n3[29] ,n119);
    dff g768(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n888), .Q(n4[17]));
    dff g769(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n990), .Q(n4[11]));
    buf g770(n5[55], 1'b0);
    nand g771(n690 ,n574 ,n507);
    nand g772(n781 ,n4[17] ,n351);
    dff g773(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n710), .Q(n3[33]));
    nor g774(n477 ,n373 ,n379);
    nor g775(n1129 ,n117 ,n119);
    nor g776(n385 ,n4[8] ,n374);
    nand g777(n834 ,n4[47] ,n668);
    not g778(n1184 ,n1183);
    xnor g779(n220 ,n4[2] ,n7[2]);
    nand g780(n862 ,n458 ,n752);
    nand g781(n1190 ,n2[13] ,n1188);
    nand g782(n419 ,n1053 ,n378);
    nor g783(n1188 ,n1167 ,n1187);
    nand g784(n150 ,n3[46] ,n149);
    not g785(n964 ,n940);
    nor g786(n367 ,n362 ,n6[0]);
    dff g787(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1034), .Q(n5[4]));
    nor g788(n145 ,n3[44] ,n144);
    nand g789(n927 ,n462 ,n827);
    not g790(n362 ,n6[2]);
    nand g791(n734 ,n482 ,n669);
    buf g792(n5[17], 1'b0);
    not g793(n193 ,n4[2]);
    dff g794(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n885), .Q(n4[20]));
    nand g795(n998 ,n782 ,n894);
    or g796(n330 ,n4[53] ,n328);
    nand g797(n669 ,n370 ,n480);
    dff g798(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n984), .Q(n4[5]));
    not g799(n481 ,n480);
    nor g800(n1157 ,n166 ,n168);
    nand g801(n459 ,n1040 ,n355);
    nand g802(n699 ,n582 ,n420);
    buf g803(n5[63], 1'b0);
    or g804(n890 ,n375 ,n747);
    nand g805(n474 ,n1111 ,n355);
    nand g806(n295 ,n4[35] ,n292);
    or g807(n1221 ,n1205 ,n2[1]);
    nand g808(n442 ,n1055 ,n355);
    nand g809(n665 ,n489 ,n479);
    nor g810(n398 ,n3[13] ,n374);
    nand g811(n1091 ,n333 ,n332);
    not g812(n955 ,n909);
    nand g813(n311 ,n4[43] ,n308);
    nand g814(n229 ,n220 ,n228);
    nand g815(n897 ,n439 ,n786);
    not g816(n953 ,n907);
    xnor g817(n1116 ,n65 ,n93);
    nand g818(n703 ,n585 ,n521);
    nand g819(n607 ,n3[18] ,n353);
    dff g820(.RN(n1209), .SN(n1225), .CK(n0), .D(n1249), .Q(n7[13]));
    xnor g821(n1138 ,n3[37] ,n132);
    nand g822(n200 ,n7[9] ,n181);
    nand g823(n636 ,n497 ,n479);
    not g824(n184 ,n4[1]);
    nand g825(n723 ,n605 ,n543);
    nand g826(n521 ,n1141 ,n354);
    nand g827(n659 ,n374 ,n414);
    nand g828(n472 ,n1063 ,n354);
    or g829(n635 ,n380 ,n390);
    dff g830(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n703), .Q(n3[40]));
    nand g831(n915 ,n551 ,n813);
    nand g832(n449 ,n1046 ,n356);
    nand g833(n842 ,n4[54] ,n351);
    nand g834(n455 ,n1157 ,n354);
    nand g835(n299 ,n4[37] ,n296);
    or g836(n493 ,n7[6] ,n374);
    xnor g837(n1258 ,n2[4] ,n1173);
    nand g838(n424 ,n1089 ,n379);
    nand g839(n910 ,n468 ,n745);
    nand g840(n422 ,n1147 ,n354);
    nand g841(n852 ,n4[6] ,n737);
    xnor g842(n219 ,n4[1] ,n7[1]);
    nand g843(n287 ,n4[31] ,n284);
    nor g844(n110 ,n3[24] ,n109);
    nand g845(n552 ,n1109 ,n354);
    not g846(n100 ,n99);
    xnor g847(n51 ,n7[9] ,n3[9]);
    nand g848(n1056 ,n263 ,n262);
    or g849(n264 ,n4[20] ,n262);
    xnor g850(n1041 ,n226 ,n232);
    dff g851(.RN(n1220), .SN(n1238), .CK(n0), .D(n1260), .Q(n7[2]));
    or g852(n286 ,n4[31] ,n284);
    or g853(n314 ,n4[45] ,n312);
    nand g854(n572 ,n3[55] ,n353);
    xnor g855(n1154 ,n3[53] ,n160);
    nor g856(n1137 ,n131 ,n133);
    nand g857(n591 ,n3[34] ,n353);
    nand g858(n556 ,n1073 ,n378);
    xor g859(n1023 ,n613 ,n977);
    nand g860(n989 ,n848 ,n948);
    dff g861(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1026), .Q(n5[9]));
    nand g862(n823 ,n4[56] ,n668);
    nand g863(n507 ,n1154 ,n355);
    nand g864(n1055 ,n261 ,n260);
    nand g865(n498 ,n1163 ,n379);
    nor g866(n380 ,n370 ,n366);
    nand g867(n745 ,n7[0] ,n634);
    xnor g868(n1103 ,n59 ,n67);
    nand g869(n571 ,n3[56] ,n353);
    nand g870(n981 ,n850 ,n952);
    xnor g871(n1132 ,n3[31] ,n122);
    not g872(n161 ,n160);
    nand g873(n587 ,n3[38] ,n376);
    nand g874(n863 ,n561 ,n754);
    nand g875(n568 ,n3[59] ,n353);
    nand g876(n975 ,n5[10] ,n890);
    not g877(n1203 ,n1202);
    nand g878(n833 ,n4[48] ,n351);
    nand g879(n611 ,n3[61] ,n353);
    nand g880(n967 ,n5[2] ,n890);
    nand g881(n1078 ,n307 ,n306);
    nand g882(n710 ,n592 ,n528);
    nand g883(n247 ,n212 ,n246);
    nand g884(n812 ,n3[15] ,n649);
    nand g885(n719 ,n601 ,n539);
    xnor g886(n215 ,n4[15] ,n7[15]);
    not g887(n944 ,n898);
    nand g888(n697 ,n581 ,n422);
    nand g889(n446 ,n1047 ,n355);
    nand g890(n602 ,n3[23] ,n376);
    nand g891(n909 ,n457 ,n803);
    xnor g892(n63 ,n7[13] ,n3[13]);
    nand g893(n565 ,n3[45] ,n376);
    xnor g894(n1046 ,n214 ,n242);
    nor g895(n476 ,n1 ,n372);
    or g896(n657 ,n476 ,n394);
    nand g897(n75 ,n44 ,n74);
    nand g898(n426 ,n1102 ,n379);
    nand g899(n882 ,n444 ,n810);
    nor g900(n1161 ,n173 ,n175);
    nand g901(n798 ,n7[8] ,n630);
    nand g902(n794 ,n7[10] ,n626);
    not g903(n175 ,n174);
    buf g904(n5[27], 1'b0);
    nand g905(n106 ,n3[21] ,n105);
    nand g906(n543 ,n1121 ,n354);
    nand g907(n1068 ,n287 ,n286);
    or g908(n620 ,n380 ,n408);
    dff g909(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n865), .Q(n4[36]));
    nand g910(n548 ,n1117 ,n378);
    or g911(n622 ,n380 ,n401);
    nand g912(n692 ,n576 ,n435);
    nand g913(n830 ,n4[50] ,n351);
    dff g914(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n864), .Q(n4[37]));
    nand g915(n1173 ,n2[3] ,n1172);
    xnor g916(n1131 ,n3[30] ,n120);
    buf g917(n5[58], 1'b0);
    nand g918(n848 ,n4[10] ,n733);
    nand g919(n1239 ,n8[1] ,n8[0]);
    or g920(n645 ,n476 ,n398);
    nand g921(n982 ,n851 ,n953);
    dff g922(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1005), .Q(n3[14]));
    nand g923(n853 ,n4[5] ,n738);
    or g924(n27 ,n3[4] ,n7[4]);
    dff g925(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n699), .Q(n3[44]));
    nor g926(n389 ,n3[8] ,n374);
    nand g927(n72 ,n27 ,n71);
    nand g928(n828 ,n4[52] ,n351);
    nand g929(n81 ,n42 ,n80);
    not g930(n355 ,n357);
    dff g931(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n980), .Q(n3[1]));
    or g932(n648 ,n476 ,n403);
    nor g933(n203 ,n187 ,n4[0]);
    dff g934(.RN(n1205), .SN(1'b1), .CK(n0), .D(n1265), .Q(n8[4]));
    nor g935(n1145 ,n145 ,n147);
    dff g936(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1023), .Q(n5[12]));
    nand g937(n820 ,n4[58] ,n351);
    nand g938(n764 ,n4[29] ,n668);
    nand g939(n1094 ,n339 ,n338);
    dff g940(.RN(n1213), .SN(n1230), .CK(n0), .D(n1254), .Q(n7[8]));
    nand g941(n269 ,n4[22] ,n266);
    nand g942(n994 ,n845 ,n944);
    dff g943(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n681), .Q(n3[62]));
    nand g944(n1036 ,n1018 ,n1032);
    not g945(n179 ,n4[14]);
    buf g946(n5[50], 1'b0);
    nand g947(n847 ,n4[11] ,n732);
    not g948(n194 ,n4[13]);
    or g949(n1218 ,n1205 ,n2[4]);
    nand g950(n768 ,n3[13] ,n646);
    nand g951(n1197 ,n8[2] ,n1196);
    nand g952(n933 ,n529 ,n833);
    nand g953(n313 ,n4[44] ,n310);
    or g954(n494 ,n7[13] ,n374);
    nand g955(n547 ,n1133 ,n378);
    nand g956(n451 ,n1045 ,n356);
    nand g957(n881 ,n430 ,n773);
    dff g958(.RN(n1212), .SN(n1229), .CK(n0), .D(n1253), .Q(n7[9]));
    nand g959(n94 ,n32 ,n93);
    xnor g960(n1130 ,n3[29] ,n118);
    nand g961(n40 ,n3[3] ,n7[3]);
    not g962(n947 ,n901);
    nand g963(n553 ,n1072 ,n378);
    nand g964(n729 ,n483 ,n669);
    dff g965(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n862), .Q(n4[39]));
    not g966(n961 ,n920);
    xor g967(n1035 ,n674 ,n970);
    nand g968(n77 ,n48 ,n76);
    nor g969(n1181 ,n1166 ,n1180);
    xnor g970(n1255 ,n2[7] ,n1178);
    nand g971(n916 ,n515 ,n814);
    dff g972(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n711), .Q(n3[32]));
    nand g973(n315 ,n4[45] ,n312);
    or g974(n1032 ,n477 ,n1017);
    or g975(n483 ,n7[14] ,n374);
    nand g976(n1192 ,n2[14] ,n1191);
    or g977(n652 ,n380 ,n391);
    nand g978(n771 ,n4[25] ,n351);
    nand g979(n83 ,n46 ,n82);
    nand g980(n800 ,n7[11] ,n640);
    or g981(n344 ,n4[60] ,n342);
    or g982(n495 ,n7[12] ,n374);
    nand g983(n241 ,n224 ,n240);
    nand g984(n849 ,n4[9] ,n734);
    dff g985(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n689), .Q(n3[54]));
    nand g986(n592 ,n3[33] ,n376);
    or g987(n627 ,n476 ,n382);
    or g988(n282 ,n4[29] ,n280);
    nand g989(n357 ,n367 ,n365);
    nand g990(n545 ,n1119 ,n354);
    or g991(n1220 ,n1205 ,n2[2]);
    nand g992(n428 ,n1061 ,n356);
    or g993(n258 ,n4[17] ,n257);
    nor g994(n396 ,n3[11] ,n374);
    nand g995(n504 ,n1080 ,n356);
    nor g996(n1257 ,n1175 ,n1177);
    nor g997(n377 ,n369 ,n371);
    nor g998(n403 ,n3[15] ,n374);
    not g999(n168 ,n167);
    or g1000(n628 ,n380 ,n387);
    nand g1001(n801 ,n3[1] ,n631);
    nand g1002(n791 ,n3[3] ,n623);
    dff g1003(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n935), .Q(n4[47]));
    dff g1004(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n694), .Q(n3[49]));
    nand g1005(n1240 ,n8[3] ,n8[2]);
    nand g1006(n851 ,n4[7] ,n736);
    buf g1007(n5[45], 1'b0);
    xnor g1008(n1262 ,n1204 ,n8[7]);
    dff g1009(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n722), .Q(n3[21]));
    not g1010(n360 ,n7[8]);
    nand g1011(n887 ,n442 ,n780);
    nand g1012(n1087 ,n325 ,n324);
    nand g1013(n567 ,n3[60] ,n376);
    nand g1014(n660 ,n484 ,n479);
    not g1015(n962 ,n928);
    nand g1016(n554 ,n1114 ,n378);
    not g1017(n1186 ,n1185);
    nand g1018(n908 ,n467 ,n802);
    nand g1019(n598 ,n3[27] ,n376);
    nand g1020(n918 ,n419 ,n783);
    nand g1021(n252 ,n208 ,n251);
    xnor g1022(n1148 ,n3[47] ,n150);
    nand g1023(n273 ,n4[24] ,n270);
    nand g1024(n900 ,n562 ,n790);
    nand g1025(n913 ,n473 ,n748);
    nand g1026(n898 ,n550 ,n788);
    nand g1027(n785 ,n3[4] ,n660);
    or g1028(n653 ,n476 ,n393);
    nand g1029(n741 ,n496 ,n669);
    nand g1030(n1064 ,n279 ,n278);
    dff g1031(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1007), .Q(n3[11]));
    nand g1032(n815 ,n4[62] ,n351);
    nand g1033(n1083 ,n317 ,n316);
    nand g1034(n1238 ,n1 ,n2[2]);
    dff g1035(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n413), .Q(n6[1]));
    or g1036(n274 ,n4[25] ,n272);
    nand g1037(n1088 ,n327 ,n326);
    nand g1038(n348 ,n4[61] ,n344);
    nand g1039(n86 ,n30 ,n85);
    nand g1040(n199 ,n7[7] ,n189);
    nand g1041(n1235 ,n1 ,n2[3]);
    buf g1042(n5[21], 1'b0);
    nand g1043(n523 ,n1139 ,n378);
    nand g1044(n500 ,n1161 ,n355);
    dff g1045(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n659), .Q(n6[2]));
    nor g1046(n1246 ,n1241 ,n1245);
    nand g1047(n732 ,n490 ,n669);
    nand g1048(n965 ,n5[15] ,n890);
    dff g1049(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n860), .Q(n4[41]));
    nand g1050(n797 ,n7[1] ,n629);
    nand g1051(n683 ,n567 ,n500);
    nand g1052(n899 ,n441 ,n789);
    nor g1053(n165 ,n11 ,n164);
    dff g1054(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n988), .Q(n4[1]));
    nand g1055(n574 ,n3[53] ,n376);
    nand g1056(n136 ,n3[38] ,n135);
    nand g1057(n430 ,n1060 ,n356);
    not g1058(n112 ,n111);
    nand g1059(n265 ,n4[20] ,n262);
    nand g1060(n506 ,n1155 ,n355);
    dff g1061(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n873), .Q(n4[30]));
    nand g1062(n874 ,n418 ,n764);
    nand g1063(n45 ,n3[1] ,n7[1]);
    dff g1064(.RN(n1210), .SN(n1227), .CK(n0), .D(n1251), .Q(n7[11]));
    nor g1065(n138 ,n3[40] ,n137);
    nand g1066(n879 ,n429 ,n770);
    dff g1067(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n685), .Q(n3[58]));
    nand g1068(n902 ,n446 ,n794);
    nand g1069(n329 ,n4[52] ,n326);
    nand g1070(n995 ,n844 ,n943);
    nor g1071(n382 ,n3[2] ,n374);
    nand g1072(n227 ,n203 ,n219);
    nand g1073(n71 ,n40 ,n70);
    nand g1074(n934 ,n425 ,n800);
    nand g1075(n656 ,n491 ,n479);
    nand g1076(n508 ,n1094 ,n354);
    nor g1077(n386 ,n4[0] ,n374);
    nand g1078(n570 ,n3[57] ,n353);
    nand g1079(n92 ,n26 ,n91);
    xnor g1080(n222 ,n4[12] ,n7[12]);
    nand g1081(n931 ,n445 ,n830);
    nand g1082(n722 ,n604 ,n542);
    not g1083(n379 ,n357);
    nand g1084(n819 ,n4[59] ,n668);
    not g1085(n945 ,n899);
    nand g1086(n676 ,n7[3] ,n478);
    nand g1087(n228 ,n198 ,n227);
    nand g1088(n671 ,n7[8] ,n478);
    nor g1089(n152 ,n3[48] ,n151);
    not g1090(n188 ,n4[15]);
    nand g1091(n1178 ,n2[6] ,n1177);
    or g1092(n489 ,n7[7] ,n374);
    dff g1093(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n878), .Q(n4[25]));
    not g1094(n356 ,n357);
    nand g1095(n425 ,n1112 ,n379);
    nand g1096(n153 ,n3[48] ,n151);
    nor g1097(n641 ,n380 ,n399);
    not g1098(n192 ,n4[4]);
    dff g1099(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n714), .Q(n3[29]));
    not g1100(n347 ,n346);
    xnor g1101(n1259 ,n2[3] ,n1171);
    buf g1102(n5[62], 1'b0);
    dff g1103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n932), .Q(n4[49]));
    dff g1104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n708), .Q(n3[35]));
    nor g1105(n402 ,n4[4] ,n374);
    nor g1106(n117 ,n3[28] ,n116);
    dff g1107(.RN(n1207), .SN(n1226), .CK(n0), .D(n1250), .Q(n7[12]));
    nand g1108(n770 ,n7[6] ,n664);
    or g1109(n626 ,n380 ,n395);
    nand g1110(n714 ,n596 ,n534);
    nand g1111(n855 ,n4[3] ,n740);
    not g1112(n147 ,n146);
    nand g1113(n1065 ,n281 ,n280);
    nor g1114(n807 ,n359 ,n642);
    nand g1115(n802 ,n7[6] ,n633);
    or g1116(n632 ,n380 ,n407);
    nand g1117(n501 ,n1160 ,n355);
    nor g1118(n1174 ,n1165 ,n1173);
    xnor g1119(n1047 ,n213 ,n244);
    or g1120(n342 ,n4[59] ,n340);
    nand g1121(n618 ,n7[11] ,n478);
    nand g1122(n974 ,n5[9] ,n890);
    nor g1123(n1201 ,n8[5] ,n1200);
    nand g1124(n576 ,n3[51] ,n353);
    xor g1125(n1053 ,n256 ,n4[16]);
    nand g1126(n461 ,n1058 ,n378);
    nand g1127(n44 ,n3[5] ,n7[5]);
    xnor g1128(n58 ,n7[8] ,n3[8]);
    nand g1129(n464 ,n1057 ,n356);
    nand g1130(n971 ,n5[6] ,n890);
    nand g1131(n608 ,n3[17] ,n353);
    nand g1132(n171 ,n3[58] ,n170);
    xnor g1133(n1135 ,n3[34] ,n127);
    dff g1134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n883), .Q(n4[21]));
    dff g1135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n726), .Q(n3[17]));
    nand g1136(n661 ,n492 ,n479);
    not g1137(n1177 ,n1176);
    dff g1138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1029), .Q(n5[6]));
    nand g1139(n466 ,n1096 ,n354);
    or g1140(n372 ,n6[2] ,n364);
    nand g1141(n670 ,n368 ,n480);
    nand g1142(n339 ,n4[57] ,n336);
    dff g1143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n684), .Q(n3[59]));
    nand g1144(n1000 ,n809 ,n892);
    nand g1145(n209 ,n7[3] ,n190);
    dff g1146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n680), .Q(n3[63]));
    dff g1147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n696), .Q(n3[47]));
    nand g1148(n854 ,n4[4] ,n739);
    or g1149(n26 ,n3[14] ,n7[14]);
    nor g1150(n1153 ,n159 ,n161);
    nand g1151(n84 ,n33 ,n83);
    nand g1152(n1176 ,n2[5] ,n1174);
    nand g1153(n559 ,n1074 ,n378);
    nand g1154(n1245 ,n8[4] ,n1244);
    nand g1155(n544 ,n1120 ,n354);
    not g1156(n958 ,n912);
    nand g1157(n1058 ,n267 ,n266);
    xor g1158(n1101 ,n7[0] ,n3[0]);
    nand g1159(n343 ,n4[59] ,n340);
    nand g1160(n716 ,n598 ,n536);
    nand g1161(n601 ,n3[24] ,n376);
    nand g1162(n420 ,n1145 ,n356);
    dff g1163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n700), .Q(n3[43]));
    xnor g1164(n53 ,n7[4] ,n3[4]);
    nand g1165(n557 ,n1164 ,n354);
    dff g1166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n683), .Q(n3[60]));
    nor g1167(n137 ,n14 ,n136);
    nand g1168(n503 ,n1158 ,n379);
    nand g1169(n694 ,n578 ,n511);
    nand g1170(n935 ,n514 ,n834);
    xnor g1171(n65 ,n7[15] ,n3[15]);
    dff g1172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n718), .Q(n3[25]));
    xnor g1173(n223 ,n4[5] ,n7[5]);
    nand g1174(n450 ,n1140 ,n355);
    nand g1175(n837 ,n4[45] ,n668);
    xnor g1176(n1160 ,n3[59] ,n171);
    nor g1177(n394 ,n3[12] ,n374);
    nand g1178(n673 ,n7[6] ,n478);
    nand g1179(n976 ,n5[11] ,n890);
    nor g1180(n346 ,n4[61] ,n344);
    xnor g1181(n1111 ,n60 ,n83);
    nand g1182(n118 ,n3[28] ,n116);
    nand g1183(n462 ,n1090 ,n356);
    nand g1184(n990 ,n847 ,n947);
    nand g1185(n780 ,n4[18] ,n351);
    or g1186(n662 ,n476 ,n383);
    xnor g1187(n1038 ,n219 ,n203);
    or g1188(n306 ,n4[41] ,n304);
    dff g1189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n701), .Q(n3[42]));
    nand g1190(n746 ,n7[0] ,n644);
    nand g1191(n586 ,n3[39] ,n353);
    or g1192(n33 ,n3[10] ,n7[10]);
    nand g1193(n779 ,n4[19] ,n668);
    dff g1194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n716), .Q(n3[27]));
    nand g1195(n966 ,n5[1] ,n890);
    nand g1196(n702 ,n612 ,n520);
    xnor g1197(n1110 ,n51 ,n81);
    nand g1198(n208 ,n7[13] ,n194);
    nand g1199(n696 ,n580 ,n513);
    or g1200(n30 ,n3[11] ,n7[11]);
    dff g1201(.RN(n1205), .SN(1'b1), .CK(n0), .D(n1206), .Q(n8[0]));
    nand g1202(n651 ,n483 ,n479);
    nand g1203(n930 ,n448 ,n829);
    or g1204(n292 ,n4[34] ,n290);
    nand g1205(n922 ,n512 ,n820);
    nand g1206(n1232 ,n1 ,n2[6]);
    nor g1207(n655 ,n476 ,n389);
    nand g1208(n721 ,n603 ,n541);
    nand g1209(n261 ,n4[18] ,n258);
    xnor g1210(n1146 ,n3[45] ,n146);
    dff g1211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n938), .Q(n4[44]));
    nand g1212(n536 ,n1128 ,n354);
    nand g1213(n20 ,n3[11] ,n7[11]);
    not g1214(n354 ,n357);
    nand g1215(n728 ,n485 ,n669);
    nand g1216(n48 ,n3[6] ,n7[6]);
    not g1217(n18 ,n3[31]);
    dff g1218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n682), .Q(n3[61]));
    or g1219(n326 ,n4[51] ,n324);
    xnor g1220(n1158 ,n3[57] ,n167);
    dff g1221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n882), .Q(n4[22]));
    dff g1222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n992), .Q(n4[12]));
    xnor g1223(n1260 ,n2[2] ,n1169);
    nand g1224(n174 ,n3[60] ,n172);
    or g1225(n625 ,n380 ,n388);
    nand g1226(n871 ,n423 ,n762);
    or g1227(n328 ,n4[52] ,n326);
    nand g1228(n155 ,n3[49] ,n154);
    nand g1229(n1073 ,n297 ,n296);
    xnor g1230(n1106 ,n54 ,n73);
    nand g1231(n1080 ,n311 ,n310);
    or g1232(n304 ,n4[40] ,n302);
    dff g1233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1022), .Q(n5[13]));
    nand g1234(n516 ,n1146 ,n356);
    nand g1235(n167 ,n3[56] ,n165);
    not g1236(n353 ,n352);
    not g1237(n1166 ,n2[8]);
    nand g1238(n291 ,n4[33] ,n288);
    dff g1239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n727), .Q(n3[16]));
    buf g1240(n5[51], 1'b0);
    nand g1241(n877 ,n472 ,n769);
    dff g1242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n981), .Q(n4[8]));
    xnor g1243(n55 ,n7[6] ,n3[6]);
    nor g1244(n393 ,n3[3] ,n374);
    nor g1245(n383 ,n3[5] ,n374);
    nor g1246(n400 ,n3[1] ,n374);
    nand g1247(n1070 ,n291 ,n290);
    not g1248(n1170 ,n1169);
    nand g1249(n561 ,n1075 ,n356);
    nand g1250(n88 ,n31 ,n87);
    nand g1251(n87 ,n20 ,n86);
    nand g1252(n589 ,n3[36] ,n353);
    nand g1253(n584 ,n3[42] ,n376);
    nand g1254(n1225 ,n1 ,n2[13]);
    or g1255(n633 ,n380 ,n381);
    or g1256(n31 ,n3[12] ,n7[12]);
    nand g1257(n232 ,n209 ,n231);
    nand g1258(n1061 ,n273 ,n272);
    nand g1259(n889 ,n787 ,n785);
    nand g1260(n50 ,n3[0] ,n7[0]);
    xnor g1261(n1248 ,n2[14] ,n1190);
    nand g1262(n429 ,n1107 ,n355);
    nand g1263(n928 ,n751 ,n825);
    dff g1264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1002), .Q(n3[9]));
    or g1265(n298 ,n4[37] ,n296);
    xnor g1266(n1104 ,n52 ,n69);
    not g1267(n17 ,n3[23]);
    nand g1268(n551 ,n1115 ,n354);
    nor g1269(n102 ,n9 ,n101);
    xnor g1270(n1151 ,n3[50] ,n155);
    nand g1271(n432 ,n1106 ,n356);
    nand g1272(n1066 ,n283 ,n282);
    nand g1273(n555 ,n1071 ,n354);
    or g1274(n338 ,n4[57] ,n336);
    xnor g1275(n1162 ,n3[61] ,n174);
    nor g1276(n409 ,n3[4] ,n374);
    or g1277(n302 ,n4[39] ,n300);
    nand g1278(n69 ,n49 ,n68);
    nand g1279(n479 ,n376 ,n374);
    nand g1280(n439 ,n1051 ,n379);
    nand g1281(n271 ,n4[23] ,n268);
    nand g1282(n341 ,n4[58] ,n338);
    nand g1283(n747 ,n357 ,n670);
    nand g1284(n237 ,n225 ,n236);
    not g1285(n126 ,n125);
    nor g1286(n411 ,n3[0] ,n374);
    buf g1287(n5[33], 1'b0);
    nand g1288(n767 ,n4[27] ,n668);
    or g1289(n24 ,n3[6] ,n7[6]);
    nand g1290(n230 ,n204 ,n229);
    dff g1291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n867), .Q(n4[34]));
    nand g1292(n39 ,n3[13] ,n7[13]);
    nand g1293(n70 ,n22 ,n69);
    nand g1294(n737 ,n493 ,n669);
    dff g1295(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n887), .Q(n4[18]));
    not g1296(n181 ,n4[9]);
    buf g1297(n5[18], 1'b0);
    nand g1298(n333 ,n4[54] ,n330);
    or g1299(n294 ,n4[35] ,n292);
    nor g1300(n1168 ,n2[1] ,n1246);
    dff g1301(.RN(n1205), .SN(1'b1), .CK(n0), .D(n1264), .Q(n8[5]));
    dff g1302(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n861), .Q(n4[40]));
    buf g1303(n5[48], 1'b0);
    or g1304(n296 ,n4[36] ,n294);
    or g1305(n1213 ,n1205 ,n2[8]);
    nand g1306(n646 ,n494 ,n479);
    xor g1307(n1026 ,n679 ,n974);
    nand g1308(n85 ,n47 ,n84);
    nor g1309(n395 ,n4[10] ,n374);
    nand g1310(n433 ,n1056 ,n355);
    nand g1311(n512 ,n1095 ,n356);
    nand g1312(n991 ,n858 ,n958);
    xnor g1313(n1156 ,n3[55] ,n164);
    nor g1314(n23 ,n3[1] ,n7[1]);
    nand g1315(n68 ,n25 ,n67);
    xnor g1316(n1127 ,n3[26] ,n113);
    buf g1317(n5[56], 1'b0);
    dff g1318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n697), .Q(n3[46]));
    nand g1319(n444 ,n1059 ,n355);
    nand g1320(n579 ,n3[48] ,n376);
    nand g1321(n880 ,n428 ,n772);
    nand g1322(n983 ,n852 ,n954);
    not g1323(n121 ,n120);
    buf g1324(n5[44], 1'b0);
    xnor g1325(n1142 ,n3[41] ,n139);
    dff g1326(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n987), .Q(n3[2]));
    nand g1327(n826 ,n3[14] ,n651);
    nand g1328(n985 ,n804 ,n956);
    nand g1329(n178 ,n3[62] ,n177);
    nand g1330(n1076 ,n303 ,n302);
    nand g1331(n686 ,n570 ,n503);
    dff g1332(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n933), .Q(n4[48]));
    nand g1333(n528 ,n1134 ,n354);
    or g1334(n284 ,n4[30] ,n282);
    nand g1335(n754 ,n4[38] ,n668);
    xnor g1336(n1250 ,n2[12] ,n1187);
    nor g1337(n387 ,n4[9] ,n374);
    buf g1338(n5[24], 1'b0);
    dff g1339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n913), .Q(n4[42]));
    xnor g1340(n213 ,n4[10] ,n7[10]);
    dff g1341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n985), .Q(n3[0]));
    nand g1342(n122 ,n3[30] ,n121);
    or g1343(n308 ,n4[42] ,n306);
    nand g1344(n289 ,n4[32] ,n286);
    nand g1345(n162 ,n3[53] ,n161);
    nand g1346(n514 ,n1084 ,n355);
    dff g1347(.RN(n1217), .SN(n1233), .CK(n0), .D(n1257), .Q(n7[5]));
    xor g1348(n1034 ,n675 ,n969);
    nand g1349(n926 ,n558 ,n842);
    dff g1350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n918), .Q(n4[16]));
    xnor g1351(n1143 ,n3[42] ,n141);
    nand g1352(n414 ,n6[2] ,n353);
    nand g1353(n1067 ,n285 ,n284);
    nand g1354(n240 ,n199 ,n239);
    dff g1355(.RN(n1211), .SN(n1228), .CK(n0), .D(n1252), .Q(n7[10]));
    not g1356(n177 ,n176);
    nand g1357(n583 ,n3[43] ,n376);
    nand g1358(n527 ,n1135 ,n354);
    nand g1359(n805 ,n7[4] ,n637);
    nand g1360(n529 ,n1085 ,n378);
    nor g1361(n778 ,n360 ,n655);
    nand g1362(n520 ,n1142 ,n355);
    not g1363(n15 ,n3[43]);
    dff g1364(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n693), .Q(n3[50]));
    or g1365(n638 ,n476 ,n410);
    not g1366(n1205 ,n1);
    nand g1367(n525 ,n1137 ,n354);
    nor g1368(n1125 ,n110 ,n112);
    nand g1369(n824 ,n4[55] ,n351);
    nand g1370(n1237 ,n1 ,n2[0]);
    nand g1371(n756 ,n3[8] ,n667);
    nand g1372(n1199 ,n8[3] ,n1198);
    nand g1373(n546 ,n1118 ,n354);
    nand g1374(n467 ,n1043 ,n378);
    xnor g1375(n1118 ,n3[17] ,n97);
    xnor g1376(n225 ,n4[6] ,n7[6]);
    buf g1377(n5[34], 1'b0);
    nand g1378(n1183 ,n2[9] ,n1181);
    nand g1379(n920 ,n554 ,n817);
    xnor g1380(n52 ,n7[3] ,n3[3]);
    nand g1381(n303 ,n4[39] ,n300);
    nand g1382(n513 ,n1148 ,n355);
    buf g1383(n5[46], 1'b0);
    nand g1384(n763 ,n4[30] ,n668);
    nand g1385(n95 ,n43 ,n94);
    nand g1386(n143 ,n3[42] ,n142);
    dff g1387(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n723), .Q(n3[20]));
    nand g1388(n860 ,n470 ,n749);
    nand g1389(n941 ,n522 ,n816);
    nand g1390(n924 ,n509 ,n823);
    nand g1391(n615 ,n7[14] ,n478);
    nand g1392(n285 ,n4[30] ,n282);
    not g1393(n154 ,n153);
    nand g1394(n205 ,n7[10] ,n195);
    nor g1395(n1141 ,n138 ,n140);
    nand g1396(n748 ,n4[42] ,n351);
    xnor g1397(n216 ,n4[14] ,n7[14]);
    not g1398(n149 ,n148);
    not g1399(n1014 ,n1009);
    xnor g1400(n214 ,n4[9] ,n7[9]);
    dff g1401(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n712), .Q(n3[31]));
    or g1402(n666 ,n476 ,n405);
    buf g1403(n5[22], 1'b0);
    dff g1404(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n707), .Q(n3[36]));
    or g1405(n332 ,n4[54] ,n330);
    nand g1406(n79 ,n36 ,n78);
    nand g1407(n108 ,n3[22] ,n107);
    xnor g1408(n1049 ,n222 ,n248);
    nand g1409(n1017 ,n7[0] ,n1012);
    dff g1410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n717), .Q(n3[26]));
    dff g1411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n720), .Q(n3[23]));
    or g1412(n1211 ,n1205 ,n2[10]);
    nand g1413(n970 ,n5[5] ,n890);
    or g1414(n621 ,n476 ,n409);
    xnor g1415(n1147 ,n3[46] ,n148);
    nand g1416(n588 ,n3[37] ,n376);
    nor g1417(n172 ,n10 ,n171);
    nand g1418(n762 ,n4[31] ,n668);
    nand g1419(n758 ,n4[35] ,n668);
    nor g1420(n668 ,n380 ,n481);
    buf g1421(n5[47], 1'b0);
    nand g1422(n1062 ,n275 ,n274);
    dff g1423(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n706), .Q(n3[37]));
    or g1424(n66 ,n50 ,n23);
    dff g1425(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n881), .Q(n4[23]));
    nand g1426(n939 ,n504 ,n839);
    nand g1427(n776 ,n4[21] ,n668);
    or g1428(n1212 ,n1205 ,n2[9]);
    dff g1429(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n986), .Q(n4[9]));
    nor g1430(n408 ,n4[14] ,n374);
    not g1431(n156 ,n155);
    nand g1432(n1012 ,n5[0] ,n890);
    xor g1433(n1029 ,n673 ,n971);
    dff g1434(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n917), .Q(n4[62]));
    nor g1435(n407 ,n4[7] ,n374);
    nor g1436(n365 ,n6[1] ,n1);
    nand g1437(n921 ,n466 ,n819);
    nand g1438(n371 ,n6[1] ,n358);
    not g1439(n893 ,n879);
    nand g1440(n718 ,n600 ,n538);
    dff g1441(.RN(n1221), .SN(n1236), .CK(n0), .D(n1261), .Q(n7[1]));
    buf g1442(n5[43], 1'b0);
    not g1443(n98 ,n97);
    nand g1444(n705 ,n587 ,n523);
    dff g1445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1004), .Q(n3[15]));
    xnor g1446(n1119 ,n3[18] ,n99);
    not g1447(n959 ,n914);
    xnor g1448(n57 ,n7[1] ,n3[1]);
    nand g1449(n687 ,n571 ,n455);
    xnor g1450(n1155 ,n3[54] ,n162);
    nand g1451(n67 ,n45 ,n66);
    dff g1452(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n692), .Q(n3[51]));
    nand g1453(n465 ,n1039 ,n356);
    nand g1454(n468 ,n1101 ,n356);
    nand g1455(n1195 ,n8[1] ,n8[0]);
    nor g1456(n404 ,n3[6] ,n374);
    xnor g1457(n1267 ,n8[2] ,n1195);
    nand g1458(n263 ,n4[19] ,n260);
    nand g1459(n790 ,n7[12] ,n622);
    nand g1460(n1002 ,n821 ,n891);
    dff g1461(.RN(n1215), .SN(n1232), .CK(n0), .D(n1256), .Q(n7[6]));
    nand g1462(n678 ,n7[1] ,n478);
    nand g1463(n772 ,n4[24] ,n351);
    nand g1464(n846 ,n4[12] ,n731);
    nand g1465(n317 ,n4[46] ,n314);
    dff g1466(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n982), .Q(n4[7]));
    nand g1467(n1057 ,n265 ,n264);
    nand g1468(n132 ,n3[36] ,n130);
    nand g1469(n251 ,n218 ,n250);
    nand g1470(n996 ,n438 ,n895);
    nand g1471(n688 ,n572 ,n505);
    not g1472(n1244 ,n1243);
    dff g1473(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n941), .Q(n4[61]));
    not g1474(n9 ,n3[19]);
    nand g1475(n577 ,n3[50] ,n376);
    nand g1476(n37 ,n3[12] ,n7[12]);
    xor g1477(n1100 ,n4[63] ,n349);
    nand g1478(n858 ,n4[0] ,n743);
endmodule
