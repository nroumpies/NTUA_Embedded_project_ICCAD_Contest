module top (n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [63:0] n6;
    wire [63:0] n7;
    wire [63:0] n8;
    wire [63:0] n9;
    wire [63:0] n10;
    wire [63:0] n11;
    wire [2:0] n12;
    wire [3:0] n13;
    wire [15:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
    wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
    wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
    wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
    wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
    wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
    wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
    wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
    wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
    wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
    wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
    wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
    wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
    wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
    wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
    wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
    wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
    wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
    wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
    wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
    wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
    wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
    wire n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742;
    wire n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750;
    wire n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758;
    wire n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766;
    wire n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774;
    wire n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782;
    wire n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790;
    wire n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798;
    wire n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806;
    wire n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814;
    wire n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822;
    wire n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
    wire n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838;
    wire n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846;
    wire n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854;
    wire n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
    wire n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870;
    wire n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878;
    wire n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886;
    wire n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894;
    wire n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902;
    wire n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910;
    wire n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918;
    wire n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
    wire n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934;
    wire n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
    wire n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950;
    wire n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958;
    wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
    wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974;
    wire n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982;
    wire n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990;
    wire n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998;
    wire n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
    wire n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014;
    wire n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022;
    wire n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;
    wire n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038;
    wire n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046;
    wire n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054;
    wire n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062;
    wire n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070;
    wire n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078;
    wire n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086;
    wire n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094;
    wire n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102;
    wire n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110;
    wire n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118;
    wire n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126;
    wire n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134;
    wire n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142;
    wire n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150;
    wire n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158;
    wire n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166;
    wire n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174;
    wire n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182;
    wire n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190;
    wire n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198;
    wire n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206;
    wire n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214;
    wire n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222;
    wire n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230;
    wire n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238;
    wire n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246;
    wire n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254;
    wire n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262;
    wire n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270;
    wire n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278;
    wire n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286;
    wire n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294;
    wire n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302;
    wire n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310;
    wire n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318;
    wire n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326;
    wire n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334;
    wire n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342;
    wire n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350;
    wire n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358;
    wire n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366;
    wire n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374;
    wire n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382;
    wire n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390;
    wire n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398;
    wire n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406;
    wire n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414;
    wire n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422;
    wire n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430;
    wire n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438;
    wire n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446;
    wire n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454;
    wire n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462;
    wire n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470;
    wire n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478;
    wire n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486;
    wire n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494;
    wire n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502;
    wire n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510;
    wire n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518;
    wire n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526;
    wire n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534;
    wire n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542;
    wire n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550;
    wire n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558;
    wire n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566;
    wire n2567;
    nor g0(n883 ,n2510 ,n11[37]);
    dff g1(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1973), .Q(n8[7]));
    nor g2(n861 ,n648 ,n860);
    nand g3(n1616 ,n1306 ,n1487);
    xnor g4(n4[19] ,n2112 ,n8[19]);
    nand g5(n1454 ,n2249 ,n1289);
    xnor g6(n2555 ,n710 ,n871);
    xnor g7(n1000 ,n11[37] ,n2542);
    nand g8(n1018 ,n938 ,n1017);
    xnor g9(n2559 ,n706 ,n875);
    nor g10(n1080 ,n915 ,n1079);
    nand g11(n1732 ,n1233 ,n1499);
    xnor g12(n5[2] ,n2110 ,n6[2]);
    xnor g13(n437 ,n11[40] ,n2187);
    nand g14(n538 ,n368 ,n537);
    xnor g15(n2444 ,n2066 ,n2445);
    xnor g16(n5[5] ,n2102 ,n6[5]);
    xnor g17(n2412 ,n986 ,n1080);
    dff g18(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1900), .Q(n6[43]));
    nand g19(n1854 ,n1443 ,n1656);
    xnor g20(n2183 ,n2[67] ,n2078);
    or g21(n1303 ,n8[50] ,n1193);
    nand g22(n1430 ,n2266 ,n1289);
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1970), .Q(n8[9]));
    nor g24(n1031 ,n989 ,n1030);
    xnor g25(n2327 ,n2078 ,n2[19]);
    or g26(n1392 ,n6[32] ,n1292);
    nor g27(n1164 ,n9[53] ,n1155);
    xnor g28(n2163 ,n594 ,n384);
    nand g29(n597 ,n402 ,n596);
    xnor g30(n2506 ,n2065 ,n2507);
    nor g31(n817 ,n659 ,n816);
    nand g32(n1694 ,n1288 ,n1501);
    nand g33(n2020 ,n9[57] ,n1914);
    xnor g34(n2344 ,n2065 ,n2[36]);
    or g35(n1219 ,n6[4] ,n1196);
    or g36(n1376 ,n7[51] ,n1199);
    xnor g37(n2502 ,n2503 ,n2068);
    xnor g38(n2498 ,n2499 ,n2067);
    or g39(n1228 ,n7[24] ,n1195);
    nand g40(n241 ,n67 ,n240);
    nor g41(n776 ,n731 ,n775);
    xnor g42(n3[5] ,n2102 ,n7[5]);
    nand g43(n937 ,n2448 ,n11[38]);
    xnor g44(n409 ,n11[36] ,n2231);
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1916), .Q(n8[43]));
    nand g46(n105 ,n2353 ,n11[45]);
    not g47(n500 ,n499);
    nand g48(n1698 ,n1298 ,n1489);
    nor g49(n1120 ,n881 ,n1119);
    nand g50(n336 ,n2219 ,n11[40]);
    xnor g51(n2237 ,n2[121] ,n2071);
    nand g52(n1807 ,n1296 ,n1486);
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1979), .Q(n8[2]));
    nand g54(n938 ,n2450 ,n11[39]);
    not g55(n942 ,n941);
    nor g56(n1097 ,n949 ,n1096);
    or g57(n1286 ,n8[6] ,n1197);
    nor g58(n1035 ,n993 ,n1034);
    xnor g59(n176 ,n11[41] ,n2365);
    xnor g60(n944 ,n11[43] ,n2554);
    xnor g61(n2272 ,n147 ,n246);
    nand g62(n1480 ,n2377 ,n1289);
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2012), .Q(n13[0]));
    or g64(n1267 ,n6[59] ,n1186);
    nor g65(n925 ,n2556 ,n11[44]);
    or g66(n1345 ,n6[27] ,n1186);
    nand g67(n1545 ,n2144 ,n1289);
    nand g68(n1483 ,n2421 ,n1289);
    not g69(n444 ,n443);
    nand g70(n1469 ,n2428 ,n1289);
    xnor g71(n2476 ,n2066 ,n2477);
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2005), .Q(n7[47]));
    nand g73(n2062 ,n2027 ,n2044);
    nor g74(n1102 ,n928 ,n1101);
    nor g75(n881 ,n2552 ,n11[42]);
    xnor g76(n2261 ,n184 ,n224);
    nand g77(n343 ,n2230 ,n11[35]);
    nand g78(n1781 ,n1359 ,n1493);
    nand g79(n1418 ,n2276 ,n1289);
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1885), .Q(n6[51]));
    xnor g81(n2173 ,n614 ,n439);
    xnor g82(n2246 ,n177 ,n194);
    nand g83(n11[42] ,n2076 ,n2071);
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1920), .Q(n6[36]));
    nand g85(n1802 ,n1352 ,n1493);
    nand g86(n85 ,n2327 ,n11[35]);
    nor g87(n666 ,n2[35] ,n2[99]);
    or g88(n1326 ,n8[27] ,n1186);
    nand g89(n1606 ,n2293 ,n1289);
    xnor g90(n5[27] ,n2105 ,n6[27]);
    nand g91(n1683 ,n1276 ,n1495);
    nand g92(n79 ,n2317 ,n11[41]);
    nor g93(n1107 ,n987 ,n1106);
    nor g94(n1112 ,n929 ,n1111);
    xnor g95(n4[61] ,n2103 ,n8[61]);
    nand g96(n2041 ,n10[6] ,n2031);
    nand g97(n1686 ,n1274 ,n1492);
    or g98(n29 ,n2312 ,n11[36]);
    not g99(n394 ,n393);
    or g100(n37 ,n2327 ,n11[35]);
    nand g101(n306 ,n108 ,n305);
    nand g102(n1858 ,n1447 ,n1659);
    nand g103(n316 ,n2370 ,n315);
    nand g104(n1551 ,n2381 ,n1289);
    nor g105(n1072 ,n895 ,n1071);
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2062), .Q(n10[1]));
    xnor g107(n2463 ,n735 ,n779);
    nand g108(n2036 ,n10[11] ,n2031);
    nand g109(n1743 ,n1330 ,n1489);
    xnor g110(n2224 ,n2[108] ,n2079);
    nand g111(n1404 ,n2285 ,n1289);
    nor g112(n1498 ,n1168 ,n1291);
    nand g113(n575 ,n387 ,n574);
    nand g114(n1925 ,n1531 ,n1723);
    nand g115(n1818 ,n1551 ,n1807);
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1996), .Q(n6[11]));
    xnor g117(n407 ,n11[33] ,n2212);
    nor g118(n785 ,n632 ,n784);
    nand g119(n1533 ,n2152 ,n1289);
    xnor g120(n3[21] ,n2102 ,n7[21]);
    nor g121(n662 ,n2[41] ,n2[105]);
    nand g122(n224 ,n128 ,n223);
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1941), .Q(n6[29]));
    nor g124(n1195 ,n1141 ,n1155);
    xnor g125(n2198 ,n2[82] ,n2068);
    nand g126(n243 ,n30 ,n242);
    nor g127(n812 ,n696 ,n811);
    xnor g128(n2347 ,n2074 ,n2[39]);
    xnor g129(n2443 ,n717 ,n759);
    xnor g130(n973 ,n11[44] ,n2524);
    nand g131(n1919 ,n1421 ,n1719);
    xnor g132(n694 ,n2[45] ,n2[109]);
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1827), .Q(n6[7]));
    nand g134(n88 ,n2328 ,n11[36]);
    nand g135(n11[34] ,n2078 ,n2073);
    or g136(n1332 ,n6[47] ,n1194);
    nand g137(n1508 ,n2274 ,n1289);
    nand g138(n1833 ,n1419 ,n1631);
    nor g139(n805 ,n676 ,n804);
    nand g140(n533 ,n470 ,n532);
    or g141(n22 ,n2321 ,n11[45]);
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2002), .Q(n6[12]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1953), .Q(n8[18]));
    xnor g144(n4[17] ,n2114 ,n8[17]);
    not g145(n458 ,n457);
    xnor g146(n2229 ,n2[113] ,n2073);
    not g147(n2076 ,n9[59]);
    nor g148(n656 ,n2[25] ,n2[89]);
    dff g149(.RN(1'b1), .SN(n2567), .CK(n0), .D(n9[55]), .Q(n14[9]));
    nand g150(n340 ,n2215 ,n11[36]);
    nor g151(n1090 ,n921 ,n1089);
    not g152(n381 ,n380);
    xnor g153(n443 ,n11[42] ,n2189);
    xnor g154(n3[4] ,n2100 ,n7[4]);
    nand g155(n1830 ,n1416 ,n1625);
    nor g156(n1494 ,n1169 ,n1291);
    nand g157(n1664 ,n1253 ,n1487);
    nand g158(n1812 ,n1475 ,n1474);
    not g159(n2070 ,n9[56]);
    nor g160(n1147 ,n10[0] ,n10[1]);
    not g161(n492 ,n491);
    nand g162(n379 ,n2226 ,n11[31]);
    not g163(n313 ,n312);
    or g164(n1386 ,n7[44] ,n1187);
    xnor g165(n966 ,n2442 ,n11[35]);
    not g166(n1141 ,n10[8]);
    xnor g167(n447 ,n11[39] ,n2218);
    xnor g168(n981 ,n11[42] ,n2456);
    nand g169(n1762 ,n1302 ,n1499);
    xnor g170(n449 ,n11[44] ,n2191);
    nand g171(n366 ,n2221 ,n11[42]);
    or g172(n1270 ,n8[34] ,n1193);
    nand g173(n1685 ,n1269 ,n1489);
    nand g174(n1535 ,n2176 ,n1289);
    xnor g175(n3[30] ,n2113 ,n7[30]);
    nor g176(n637 ,n2[34] ,n2[98]);
    xnor g177(n2252 ,n170 ,n206);
    or g178(n62 ,n2364 ,n11[40]);
    nand g179(n1992 ,n1539 ,n1790);
    or g180(n1390 ,n7[16] ,n1292);
    or g181(n19 ,n2319 ,n11[43]);
    nand g182(n1922 ,n1413 ,n1722);
    nand g183(n1797 ,n1378 ,n1501);
    xnor g184(n692 ,n2[46] ,n2[110]);
    nor g185(n1160 ,n9[49] ,n1155);
    not g186(n490 ,n489);
    nand g187(n1521 ,n2170 ,n1289);
    nand g188(n1915 ,n1177 ,n1814);
    or g189(n1275 ,n6[52] ,n1196);
    not g190(n412 ,n411);
    nand g191(n568 ,n334 ,n567);
    or g192(n1346 ,n8[10] ,n1198);
    xnor g193(n2537 ,n733 ,n853);
    nor g194(n1488 ,n1164 ,n1291);
    nor g195(n1081 ,n986 ,n1080);
    nand g196(n1548 ,n2141 ,n1289);
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1824), .Q(n6[8]));
    xnor g198(n693 ,n2[28] ,n2[92]);
    xnor g199(n2414 ,n995 ,n1084);
    nand g200(n2046 ,n10[4] ,n2031);
    nand g201(n2037 ,n10[10] ,n2031);
    nand g202(n1898 ,n1524 ,n1698);
    xnor g203(n2540 ,n2066 ,n2541);
    nand g204(n608 ,n370 ,n607);
    xnor g205(n2552 ,n2553 ,n2076);
    nor g206(n1012 ,n924 ,n1011);
    not g207(n1143 ,n10[4]);
    dff g208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1855), .Q(n7[13]));
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1851), .Q(n7[17]));
    nand g210(n1869 ,n1460 ,n1669);
    nand g211(n358 ,n2240 ,n11[45]);
    nand g212(n564 ,n329 ,n563);
    nand g213(n11[46] ,n2072 ,n2075);
    xnor g214(n4[62] ,n2113 ,n8[62]);
    or g215(n1249 ,n7[9] ,n1185);
    nand g216(n251 ,n24 ,n250);
    not g217(n1180 ,n1179);
    xnor g218(n5[58] ,n2101 ,n6[58]);
    not g219(n2065 ,n9[52]);
    nor g220(n1091 ,n973 ,n1090);
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1858), .Q(n7[11]));
    nand g222(n286 ,n118 ,n285);
    xnor g223(n2290 ,n142 ,n282);
    or g224(n26 ,n2339 ,n11[31]);
    nand g225(n1603 ,n2296 ,n1289);
    not g226(n2072 ,n9[47]);
    xnor g227(n471 ,n11[43] ,n2238);
    nor g228(n632 ,n2[16] ,n2[80]);
    not g229(n1294 ,n1293);
    nand g230(n1432 ,n2268 ,n1289);
    nand g231(n1631 ,n1216 ,n1493);
    xnor g232(n143 ,n11[31] ,n2355);
    nor g233(n1040 ,n888 ,n1039);
    nor g234(n1487 ,n1165 ,n1291);
    xnor g235(n951 ,n11[41] ,n2486);
    or g236(n1395 ,n8[32] ,n1292);
    or g237(n55 ,n2343 ,n11[35]);
    nand g238(n1945 ,n1568 ,n1743);
    nand g239(n1458 ,n2247 ,n1289);
    or g240(n1283 ,n6[41] ,n1185);
    or g241(n1239 ,n8[1] ,n1190);
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1907), .Q(n8[50]));
    xnor g243(n2527 ,n692 ,n843);
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1884), .Q(n6[52]));
    nand g245(n1744 ,n1345 ,n1501);
    xnor g246(n2465 ,n737 ,n781);
    nor g247(n1009 ,n966 ,n1008);
    xnor g248(n2320 ,n2079 ,n2[12]);
    nand g249(n1615 ,n2396 ,n1289);
    or g250(n1226 ,n6[35] ,n1199);
    nand g251(n341 ,n2185 ,n11[38]);
    nand g252(n213 ,n19 ,n212);
    or g253(n1372 ,n7[54] ,n1197);
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1826), .Q(n7[36]));
    nand g255(n539 ,n486 ,n538);
    nand g256(n1917 ,n1520 ,n1716);
    xnor g257(n4[27] ,n2105 ,n8[27]);
    xnor g258(n2536 ,n2078 ,n2537);
    nand g259(n1680 ,n1272 ,n1488);
    nand g260(n1777 ,n1326 ,n1501);
    nand g261(n264 ,n126 ,n263);
    nor g262(n1401 ,n1200 ,n1201);
    nand g263(n1608 ,n2382 ,n1289);
    xnor g264(n5[24] ,n2108 ,n6[24]);
    xnor g265(n2220 ,n2[104] ,n2070);
    nand g266(n2023 ,n9[54] ,n1914);
    nand g267(n604 ,n354 ,n603);
    nor g268(n681 ,n2[60] ,n2[124]);
    nor g269(n1146 ,n10[12] ,n10[13]);
    not g270(n1132 ,n10[1]);
    nand g271(n133 ,n2308 ,n9[49]);
    nand g272(n1985 ,n1420 ,n1781);
    not g273(n488 ,n487);
    nand g274(n330 ,n2214 ,n11[35]);
    xnor g275(n2128 ,n524 ,n453);
    xnor g276(n2392 ,n999 ,n1040);
    nor g277(n759 ,n683 ,n758);
    nand g278(n581 ,n462 ,n580);
    xnor g279(n141 ,n11[44] ,n2320);
    nand g280(n1607 ,n2383 ,n1289);
    nand g281(n562 ,n327 ,n561);
    nand g282(n1668 ,n1257 ,n1491);
    or g283(n51 ,n2310 ,n11[34]);
    nor g284(n663 ,n2[19] ,n2[83]);
    nor g285(n765 ,n639 ,n764);
    nand g286(n2014 ,n9[47] ,n1914);
    xnor g287(n971 ,n2446 ,n11[37]);
    nand g288(n322 ,n2204 ,n11[41]);
    nand g289(n1156 ,n13[1] ,n1129);
    nand g290(n587 ,n490 ,n586);
    or g291(n1373 ,n6[12] ,n1187);
    xnor g292(n2334 ,n2077 ,n2[26]);
    xnor g293(n4[15] ,n2115 ,n8[15]);
    nor g294(n1050 ,n905 ,n1049);
    nand g295(n572 ,n340 ,n571);
    xnor g296(n2221 ,n2[105] ,n2071);
    dff g297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1968), .Q(n8[10]));
    nand g298(n1456 ,n2119 ,n1289);
    xnor g299(n2213 ,n2[97] ,n2073);
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1872), .Q(n6[62]));
    nand g301(n1462 ,n2435 ,n1289);
    nand g302(n280 ,n99 ,n279);
    nand g303(n522 ,n352 ,n521);
    nor g304(n1066 ,n893 ,n1065);
    nor g305(n858 ,n744 ,n857);
    or g306(n1361 ,n8[28] ,n1187);
    or g307(n1281 ,n6[40] ,n1195);
    nand g308(n1406 ,n2380 ,n1289);
    nand g309(n1795 ,n1374 ,n1488);
    dff g310(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[12]), .Q(n9[60]));
    nand g311(n543 ,n492 ,n542);
    xnor g312(n2397 ,n972 ,n1050);
    nor g313(n1149 ,n10[8] ,n10[9]);
    nor g314(n650 ,n2[13] ,n2[77]);
    nand g315(n1658 ,n1244 ,n1499);
    xnor g316(n974 ,n11[37] ,n2478);
    xnor g317(n2210 ,n2[94] ,n2064);
    nand g318(n607 ,n482 ,n606);
    nand g319(n1402 ,n2419 ,n1289);
    xnor g320(n2510 ,n2069 ,n2511);
    nand g321(n11[39] ,n2070 ,n2069);
    nor g322(n661 ,n2[18] ,n2[82]);
    dff g323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2050), .Q(n10[13]));
    nand g324(n1599 ,n2146 ,n1289);
    nand g325(n1935 ,n1541 ,n1733);
    nor g326(n1491 ,n1159 ,n1291);
    nand g327(n97 ,n2356 ,n11[32]);
    xnor g328(n2468 ,n2073 ,n2469);
    or g329(n57 ,n2328 ,n11[36]);
    dff g330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1945), .Q(n8[24]));
    xnor g331(n5[25] ,n2111 ,n6[25]);
    nand g332(n1801 ,n1399 ,n1494);
    or g333(n1211 ,n7[36] ,n1196);
    xnor g334(n998 ,n11[42] ,n2520);
    dff g335(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1870), .Q(n7[0]));
    dff g336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1956), .Q(n8[17]));
    xnor g337(n691 ,n2[29] ,n2[93]);
    nor g338(n1049 ,n958 ,n1048);
    nand g339(n508 ,n338 ,n507);
    nand g340(n1702 ,n1297 ,n1488);
    nand g341(n1707 ,n1303 ,n1491);
    or g342(n1334 ,n8[20] ,n1196);
    or g343(n1247 ,n8[45] ,n1188);
    or g344(n1284 ,n8[52] ,n1196);
    nand g345(n109 ,n2320 ,n11[44]);
    xnor g346(n2239 ,n2[123] ,n2076);
    nor g347(n641 ,n2[8] ,n2[72]);
    xnor g348(n2352 ,n2079 ,n2[44]);
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1908), .Q(n6[40]));
    nand g350(n247 ,n74 ,n246);
    nand g351(n1957 ,n1528 ,n1755);
    nand g352(n1725 ,n1205 ,n1488);
    nand g353(n282 ,n105 ,n281);
    xnor g354(n397 ,n11[45] ,n2208);
    or g355(n1379 ,n8[29] ,n1188);
    xnor g356(n2296 ,n168 ,n294);
    nand g357(n298 ,n106 ,n297);
    xnor g358(n3[7] ,n2106 ,n7[7]);
    nand g359(n309 ,n25 ,n308);
    nor g360(n644 ,n2[50] ,n2[114]);
    xnor g361(n2415 ,n998 ,n1086);
    xnor g362(n479 ,n11[35] ,n2198);
    xnor g363(n4[32] ,n2107 ,n8[32]);
    nand g364(n1447 ,n2255 ,n1289);
    not g365(n438 ,n437);
    xnor g366(n2149 ,n566 ,n419);
    nand g367(n1539 ,n2300 ,n1289);
    nand g368(n1543 ,n2178 ,n1289);
    xnor g369(n996 ,n2470 ,n11[33]);
    nand g370(n619 ,n404 ,n618);
    xor g371(n2374 ,n941 ,n939);
    nand g372(n1844 ,n1430 ,n1645);
    xnor g373(n5[23] ,n2106 ,n6[23]);
    not g374(n2069 ,n9[54]);
    nand g375(n239 ,n46 ,n238);
    nand g376(n1642 ,n1231 ,n1491);
    nand g377(n613 ,n442 ,n612);
    nor g378(n893 ,n2498 ,n11[31]);
    or g379(n1223 ,n7[41] ,n1185);
    xnor g380(n3[0] ,n2098 ,n7[0]);
    xor g381(n2566 ,n2565 ,n2564);
    xnor g382(n173 ,n11[39] ,n2363);
    dff g383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1925), .Q(n6[34]));
    nand g384(n1745 ,n1343 ,n1500);
    dff g385(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1989), .Q(n7[59]));
    nand g386(n534 ,n365 ,n533);
    nand g387(n1636 ,n1258 ,n1499);
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1861), .Q(n7[8]));
    dff g389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2003), .Q(n7[49]));
    nand g390(n214 ,n44 ,n213);
    xnor g391(n970 ,n11[34] ,n2536);
    or g392(n1389 ,n7[32] ,n1292);
    nand g393(n117 ,n2339 ,n11[31]);
    nand g394(n1621 ,n1207 ,n1500);
    or g395(n1340 ,n8[22] ,n1197);
    or g396(n1301 ,n8[54] ,n1197);
    or g397(n1263 ,n6[62] ,n1192);
    xnor g398(n2528 ,n2072 ,n2529);
    nor g399(n1162 ,n9[52] ,n1155);
    nand g400(n2007 ,n1613 ,n1805);
    dff g401(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1990), .Q(n7[58]));
    xnor g402(n5[18] ,n2110 ,n6[18]);
    nor g403(n831 ,n654 ,n830);
    xnor g404(n461 ,n11[41] ,n2220);
    nor g405(n1079 ,n982 ,n1078);
    nand g406(n1423 ,n2272 ,n1289);
    nand g407(n1536 ,n2150 ,n1289);
    nand g408(n1451 ,n2161 ,n1289);
    xnor g409(n2503 ,n718 ,n819);
    nand g410(n203 ,n17 ,n202);
    xnor g411(n415 ,n11[40] ,n2235);
    nand g412(n1703 ,n1300 ,n1496);
    nand g413(n1859 ,n1448 ,n1660);
    dff g414(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2052), .Q(n10[11]));
    or g415(n756 ,n712 ,n755);
    xnor g416(n429 ,n11[40] ,n2203);
    xnor g417(n4[31] ,n2115 ,n8[31]);
    xnor g418(n166 ,n11[34] ,n2358);
    xnor g419(n4[9] ,n2111 ,n8[9]);
    xnor g420(n2241 ,n2[125] ,n2075);
    xnor g421(n961 ,n11[33] ,n2502);
    not g422(n452 ,n451);
    nor g423(n813 ,n685 ,n812);
    xnor g424(n2190 ,n2[74] ,n2077);
    nand g425(n1753 ,n1329 ,n1491);
    xnor g426(n2268 ,n183 ,n238);
    nand g427(n1682 ,n1278 ,n1500);
    dff g428(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2057), .Q(n10[7]));
    nand g429(n1871 ,n1462 ,n1671);
    nand g430(n1619 ,n1223 ,n1486);
    not g431(n428 ,n427);
    xnor g432(n2175 ,n618 ,n403);
    or g433(n1209 ,n7[37] ,n1191);
    xnor g434(n3[3] ,n2112 ,n7[3]);
    nand g435(n200 ,n94 ,n199);
    dff g436(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1991), .Q(n7[57]));
    nor g437(n1492 ,n1160 ,n1291);
    or g438(n1007 ,n963 ,n1006);
    nand g439(n1865 ,n1454 ,n1665);
    nand g440(n1687 ,n1394 ,n1494);
    nor g441(n762 ,n720 ,n761);
    xnor g442(n2534 ,n2535 ,n2068);
    xnor g443(n2136 ,n540 ,n487);
    nand g444(n541 ,n488 ,n540);
    nor g445(n1119 ,n1002 ,n1118);
    nor g446(n1019 ,n978 ,n1018);
    nor g447(n921 ,n2522 ,n11[43]);
    xnor g448(n2298 ,n172 ,n298);
    nand g449(n1519 ,n2163 ,n1289);
    xnor g450(n716 ,n2[59] ,n2[123]);
    nand g451(n2056 ,n2024 ,n2047);
    xnor g452(n2428 ,n991 ,n1112);
    or g453(n1366 ,n7[57] ,n1185);
    dff g454(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1950), .Q(n8[21]));
    nor g455(n830 ,n736 ,n829);
    xnor g456(n991 ,n11[39] ,n2546);
    xnor g457(n2367 ,n2076 ,n2[59]);
    xnor g458(n5[34] ,n2110 ,n6[34]);
    xnor g459(n485 ,n11[36] ,n2199);
    nand g460(n83 ,n2349 ,n11[41]);
    nand g461(n2039 ,n10[8] ,n2031);
    not g462(n1139 ,n10[14]);
    xnor g463(n2507 ,n724 ,n823);
    or g464(n1151 ,n13[0] ,n13[2]);
    xnor g465(n2487 ,n698 ,n803);
    xnor g466(n2233 ,n2[117] ,n2066);
    nor g467(n917 ,n2540 ,n11[36]);
    nor g468(n1024 ,n914 ,n1023);
    dff g469(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1967), .Q(n6[19]));
    nand g470(n598 ,n319 ,n597);
    xnor g471(n704 ,n2[32] ,n2[96]);
    dff g472(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1963), .Q(n6[22]));
    nand g473(n1956 ,n1560 ,n1754);
    or g474(n1246 ,n6[3] ,n1199);
    xnor g475(n2423 ,n970 ,n1102);
    nor g476(n782 ,n737 ,n781);
    not g477(n1138 ,n10[12]);
    dff g478(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1958), .Q(n8[15]));
    nand g479(n1420 ,n2387 ,n1289);
    or g480(n35 ,n2313 ,n11[37]);
    xnor g481(n457 ,n11[46] ,n2193);
    xnor g482(n2294 ,n166 ,n290);
    nor g483(n1152 ,n10[14] ,n10[15]);
    or g484(n1307 ,n8[57] ,n1185);
    nor g485(n930 ,n2542 ,n11[37]);
    xnor g486(n2466 ,n2467 ,n2067);
    nand g487(n511 ,n434 ,n510);
    nor g488(n1117 ,n983 ,n1116);
    xnor g489(n2331 ,n2074 ,n2[23]);
    nand g490(n1749 ,n1331 ,n1486);
    xor g491(n2100 ,n9[52] ,n2096);
    xnor g492(n690 ,n2[63] ,n2[127]);
    xnor g493(n978 ,n2452 ,n11[40]);
    xnor g494(n5[21] ,n2102 ,n6[21]);
    nand g495(n222 ,n77 ,n221);
    nor g496(n890 ,n2494 ,n11[45]);
    nand g497(n1909 ,n1482 ,n1709);
    xnor g498(n697 ,n2[47] ,n2[111]);
    xnor g499(n2192 ,n2[76] ,n2079);
    or g500(n1214 ,n7[34] ,n1193);
    nand g501(n506 ,n361 ,n505);
    nand g502(n546 ,n377 ,n545);
    nor g503(n1497 ,n1158 ,n1291);
    nand g504(n1591 ,n2423 ,n1289);
    xnor g505(n441 ,n11[41] ,n2236);
    or g506(n894 ,n2438 ,n11[33]);
    dff g507(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2056), .Q(n10[5]));
    nand g508(n1722 ,n1305 ,n1500);
    xnor g509(n4[36] ,n2100 ,n8[36]);
    xnor g510(n5[20] ,n2100 ,n6[20]);
    not g511(n1128 ,n1290);
    nand g512(n1440 ,n2260 ,n1289);
    nand g513(n2028 ,n9[48] ,n1914);
    dff g514(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1934), .Q(n8[32]));
    xnor g515(n2454 ,n2455 ,n2077);
    nand g516(n2086 ,n10[1] ,n11[33]);
    nor g517(n820 ,n718 ,n819);
    xnor g518(n392 ,n11[35] ,n2182);
    xnor g519(n5[26] ,n2101 ,n6[26]);
    xnor g520(n188 ,n11[39] ,n2331);
    not g521(n414 ,n413);
    nor g522(n847 ,n627 ,n846);
    or g523(n1265 ,n6[39] ,n1189);
    xor g524(n2110 ,n9[50] ,n2084);
    dff g525(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2006), .Q(n7[46]));
    nor g526(n1489 ,n1173 ,n1291);
    xnor g527(n145 ,n11[46] ,n2322);
    xnor g528(n3[26] ,n2101 ,n7[26]);
    xnor g529(n439 ,n11[42] ,n2237);
    not g530(n450 ,n449);
    or g531(n1808 ,n12[1] ,n1502);
    or g532(n1302 ,n8[12] ,n1187);
    dff g533(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1892), .Q(n6[44]));
    nand g534(n515 ,n438 ,n514);
    dff g535(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1879), .Q(n6[56]));
    nor g536(n682 ,n2[56] ,n2[120]);
    xnor g537(n3[14] ,n2113 ,n7[14]);
    nand g538(n1759 ,n1321 ,n1487);
    nand g539(n561 ,n396 ,n560);
    nand g540(n591 ,n418 ,n590);
    dff g541(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1764), .Q(n12[1]));
    dff g542(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1902), .Q(n8[54]));
    nand g543(n1693 ,n1322 ,n1498);
    nand g544(n301 ,n27 ,n300);
    dff g545(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1889), .Q(n8[62]));
    nand g546(n270 ,n120 ,n269);
    dff g547(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1933), .Q(n8[33]));
    xnor g548(n4[49] ,n2114 ,n8[49]);
    nor g549(n1167 ,n9[60] ,n1155);
    xnor g550(n138 ,n11[44] ,n2352);
    nand g551(n1825 ,n1409 ,n1624);
    nor g552(n876 ,n706 ,n875);
    nor g553(n771 ,n658 ,n770);
    nand g554(n229 ,n37 ,n228);
    dff g555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1898), .Q(n8[56]));
    xor g556(n2439 ,n712 ,n755);
    nor g557(n859 ,n674 ,n858);
    xnor g558(n181 ,n11[42] ,n2366);
    xnor g559(n2188 ,n2[72] ,n2070);
    nand g560(n2034 ,n10[13] ,n2031);
    nor g561(n1166 ,n9[47] ,n1155);
    nand g562(n363 ,n2195 ,n11[32]);
    nand g563(n1478 ,n2151 ,n1289);
    or g564(n56 ,n2326 ,n11[34]);
    xnor g565(n987 ,n11[36] ,n2540);
    nand g566(n87 ,n2343 ,n11[35]);
    or g567(n49 ,n2329 ,n11[37]);
    xnor g568(n4[22] ,n2104 ,n8[22]);
    nand g569(n283 ,n43 ,n282);
    xnor g570(n3[8] ,n2108 ,n7[8]);
    nand g571(n1924 ,n1530 ,n1724);
    nand g572(n1986 ,n1589 ,n1785);
    dff g573(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2060), .Q(n10[3]));
    or g574(n1310 ,n8[58] ,n1198);
    nor g575(n649 ,n2[57] ,n2[121]);
    nand g576(n1468 ,n2430 ,n1289);
    or g577(n1328 ,n8[25] ,n1185);
    xnor g578(n2274 ,n134 ,n250);
    or g579(n1271 ,n6[31] ,n1194);
    nor g580(n1495 ,n1161 ,n1291);
    dff g581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1980), .Q(n8[1]));
    nand g582(n300 ,n112 ,n299);
    nand g583(n1465 ,n2164 ,n1289);
    dff g584(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1921), .Q(n8[40]));
    nand g585(n1409 ,n2281 ,n1289);
    nand g586(n329 ,n2211 ,n11[32]);
    nor g587(n1023 ,n981 ,n1022);
    nor g588(n1168 ,n9[61] ,n1155);
    nand g589(n202 ,n89 ,n201);
    or g590(n1235 ,n6[1] ,n1190);
    nand g591(n233 ,n49 ,n232);
    or g592(n39 ,n2350 ,n11[42]);
    nand g593(n369 ,n2222 ,n11[43]);
    xnor g594(n2407 ,n964 ,n1070);
    nand g595(n1852 ,n1440 ,n1653);
    nand g596(n1894 ,n1529 ,n1694);
    nand g597(n1944 ,n1548 ,n1742);
    dff g598(.RN(1'b1), .SN(n2567), .CK(n0), .D(n9[53]), .Q(n14[7]));
    nor g599(n647 ,n2[12] ,n2[76]);
    dff g600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1887), .Q(n6[47]));
    nor g601(n638 ,n2[5] ,n2[69]);
    nand g602(n279 ,n52 ,n278);
    nand g603(n1008 ,n936 ,n1007);
    xnor g604(n390 ,n11[39] ,n2186);
    xnor g605(n2425 ,n987 ,n1106);
    dff g606(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1969), .Q(n6[18]));
    xor g607(n2245 ,n178 ,n133);
    xnor g608(n3[41] ,n2111 ,n7[41]);
    xnor g609(n739 ,n2[52] ,n2[116]);
    xnor g610(n186 ,n11[34] ,n2326);
    xnor g611(n706 ,n2[62] ,n2[126]);
    nand g612(n1884 ,n1477 ,n1681);
    xnor g613(n2446 ,n2447 ,n2069);
    not g614(n400 ,n399);
    nand g615(n284 ,n113 ,n283);
    nand g616(n1592 ,n2303 ,n1289);
    xnor g617(n2530 ,n2531 ,n2067);
    xor g618(n2113 ,n9[62] ,n2082);
    nand g619(n1650 ,n1237 ,n1491);
    or g620(n1278 ,n6[55] ,n1189);
    nor g621(n1493 ,n1166 ,n1291);
    dff g622(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1995), .Q(n7[54]));
    nand g623(n1751 ,n1338 ,n1489);
    xnor g624(n2509 ,n727 ,n825);
    or g625(n1309 ,n8[43] ,n1186);
    nand g626(n1748 ,n1304 ,n1496);
    xnor g627(n992 ,n2466 ,n11[31]);
    xnor g628(n734 ,n2[13] ,n2[77]);
    xnor g629(n5[4] ,n2100 ,n6[4]);
    xnor g630(n2516 ,n2071 ,n2517);
    xnor g631(n719 ,n2[16] ,n2[80]);
    nand g632(n513 ,n391 ,n512);
    xnor g633(n136 ,n11[32] ,n2340);
    xnor g634(n171 ,n11[38] ,n2314);
    dff g635(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1952), .Q(n8[19]));
    nand g636(n1910 ,n1522 ,n1616);
    nor g637(n842 ,n694 ,n841);
    nor g638(n1158 ,n9[62] ,n1155);
    xnor g639(n746 ,n2[20] ,n2[84]);
    dff g640(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1942), .Q(n6[28]));
    nand g641(n626 ,n344 ,n625);
    xnor g642(n3[6] ,n2104 ,n7[6]);
    xnor g643(n2180 ,n2[64] ,n2067);
    or g644(n54 ,n2320 ,n11[44]);
    dff g645(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1998), .Q(n6[10]));
    nand g646(n1512 ,n2168 ,n1289);
    nand g647(n1640 ,n1225 ,n1486);
    xnor g648(n2409 ,n975 ,n1074);
    xnor g649(n177 ,n11[34] ,n2310);
    nand g650(n1582 ,n2389 ,n1289);
    or g651(n1343 ,n8[23] ,n1189);
    xnor g652(n984 ,n2458 ,n11[43]);
    nand g653(n1905 ,n1513 ,n1704);
    xnor g654(n3[58] ,n2101 ,n7[58]);
    xnor g655(n4[20] ,n2100 ,n8[20]);
    nor g656(n806 ,n695 ,n805);
    dff g657(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1891), .Q(n8[61]));
    xnor g658(n2410 ,n979 ,n1076);
    xnor g659(n4[50] ,n2110 ,n8[50]);
    dff g660(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1829), .Q(n7[34]));
    or g661(n1232 ,n7[21] ,n1191);
    nor g662(n1179 ,n13[1] ,n1155);
    nor g663(n1062 ,n890 ,n1061);
    dff g664(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[3]), .Q(n9[51]));
    nand g665(n75 ,n2346 ,n11[38]);
    nand g666(n259 ,n45 ,n258);
    nand g667(n244 ,n102 ,n243);
    nand g668(n1445 ,n2256 ,n1289);
    xnor g669(n2360 ,n2065 ,n2[52]);
    dff g670(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1852), .Q(n7[16]));
    xnor g671(n989 ,n2464 ,n11[46]);
    nand g672(n78 ,n2348 ,n11[40]);
    xnor g673(n731 ,n2[12] ,n2[76]);
    nand g674(n1425 ,n2376 ,n1289);
    xnor g675(n5[47] ,n2115 ,n6[47]);
    nand g676(n2024 ,n9[53] ,n1914);
    xnor g677(n4[58] ,n2101 ,n8[58]);
    nor g678(n1154 ,n10[4] ,n10[5]);
    nand g679(n262 ,n87 ,n261);
    nand g680(n1485 ,n2124 ,n1289);
    nand g681(n1576 ,n2123 ,n1289);
    not g682(n486 ,n485);
    xnor g683(n5[61] ,n2103 ,n6[61]);
    xnor g684(n2385 ,n1026 ,n985);
    nand g685(n1998 ,n1608 ,n1803);
    nor g686(n1109 ,n1000 ,n1108);
    xnor g687(n144 ,n11[32] ,n2356);
    xnor g688(n946 ,n11[45] ,n2558);
    or g689(n1216 ,n7[31] ,n1194);
    xnor g690(n956 ,n11[38] ,n2448);
    nand g691(n544 ,n376 ,n543);
    xnor g692(n3[16] ,n2107 ,n7[16]);
    nand g693(n1911 ,n1465 ,n1710);
    nand g694(n1419 ,n2275 ,n1289);
    nand g695(n114 ,n2337 ,n11[45]);
    nand g696(n1438 ,n2373 ,n1289);
    nor g697(n797 ,n673 ,n796);
    dff g698(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1926), .Q(n8[37]));
    nand g699(n1832 ,n1418 ,n1630);
    xnor g700(n2560 ,n2072 ,n2561);
    nand g701(n1741 ,n1327 ,n1496);
    nor g702(n655 ,n2[24] ,n2[88]);
    nand g703(n1975 ,n1579 ,n1772);
    nand g704(n2004 ,n1609 ,n1801);
    nor g705(n2031 ,n1 ,n1914);
    xnor g706(n4[8] ,n2108 ,n8[8]);
    nand g707(n1569 ,n2128 ,n1289);
    nand g708(n1929 ,n1478 ,n1728);
    nand g709(n1524 ,n2172 ,n1289);
    xnor g710(n5[40] ,n2108 ,n6[40]);
    nor g711(n642 ,n2[45] ,n2[109]);
    xnor g712(n2300 ,n174 ,n302);
    xnor g713(n401 ,n11[33] ,n2228);
    nor g714(n840 ,n700 ,n839);
    dff g715(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1845), .Q(n6[3]));
    not g716(n480 ,n479);
    nand g717(n198 ,n119 ,n197);
    xnor g718(n2391 ,n997 ,n1038);
    nand g719(n1953 ,n1558 ,n1753);
    nor g720(n810 ,n691 ,n809);
    or g721(n1261 ,n8[46] ,n1192);
    xnor g722(n2172 ,n612 ,n441);
    xnor g723(n2488 ,n2076 ,n2489);
    nor g724(n1045 ,n974 ,n1044);
    nor g725(n879 ,n2464 ,n11[46]);
    not g726(n436 ,n435);
    xnor g727(n393 ,n11[46] ,n2209);
    xnor g728(n2470 ,n2471 ,n2068);
    nand g729(n2015 ,n9[62] ,n1914);
    nor g730(n929 ,n2544 ,n11[38]);
    nand g731(n1701 ,n1301 ,n1487);
    dff g732(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1911), .Q(n8[48]));
    xnor g733(n187 ,n11[37] ,n2329);
    xnor g734(n2176 ,n620 ,n431);
    or g735(n1315 ,n8[14] ,n1192);
    nor g736(n1104 ,n918 ,n1103);
    xnor g737(n3[17] ,n2114 ,n7[17]);
    xnor g738(n1001 ,n11[36] ,n2476);
    nand g739(n1517 ,n2412 ,n1289);
    nand g740(n1967 ,n1574 ,n1769);
    nand g741(n1155 ,n13[0] ,n1145);
    dff g742(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2010), .Q(n8[46]));
    xnor g743(n2387 ,n1030 ,n989);
    xnor g744(n2271 ,n192 ,n244);
    xnor g745(n481 ,n11[38] ,n2233);
    nand g746(n1841 ,n1427 ,n1640);
    xnor g747(n2554 ,n2079 ,n2555);
    not g748(n494 ,n493);
    xnor g749(n2135 ,n538 ,n485);
    xnor g750(n162 ,n11[43] ,n2351);
    nand g751(n1771 ,n1351 ,n1491);
    xor g752(n2103 ,n9[61] ,n2093);
    dff g753(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[2]), .Q(n9[50]));
    nand g754(n602 ,n343 ,n601);
    xnor g755(n736 ,n2[39] ,n2[103]);
    xnor g756(n2204 ,n2[88] ,n2070);
    nand g757(n577 ,n448 ,n576);
    xnor g758(n3[15] ,n2115 ,n7[15]);
    nand g759(n2033 ,n10[14] ,n2031);
    nand g760(n77 ,n2323 ,n11[31]);
    nor g761(n819 ,n635 ,n818);
    xnor g762(n2324 ,n2067 ,n2[16]);
    dff g763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1951), .Q(n8[20]));
    xnor g764(n2194 ,n2[78] ,n2064);
    nand g765(n1429 ,n2267 ,n1289);
    xnor g766(n2301 ,n176 ,n304);
    nand g767(n1810 ,n1472 ,n1502);
    or g768(n1329 ,n8[18] ,n1193);
    xnor g769(n174 ,n11[40] ,n2364);
    nand g770(n1669 ,n1259 ,n1492);
    nand g771(n510 ,n339 ,n509);
    or g772(n1344 ,n8[11] ,n1186);
    dff g773(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2063), .Q(n10[4]));
    xnor g774(n150 ,n11[38] ,n2330);
    nor g775(n1083 ,n990 ,n1082);
    nand g776(n621 ,n432 ,n620);
    nand g777(n106 ,n2361 ,n11[37]);
    nand g778(n2093 ,n10[13] ,n11[45]);
    or g779(n1225 ,n7[25] ,n1185);
    nor g780(n1194 ,n1142 ,n1155);
    nand g781(n1665 ,n1254 ,n1488);
    nand g782(n1873 ,n1464 ,n1673);
    xnor g783(n4[38] ,n2104 ,n8[38]);
    not g784(n1157 ,n1156);
    nand g785(n227 ,n56 ,n226);
    not g786(n2068 ,n9[50]);
    nor g787(n1052 ,n926 ,n1051);
    xnor g788(n2424 ,n994 ,n1104);
    xnor g789(n4[39] ,n2106 ,n8[39]);
    nand g790(n1435 ,n2159 ,n1289);
    nor g791(n857 ,n660 ,n856);
    nand g792(n129 ,n2366 ,n11[42]);
    nand g793(n1822 ,n1407 ,n1621);
    nand g794(n1482 ,n2165 ,n1289);
    nor g795(n687 ,n2[59] ,n2[123]);
    nand g796(n1541 ,n2147 ,n1289);
    nor g797(n628 ,n2[29] ,n2[93]);
    nand g798(n1006 ,n894 ,n1005);
    xnor g799(n2538 ,n2065 ,n2539);
    xnor g800(n3[56] ,n2108 ,n7[56]);
    or g801(n21 ,n2360 ,n11[36]);
    nand g802(n11[35] ,n2065 ,n2068);
    xnor g803(n2539 ,n739 ,n855);
    xnor g804(n5[37] ,n2102 ,n6[37]);
    xnor g805(n2494 ,n2064 ,n2495);
    xnor g806(n721 ,n2[57] ,n2[121]);
    nor g807(n862 ,n749 ,n861);
    xnor g808(n4[0] ,n2098 ,n8[0]);
    nor g809(n1071 ,n964 ,n1070);
    nand g810(n1510 ,n2414 ,n1289);
    nor g811(n674 ,n2[53] ,n2[117]);
    nand g812(n1876 ,n1468 ,n1676);
    nor g813(n849 ,n633 ,n848);
    nand g814(n1439 ,n2261 ,n1289);
    nor g815(n1039 ,n997 ,n1038);
    xnor g816(n2337 ,n2075 ,n2[29]);
    nor g817(n1011 ,n967 ,n1010);
    xnor g818(n399 ,n11[32] ,n2211);
    nand g819(n1950 ,n1554 ,n1747);
    nor g820(n1197 ,n1144 ,n1155);
    or g821(n1279 ,n6[50] ,n1193);
    xnor g822(n2475 ,n746 ,n791);
    nand g823(n1563 ,n2131 ,n1289);
    xnor g824(n4[34] ,n2110 ,n8[34]);
    xnor g825(n149 ,n11[33] ,n2341);
    or g826(n1357 ,n8[2] ,n1193);
    nand g827(n574 ,n342 ,n573);
    nand g828(n1726 ,n1285 ,n1492);
    nand g829(n1520 ,n2409 ,n1289);
    xnor g830(n2366 ,n2077 ,n2[58]);
    nand g831(n1182 ,n1154 ,n1150);
    nand g832(n218 ,n132 ,n217);
    or g833(n1355 ,n8[4] ,n1196);
    xnor g834(n2353 ,n2075 ,n2[45]);
    nor g835(n906 ,n2538 ,n11[35]);
    nor g836(n889 ,n2528 ,n11[46]);
    or g837(n1333 ,n8[21] ,n1191);
    not g838(n2064 ,n9[62]);
    nand g839(n1556 ,n2397 ,n1289);
    xnor g840(n3[1] ,n2114 ,n7[1]);
    nand g841(n2051 ,n2030 ,n2039);
    nand g842(n1407 ,n2283 ,n1289);
    xnor g843(n2551 ,n738 ,n867);
    dff g844(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1831), .Q(n7[33]));
    xnor g845(n2248 ,n156 ,n198);
    xnor g846(n2473 ,n745 ,n789);
    nand g847(n552 ,n333 ,n551);
    nor g848(n770 ,n726 ,n769);
    nand g849(n1868 ,n1459 ,n1668);
    xnor g850(n2541 ,n744 ,n857);
    nand g851(n1547 ,n2142 ,n1289);
    dff g852(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1850), .Q(n7[18]));
    nand g853(n585 ,n476 ,n584);
    or g854(n1213 ,n6[6] ,n1197);
    nor g855(n1500 ,n1163 ,n1291);
    xnor g856(n2232 ,n2[116] ,n2065);
    xnor g857(n2405 ,n955 ,n1066);
    nand g858(n207 ,n58 ,n206);
    dff g859(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1875), .Q(n6[59]));
    not g860(n1140 ,n10[3]);
    nand g861(n273 ,n48 ,n272);
    nand g862(n1573 ,n2392 ,n1289);
    xnor g863(n2162 ,n592 ,n493);
    nor g864(n932 ,n2524 ,n11[44]);
    or g865(n1282 ,n8[36] ,n1196);
    xnor g866(n975 ,n11[36] ,n2508);
    xnor g867(n2499 ,n704 ,n815);
    nor g868(n640 ,n2[49] ,n2[113]);
    xnor g869(n749 ,n2[55] ,n2[119]);
    nor g870(n1400 ,n2372 ,n1128);
    nand g871(n130 ,n2318 ,n11[42]);
    nor g872(n1148 ,n10[2] ,n10[3]);
    nor g873(n659 ,n2[32] ,n2[96]);
    or g874(n1312 ,n8[40] ,n1195);
    xnor g875(n2408 ,n969 ,n1072);
    not g876(n496 ,n495);
    xnor g877(n4[48] ,n2107 ,n8[48]);
    xnor g878(n2479 ,n750 ,n795);
    nand g879(n624 ,n325 ,n623);
    xnor g880(n2251 ,n182 ,n204);
    xnor g881(n433 ,n11[38] ,n2185);
    dff g882(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1903), .Q(n8[53]));
    xnor g883(n752 ,n2[6] ,n2[70]);
    xnor g884(n747 ,n2[42] ,n2[106]);
    xnor g885(n5[7] ,n2106 ,n6[7]);
    nand g886(n1866 ,n1457 ,n1666);
    nand g887(n1862 ,n1455 ,n1664);
    nor g888(n1082 ,n911 ,n1081);
    nand g889(n1756 ,n1339 ,n1500);
    nand g890(n520 ,n350 ,n519);
    xnor g891(n5[17] ,n2114 ,n6[17]);
    nand g892(n1736 ,n1370 ,n1497);
    xnor g893(n2133 ,n534 ,n473);
    nand g894(n1601 ,n2297 ,n1289);
    nand g895(n100 ,n2333 ,n11[41]);
    or g896(n16 ,n2318 ,n11[42]);
    nand g897(n299 ,n68 ,n298);
    nand g898(n356 ,n2192 ,n11[45]);
    dff g899(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1982), .Q(n6[16]));
    nand g900(n2052 ,n2018 ,n2036);
    nand g901(n1555 ,n2136 ,n1289);
    nand g902(n195 ,n51 ,n194);
    nand g903(n11[38] ,n2074 ,n2066);
    or g904(n1299 ,n8[55] ,n1189);
    xnor g905(n5[14] ,n2113 ,n6[14]);
    nand g906(n1617 ,n1324 ,n1489);
    xnor g907(n4[46] ,n2113 ,n8[46]);
    nand g908(n339 ,n2184 ,n11[37]);
    nand g909(n1554 ,n2137 ,n1289);
    nor g910(n904 ,n2454 ,n11[41]);
    nor g911(n1188 ,n1136 ,n1155);
    xnor g912(n2168 ,n604 ,n459);
    xnor g913(n728 ,n2[10] ,n2[74]);
    dff g914(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1841), .Q(n7[25]));
    nand g915(n1015 ,n957 ,n1014);
    nand g916(n1857 ,n1438 ,n1644);
    not g917(n2073 ,n9[49]);
    nand g918(n348 ,n2180 ,n11[33]);
    or g919(n1250 ,n7[8] ,n1195);
    nand g920(n1937 ,n1542 ,n1736);
    xnor g921(n183 ,n11[40] ,n2332);
    nand g922(n199 ,n29 ,n198);
    nor g923(n1034 ,n910 ,n1033);
    xnor g924(n4[60] ,n2109 ,n8[60]);
    dff g925(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1966), .Q(n6[21]));
    nor g926(n778 ,n734 ,n777);
    nand g927(n623 ,n500 ,n622);
    or g928(n43 ,n2354 ,n11[46]);
    or g929(n335 ,n2181 ,n11[34]);
    nand g930(n1604 ,n2295 ,n1289);
    xnor g931(n2525 ,n694 ,n841);
    nand g932(n248 ,n110 ,n247);
    or g933(n1371 ,n6[57] ,n1185);
    nor g934(n684 ,n2[31] ,n2[95]);
    nand g935(n1005 ,n939 ,n942);
    nor g936(n633 ,n2[48] ,n2[112]);
    xor g937(n2244 ,n2308 ,n9[49]);
    xnor g938(n4[24] ,n2108 ,n8[24]);
    xnor g939(n3[54] ,n2104 ,n7[54]);
    dff g940(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2009), .Q(n8[45]));
    xnor g941(n2184 ,n2[68] ,n2065);
    xnor g942(n147 ,n11[44] ,n2336);
    dff g943(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1905), .Q(n6[41]));
    xnor g944(n2142 ,n552 ,n477);
    xnor g945(n4[12] ,n2109 ,n8[12]);
    nor g946(n919 ,n2470 ,n11[33]);
    nand g947(n1552 ,n2399 ,n1289);
    xnor g948(n733 ,n2[51] ,n2[115]);
    xnor g949(n2161 ,n590 ,n417);
    xnor g950(n469 ,n11[33] ,n2196);
    xnor g951(n167 ,n11[35] ,n2359);
    or g952(n40 ,n2355 ,n11[31]);
    xnor g953(n2267 ,n188 ,n236);
    nor g954(n1020 ,n933 ,n1019);
    nor g955(n1169 ,n9[48] ,n1155);
    nand g956(n2012 ,n1294 ,n1915);
    xnor g957(n2323 ,n2072 ,n2[15]);
    xnor g958(n2283 ,n158 ,n268);
    nor g959(n634 ,n2[15] ,n2[79]);
    xnor g960(n2328 ,n2065 ,n2[20]);
    not g961(n387 ,n386);
    nand g962(n1505 ,n2416 ,n1289);
    nand g963(n11[33] ,n2068 ,n2067);
    xnor g964(n5[16] ,n2107 ,n6[16]);
    nand g965(n357 ,n2193 ,n11[46]);
    nand g966(n2057 ,n2022 ,n2040);
    nand g967(n221 ,n34 ,n220);
    nor g968(n1065 ,n952 ,n1064);
    nand g969(n1824 ,n1406 ,n1617);
    xnor g970(n732 ,n2[38] ,n2[102]);
    nor g971(n1113 ,n991 ,n1112);
    dff g972(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1896), .Q(n6[45]));
    or g973(n1363 ,n6[14] ,n1192);
    nand g974(n11[43] ,n2079 ,n2077);
    xnor g975(n5[10] ,n2101 ,n6[10]);
    nor g976(n843 ,n642 ,n842);
    nand g977(n2091 ,n10[11] ,n11[43]);
    xnor g978(n2497 ,n699 ,n813);
    xnor g979(n5[33] ,n2114 ,n6[33]);
    nor g980(n1177 ,n13[2] ,n1156);
    xnor g981(n2193 ,n2[77] ,n2075);
    nand g982(n268 ,n75 ,n267);
    nor g983(n679 ,n2[27] ,n2[91]);
    dff g984(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1943), .Q(n8[26]));
    dff g985(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1913), .Q(n13[2]));
    xnor g986(n2249 ,n185 ,n200);
    xnor g987(n722 ,n2[48] ,n2[112]);
    xnor g988(n5[46] ,n2113 ,n6[46]);
    or g989(n1377 ,n7[50] ,n1193);
    nand g990(n1863 ,n1452 ,n1663);
    xnor g991(n154 ,n11[36] ,n2328);
    nor g992(n800 ,n702 ,n799);
    nand g993(n2092 ,n10[6] ,n11[38]);
    nand g994(n1594 ,n2302 ,n1289);
    nand g995(n1845 ,n1428 ,n1639);
    nor g996(n871 ,n687 ,n870);
    nand g997(n230 ,n85 ,n229);
    dff g998(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2001), .Q(n7[50]));
    nand g999(n293 ,n71 ,n292);
    xnor g1000(n4[26] ,n2101 ,n8[26]);
    xnor g1001(n2226 ,n2[110] ,n2064);
    nand g1002(n378 ,n2224 ,n11[45]);
    nand g1003(n1627 ,n1212 ,n1495);
    nand g1004(n2095 ,n10[10] ,n11[42]);
    nor g1005(n905 ,n2482 ,n11[39]);
    nor g1006(n822 ,n705 ,n821);
    or g1007(n1380 ,n8[30] ,n1192);
    nand g1008(n504 ,n335 ,n503);
    xor g1009(n2105 ,n9[59] ,n2091);
    dff g1010(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1946), .Q(n8[23]));
    xnor g1011(n2489 ,n695 ,n805);
    nor g1012(n1043 ,n1001 ,n1042);
    nand g1013(n1443 ,n2258 ,n1289);
    xnor g1014(n5[1] ,n2114 ,n6[1]);
    dff g1015(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1988), .Q(n7[60]));
    nand g1016(n1755 ,n1396 ,n1494);
    or g1017(n1349 ,n8[8] ,n1195);
    nand g1018(n1516 ,n2166 ,n1289);
    nand g1019(n1993 ,n1598 ,n1793);
    nand g1020(n1657 ,n1243 ,n1498);
    or g1021(n18 ,n2331 ,n11[39]);
    nor g1022(n678 ,n2[38] ,n2[102]);
    xnor g1023(n3[20] ,n2100 ,n7[20]);
    nand g1024(n1564 ,n2130 ,n1289);
    xnor g1025(n2565 ,n9[60] ,n14[15]);
    nand g1026(n1515 ,n2415 ,n1289);
    nand g1027(n2059 ,n2028 ,n2042);
    xnor g1028(n695 ,n2[27] ,n2[91]);
    dff g1029(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1927), .Q(n8[36]));
    nand g1030(n1612 ,n2290 ,n1289);
    xnor g1031(n2338 ,n2064 ,n2[30]);
    nand g1032(n1932 ,n1538 ,n1734);
    xnor g1033(n2517 ,n742 ,n833);
    xnor g1034(n990 ,n11[40] ,n2516);
    xnor g1035(n134 ,n11[46] ,n2338);
    nand g1036(n194 ,n121 ,n193);
    xnor g1037(n2126 ,n520 ,n445);
    xnor g1038(n2314 ,n2069 ,n2[6]);
    nor g1039(n935 ,n2442 ,n11[35]);
    nand g1040(n377 ,n2202 ,n11[39]);
    or g1041(n1297 ,n8[53] ,n1191);
    nor g1042(n788 ,n743 ,n787);
    nor g1043(n828 ,n732 ,n827);
    or g1044(n1388 ,n6[19] ,n1199);
    xnor g1045(n2208 ,n2[92] ,n2079);
    xnor g1046(n2419 ,n954 ,n1094);
    nand g1047(n1452 ,n2251 ,n1289);
    xnor g1048(n178 ,n11[33] ,n2309);
    xnor g1049(n4[57] ,n2111 ,n8[57]);
    xnor g1050(n2309 ,n2073 ,n2[1]);
    or g1051(n1280 ,n8[51] ,n1199);
    dff g1052(.RN(1'b1), .SN(n2567), .CK(n0), .D(n14[2]), .Q(n14[3]));
    xnor g1053(n146 ,n11[45] ,n2321);
    or g1054(n1304 ,n6[26] ,n1198);
    nand g1055(n373 ,n2227 ,n11[32]);
    xnor g1056(n2170 ,n608 ,n501);
    nand g1057(n1711 ,n1265 ,n1500);
    xnor g1058(n2459 ,n731 ,n775);
    xnor g1059(n2394 ,n974 ,n1044);
    or g1060(n1317 ,n6[34] ,n1193);
    xnor g1061(n2278 ,n151 ,n258);
    nor g1062(n829 ,n678 ,n828);
    xnor g1063(n2098 ,n2067 ,n2080);
    nand g1064(n1672 ,n1263 ,n1497);
    nand g1065(n1696 ,n1316 ,n1499);
    dff g1066(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2058), .Q(n10[6]));
    not g1067(n406 ,n405);
    xnor g1068(n2321 ,n2075 ,n2[13]);
    xnor g1069(n729 ,n2[61] ,n2[125]);
    nand g1070(n208 ,n82 ,n207);
    xnor g1071(n3[13] ,n2103 ,n7[13]);
    xnor g1072(n2284 ,n159 ,n270);
    nand g1073(n600 ,n320 ,n599);
    or g1074(n1335 ,n8[19] ,n1199);
    nand g1075(n1699 ,n1311 ,n1501);
    nand g1076(n609 ,n502 ,n608);
    not g1077(n402 ,n401);
    nor g1078(n1187 ,n1138 ,n1155);
    xnor g1079(n2523 ,n700 ,n839);
    nand g1080(n1908 ,n1517 ,n1708);
    not g1081(n454 ,n453);
    xnor g1082(n983 ,n11[41] ,n2550);
    nand g1083(n1678 ,n1318 ,n1487);
    nand g1084(n312 ,n2368 ,n310);
    xnor g1085(n741 ,n2[8] ,n2[72]);
    nand g1086(n1738 ,n1361 ,n1499);
    nand g1087(n1427 ,n2269 ,n1289);
    nor g1088(n673 ,n2[22] ,n2[86]);
    nand g1089(n1437 ,n2374 ,n1289);
    xnor g1090(n2379 ,n1014 ,n956);
    xnor g1091(n2480 ,n2481 ,n2074);
    nand g1092(n290 ,n127 ,n289);
    nor g1093(n1190 ,n1132 ,n1155);
    xnor g1094(n964 ,n11[34] ,n2504);
    nor g1095(n1075 ,n975 ,n1074);
    nand g1096(n2006 ,n1612 ,n1804);
    nor g1097(n1077 ,n979 ,n1076);
    nand g1098(n223 ,n60 ,n222);
    xnor g1099(n3[47] ,n2115 ,n7[47]);
    dff g1100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1986), .Q(n7[61]));
    nor g1101(n1030 ,n913 ,n1029);
    or g1102(n1327 ,n8[26] ,n1198);
    nand g1103(n1587 ,n2307 ,n1289);
    nand g1104(n509 ,n389 ,n508);
    xnor g1105(n2432 ,n944 ,n1120);
    not g1106(n426 ,n425);
    xnor g1107(n427 ,n11[36] ,n2215);
    nand g1108(n535 ,n474 ,n534);
    xnor g1109(n139 ,n11[31] ,n2323);
    nor g1110(n918 ,n2536 ,n11[34]);
    nand g1111(n265 ,n72 ,n264);
    xnor g1112(n5[63] ,n2099 ,n6[63]);
    xnor g1113(n4[5] ,n2102 ,n8[5]);
    xnor g1114(n495 ,n11[45] ,n2224);
    nor g1115(n1126 ,n902 ,n1125);
    nor g1116(n786 ,n740 ,n785);
    nand g1117(n530 ,n359 ,n529);
    not g1118(n1130 ,n10[9]);
    or g1119(n72 ,n2345 ,n11[37]);
    xnor g1120(n5[56] ,n2108 ,n6[56]);
    xnor g1121(n5[12] ,n2109 ,n6[12]);
    dff g1122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1838), .Q(n7[27]));
    nand g1123(n263 ,n38 ,n262);
    xnor g1124(n955 ,n2500 ,n11[32]);
    xnor g1125(n4[10] ,n2101 ,n8[10]);
    nand g1126(n939 ,n2436 ,n9[49]);
    nand g1127(n1990 ,n1594 ,n1788);
    nand g1128(n337 ,n2236 ,n11[41]);
    nand g1129(n102 ,n2334 ,n11[42]);
    not g1130(n1134 ,n10[11]);
    nand g1131(n1645 ,n1224 ,n1487);
    nand g1132(n292 ,n104 ,n291);
    xnor g1133(n2157 ,n582 ,n467);
    nand g1134(n612 ,n362 ,n611);
    or g1135(n505 ,n392 ,n504);
    nand g1136(n2002 ,n1602 ,n1792);
    nand g1137(n206 ,n125 ,n205);
    xnor g1138(n2132 ,n532 ,n469);
    dff g1139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1822), .Q(n7[39]));
    xnor g1140(n2377 ,n1010 ,n967);
    nand g1141(n1705 ,n1284 ,n1490);
    nand g1142(n1565 ,n2129 ,n1289);
    xnor g1143(n2310 ,n2068 ,n2[2]);
    xnor g1144(n499 ,n11[46] ,n2241);
    xnor g1145(n737 ,n2[15] ,n2[79]);
    nand g1146(n1867 ,n1458 ,n1667);
    nor g1147(n2304 ,n313 ,n311);
    nor g1148(n653 ,n2[61] ,n2[125]);
    nand g1149(n1890 ,n1503 ,n1691);
    xnor g1150(n2145 ,n558 ,n393);
    xnor g1151(n2240 ,n2[124] ,n2079);
    not g1152(n977 ,n976);
    xnor g1153(n2189 ,n2[73] ,n2071);
    or g1154(n1251 ,n8[35] ,n1199);
    nand g1155(n576 ,n331 ,n575);
    dff g1156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1978), .Q(n6[17]));
    nand g1157(n1787 ,n1364 ,n1501);
    xnor g1158(n156 ,n11[36] ,n2312);
    nand g1159(n2044 ,n10[1] ,n2031);
    dff g1160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1860), .Q(n7[9]));
    xnor g1161(n742 ,n2[41] ,n2[105]);
    dff g1162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2048), .Q(n10[15]));
    dff g1163(.RN(1'b1), .SN(n2567), .CK(n0), .D(n2566), .Q(n14[0]));
    nand g1164(n308 ,n129 ,n307);
    nand g1165(n128 ,n2324 ,n11[32]);
    xnor g1166(n2545 ,n749 ,n861);
    nand g1167(n1948 ,n1553 ,n1748);
    xnor g1168(n2171 ,n610 ,n415);
    xnor g1169(n4[51] ,n2112 ,n8[51]);
    nand g1170(n95 ,n2360 ,n11[36]);
    nand g1171(n578 ,n353 ,n577);
    nand g1172(n1578 ,n2122 ,n1289);
    nand g1173(n1836 ,n1422 ,n1635);
    nand g1174(n1647 ,n1234 ,n1490);
    nor g1175(n646 ,n2[37] ,n2[101]);
    nor g1176(n1067 ,n955 ,n1066);
    nand g1177(n2061 ,n2029 ,n2043);
    dff g1178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1987), .Q(n6[14]));
    xnor g1179(n2329 ,n2066 ,n2[21]);
    nand g1180(n1620 ,n1206 ,n1489);
    nand g1181(n110 ,n2336 ,n11[44]);
    xnor g1182(n2562 ,n12[2] ,n1127);
    xnor g1183(n724 ,n2[36] ,n2[100]);
    xnor g1184(n2155 ,n578 ,n455);
    nor g1185(n1108 ,n917 ,n1107);
    nand g1186(n1581 ,n2120 ,n1289);
    xnor g1187(n140 ,n11[45] ,n2353);
    nor g1188(n1189 ,n1135 ,n1155);
    nor g1189(n1098 ,n899 ,n1097);
    not g1190(n1815 ,n1811);
    xnor g1191(n3[43] ,n2105 ,n7[43]);
    nand g1192(n1716 ,n1240 ,n1488);
    xnor g1193(n190 ,n11[41] ,n2333);
    xnor g1194(n3[39] ,n2106 ,n7[39]);
    xnor g1195(n182 ,n11[39] ,n2315);
    xnor g1196(n701 ,n2[54] ,n2[118]);
    or g1197(n28 ,n2358 ,n11[34]);
    nand g1198(n1675 ,n1267 ,n1501);
    or g1199(n45 ,n2342 ,n11[34]);
    nand g1200(n1639 ,n1246 ,n1495);
    xnor g1201(n2413 ,n990 ,n1082);
    nand g1202(n1613 ,n2289 ,n1289);
    dff g1203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1961), .Q(n8[14]));
    xnor g1204(n487 ,n11[37] ,n2200);
    xnor g1205(n5[30] ,n2113 ,n6[30]);
    nand g1206(n1568 ,n2140 ,n1289);
    dff g1207(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[15]), .Q(n9[47]));
    nand g1208(n2087 ,n10[8] ,n11[40]);
    xnor g1209(n463 ,n11[31] ,n2194);
    xnor g1210(n715 ,n2[3] ,n2[67]);
    nor g1211(n1165 ,n9[54] ,n1155);
    xnor g1212(n2435 ,n940 ,n1126);
    nand g1213(n2010 ,n1453 ,n1713);
    dff g1214(.RN(n2567), .SN(1'b1), .CK(n0), .D(n9[51]), .Q(n9[52]));
    nor g1215(n900 ,n2508 ,n11[36]);
    nand g1216(n1586 ,n2116 ,n1289);
    xnor g1217(n949 ,n2530 ,n11[31]);
    nand g1218(n285 ,n40 ,n284);
    nor g1219(n1029 ,n988 ,n1028);
    not g1220(n2075 ,n9[61]);
    nor g1221(n1914 ,n12[2] ,n1808);
    nand g1222(n101 ,n2310 ,n11[34]);
    nor g1223(n658 ,n2[9] ,n2[73]);
    xnor g1224(n3[38] ,n2104 ,n7[38]);
    nand g1225(n367 ,n2197 ,n11[34]);
    or g1226(n1234 ,n7[20] ,n1196);
    xnor g1227(n5[28] ,n2109 ,n6[28]);
    xnor g1228(n2325 ,n2073 ,n2[17]);
    nand g1229(n1960 ,n1567 ,n1687);
    or g1230(n74 ,n2336 ,n11[44]);
    xnor g1231(n388 ,n11[37] ,n2184);
    dff g1232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1917), .Q(n6[37]));
    nor g1233(n896 ,n2554 ,n11[43]);
    nor g1234(n798 ,n753 ,n797);
    xnor g1235(n191 ,n11[42] ,n2334);
    xnor g1236(n2292 ,n144 ,n286);
    nand g1237(n1839 ,n1426 ,n1638);
    nor g1238(n1054 ,n934 ,n1053);
    xnor g1239(n2234 ,n2[118] ,n2069);
    nor g1240(n672 ,n2[46] ,n2[110]);
    xnor g1241(n2376 ,n1008 ,n966);
    nand g1242(n1906 ,n1484 ,n1706);
    nor g1243(n1055 ,n959 ,n1054);
    nor g1244(n1486 ,n1172 ,n1291);
    xnor g1245(n2356 ,n2067 ,n2[48]);
    nand g1246(n108 ,n2365 ,n11[41]);
    nand g1247(n1982 ,n1585 ,n1776);
    or g1248(n65 ,n2311 ,n11[35]);
    nor g1249(n804 ,n698 ,n803);
    nand g1250(n548 ,n332 ,n547);
    or g1251(n70 ,n2340 ,n11[32]);
    nand g1252(n1995 ,n1600 ,n1794);
    nand g1253(n1414 ,n2278 ,n1289);
    or g1254(n1300 ,n6[42] ,n1198);
    nand g1255(n1575 ,n2390 ,n1289);
    xnor g1256(n2461 ,n734 ,n777);
    xnor g1257(n997 ,n11[34] ,n2472);
    nor g1258(n1068 ,n892 ,n1067);
    xnor g1259(n2312 ,n2065 ,n2[4]);
    xnor g1260(n2250 ,n171 ,n202);
    or g1261(n1313 ,n7[38] ,n1197);
    xnor g1262(n2223 ,n2[107] ,n2076);
    nand g1263(n1681 ,n1275 ,n1490);
    nor g1264(n675 ,n2[43] ,n2[107]);
    nand g1265(n216 ,n109 ,n215);
    xnor g1266(n2350 ,n2077 ,n2[42]);
    nand g1267(n1453 ,n2162 ,n1289);
    xnor g1268(n5[50] ,n2110 ,n6[50]);
    xnor g1269(n2282 ,n157 ,n266);
    dff g1270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1816), .Q(n6[39]));
    nand g1271(n1747 ,n1333 ,n1488);
    or g1272(n1352 ,n7[47] ,n1194);
    xnor g1273(n137 ,n11[32] ,n2324);
    xnor g1274(n5[31] ,n2115 ,n6[31]);
    or g1275(n1305 ,n8[39] ,n1189);
    dff g1276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1955), .Q(n6[24]));
    nor g1277(n848 ,n722 ,n847);
    xnor g1278(n988 ,n2462 ,n11[45]);
    nand g1279(n1835 ,n1480 ,n1632);
    xnor g1280(n2259 ,n139 ,n220);
    nand g1281(n1540 ,n2148 ,n1289);
    nand g1282(n1724 ,n1208 ,n1487);
    nand g1283(n1899 ,n1514 ,n1700);
    dff g1284(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1839), .Q(n7[26]));
    nand g1285(n1752 ,n1335 ,n1495);
    nand g1286(n11[40] ,n2071 ,n2074);
    xor g1287(n2104 ,n9[54] ,n2092);
    nand g1288(n1926 ,n1532 ,n1725);
    nand g1289(n1776 ,n1397 ,n1494);
    or g1290(n66 ,n2322 ,n11[46]);
    xnor g1291(n2518 ,n2077 ,n2519);
    dff g1292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1924), .Q(n8[38]));
    nand g1293(n755 ,n631 ,n754);
    xnor g1294(n2417 ,n973 ,n1090);
    nand g1295(n1947 ,n1552 ,n1744);
    nand g1296(n287 ,n31 ,n286);
    nand g1297(n2084 ,n10[2] ,n11[34]);
    nand g1298(n1847 ,n1437 ,n1642);
    xnor g1299(n435 ,n11[37] ,n2216);
    nand g1300(n302 ,n122 ,n301);
    xnor g1301(n5[19] ,n2112 ,n6[19]);
    xnor g1302(n2464 ,n2072 ,n2465);
    nand g1303(n354 ,n2231 ,n11[36]);
    dff g1304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1883), .Q(n6[50]));
    nand g1305(n1994 ,n1597 ,n1791);
    xnor g1306(n2156 ,n580 ,n461);
    xnor g1307(n2273 ,n148 ,n248);
    nand g1308(n1813 ,n1347 ,n1490);
    nor g1309(n794 ,n748 ,n793);
    or g1310(n1367 ,n8[62] ,n1192);
    xnor g1311(n2411 ,n982 ,n1078);
    nand g1312(n1424 ,n2271 ,n1289);
    nand g1313(n372 ,n2223 ,n11[44]);
    nand g1314(n116 ,n2338 ,n11[46]);
    xnor g1315(n2456 ,n2076 ,n2457);
    xnor g1316(n699 ,n2[31] ,n2[95]);
    dff g1317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1938), .Q(n8[29]));
    nand g1318(n1677 ,n1371 ,n1486);
    nand g1319(n1504 ,n2417 ,n1289);
    xnor g1320(n2526 ,n2064 ,n2527);
    dff g1321(.RN(1'b1), .SN(n2567), .CK(n0), .D(n14[14]), .Q(n14[15]));
    xnor g1322(n3[63] ,n2099 ,n7[63]);
    nor g1323(n1290 ,n1 ,n1180);
    nand g1324(n1626 ,n1211 ,n1490);
    nand g1325(n1709 ,n1277 ,n1492);
    or g1326(n1350 ,n8[7] ,n1189);
    nand g1327(n1850 ,n1436 ,n1650);
    xnor g1328(n2123 ,n514 ,n437);
    dff g1329(.RN(1'b1), .SN(n2567), .CK(n0), .D(n14[9]), .Q(n14[10]));
    nand g1330(n1730 ,n1320 ,n1492);
    nand g1331(n2045 ,n10[3] ,n2031);
    or g1332(n1288 ,n8[59] ,n1186);
    nand g1333(n1877 ,n1610 ,n1677);
    xnor g1334(n982 ,n11[38] ,n2512);
    nor g1335(n772 ,n728 ,n771);
    nand g1336(n1464 ,n2433 ,n1289);
    nand g1337(n1514 ,n2171 ,n1289);
    dff g1338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1840), .Q(n6[4]));
    nor g1339(n926 ,n2484 ,n11[40]);
    nor g1340(n1115 ,n953 ,n1114);
    nand g1341(n1828 ,n1412 ,n1627);
    dff g1342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1867), .Q(n7[3]));
    or g1343(n1217 ,n6[29] ,n1188);
    xnor g1344(n2181 ,n2[65] ,n2073);
    nand g1345(n1663 ,n1252 ,n1500);
    nand g1346(n1634 ,n1219 ,n1490);
    nand g1347(n2011 ,n1565 ,n1760);
    or g1348(n1320 ,n8[33] ,n1190);
    xnor g1349(n3[50] ,n2110 ,n7[50]);
    xnor g1350(n161 ,n11[42] ,n2350);
    nand g1351(n220 ,n76 ,n219);
    dff g1352(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1906), .Q(n8[51]));
    nand g1353(n355 ,n2191 ,n11[44]);
    nand g1354(n364 ,n2232 ,n11[37]);
    dff g1355(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1847), .Q(n6[2]));
    nand g1356(n1723 ,n1317 ,n1491);
    nand g1357(n1595 ,n2301 ,n1289);
    nand g1358(n288 ,n97 ,n287);
    xnor g1359(n4[40] ,n2108 ,n8[40]);
    xnor g1360(n727 ,n2[37] ,n2[101]);
    nand g1361(n936 ,n2440 ,n11[34]);
    nand g1362(n1770 ,n1286 ,n1487);
    or g1363(n1253 ,n7[6] ,n1197);
    nand g1364(n1416 ,n2378 ,n1289);
    nand g1365(n11[36] ,n2066 ,n2078);
    xnor g1366(n2429 ,n953 ,n1114);
    nand g1367(n81 ,n2325 ,n11[33]);
    xnor g1368(n3[57] ,n2111 ,n7[57]);
    nand g1369(n252 ,n116 ,n251);
    dff g1370(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2021), .Q(n13[1]));
    or g1371(n1337 ,n8[61] ,n1188);
    nand g1372(n1788 ,n1204 ,n1496);
    nand g1373(n82 ,n2316 ,n11[40]);
    nand g1374(n1964 ,n1569 ,n1762);
    not g1375(n1137 ,n10[2]);
    nand g1376(n512 ,n341 ,n511);
    nand g1377(n1638 ,n1222 ,n1496);
    xnor g1378(n3[40] ,n2108 ,n7[40]);
    nor g1379(n1037 ,n996 ,n1036);
    xnor g1380(n2354 ,n2064 ,n2[46]);
    nand g1381(n1624 ,n1209 ,n1488);
    nand g1382(n1656 ,n1242 ,n1497);
    nand g1383(n349 ,n2186 ,n11[39]);
    nor g1384(n880 ,n2488 ,n11[42]);
    nor g1385(n767 ,n671 ,n766);
    not g1386(n482 ,n481);
    xnor g1387(n2457 ,n730 ,n773);
    nor g1388(n657 ,n2[17] ,n2[81]);
    xnor g1389(n3[61] ,n2103 ,n7[61]);
    nor g1390(n1094 ,n886 ,n1093);
    or g1391(n1338 ,n6[24] ,n1195);
    xnor g1392(n3[52] ,n2100 ,n7[52]);
    nand g1393(n338 ,n2183 ,n11[36]);
    nor g1394(n811 ,n628 ,n810);
    xnor g1395(n2141 ,n550 ,n405);
    not g1396(n434 ,n433);
    dff g1397(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1843), .Q(n7[23]));
    nand g1398(n253 ,n26 ,n252);
    nand g1399(n1798 ,n1376 ,n1495);
    nand g1400(n2022 ,n9[55] ,n1914);
    nand g1401(n622 ,n358 ,n621);
    or g1402(n1319 ,n8[17] ,n1190);
    dff g1403(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1937), .Q(n6[30]));
    or g1404(n1322 ,n6[45] ,n1188);
    nor g1405(n886 ,n2526 ,n11[45]);
    or g1406(n1316 ,n6[44] ,n1187);
    xnor g1407(n155 ,n11[37] ,n2345);
    xnor g1408(n4[43] ,n2105 ,n8[43]);
    xnor g1409(n2512 ,n2074 ,n2513);
    nor g1410(n1114 ,n907 ,n1113);
    nor g1411(n773 ,n645 ,n772);
    xnor g1412(n2484 ,n2071 ,n2485);
    nand g1413(n1676 ,n1268 ,n1496);
    or g1414(n1375 ,n7[52] ,n1196);
    xnor g1415(n2558 ,n2064 ,n2559);
    not g1416(n408 ,n407);
    or g1417(n1321 ,n6[22] ,n1197);
    nand g1418(n1673 ,n1264 ,n1498);
    xnor g1419(n2256 ,n141 ,n214);
    nand g1420(n310 ,n115 ,n309);
    nand g1421(n2021 ,n1128 ,n1915);
    nor g1422(n671 ,n2[7] ,n2[71]);
    xnor g1423(n2207 ,n2[91] ,n2076);
    nor g1424(n1014 ,n898 ,n1013);
    or g1425(n1306 ,n6[38] ,n1197);
    xnor g1426(n2393 ,n1001 ,n1042);
    nand g1427(n123 ,n2345 ,n11[37]);
    xnor g1428(n2496 ,n2072 ,n2497);
    nand g1429(n1763 ,n1344 ,n1501);
    xnor g1430(n2266 ,n150 ,n234);
    nor g1431(n1021 ,n980 ,n1020);
    nor g1432(n882 ,n2492 ,n11[44]);
    nand g1433(n1792 ,n1373 ,n1499);
    xnor g1434(n986 ,n11[39] ,n2514);
    xor g1435(n2109 ,n9[60] ,n2085);
    dff g1436(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1862), .Q(n7[6]));
    nand g1437(n1593 ,n2386 ,n1289);
    xor g1438(n2563 ,n12[1] ,n12[0]);
    nand g1439(n1572 ,n2125 ,n1289);
    nor g1440(n643 ,n2[42] ,n2[106]);
    xnor g1441(n994 ,n11[35] ,n2538);
    nand g1442(n219 ,n66 ,n218);
    nand g1443(n1712 ,n1260 ,n1493);
    xnor g1444(n2125 ,n518 ,n443);
    xnor g1445(n748 ,n2[21] ,n2[85]);
    or g1446(n1277 ,n8[49] ,n1190);
    nor g1447(n913 ,n2462 ,n11[45]);
    nor g1448(n852 ,n725 ,n851);
    nand g1449(n119 ,n2311 ,n11[35]);
    or g1450(n1215 ,n7[33] ,n1190);
    or g1451(n41 ,n2337 ,n11[45]);
    xnor g1452(n2381 ,n1018 ,n978);
    nand g1453(n1735 ,n1380 ,n1497);
    nor g1454(n1196 ,n1143 ,n1155);
    or g1455(n15 ,n2341 ,n11[33]);
    or g1456(n1273 ,n7[30] ,n1192);
    xnor g1457(n2378 ,n1012 ,n971);
    xnor g1458(n2355 ,n2072 ,n2[47]);
    nor g1459(n1013 ,n971 ,n1012);
    xnor g1460(n2119 ,n506 ,n425);
    nand g1461(n517 ,n383 ,n516);
    xor g1462(n2102 ,n9[53] ,n2094);
    xnor g1463(n753 ,n2[23] ,n2[87]);
    nor g1464(n783 ,n634 ,n782);
    dff g1465(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1830), .Q(n6[6]));
    xnor g1466(n3[35] ,n2112 ,n7[35]);
    nand g1467(n1585 ,n2388 ,n1289);
    xnor g1468(n2388 ,n1032 ,n992);
    xnor g1469(n2120 ,n508 ,n388);
    xnor g1470(n979 ,n11[37] ,n2510);
    nand g1471(n1907 ,n1516 ,n1707);
    nand g1472(n588 ,n372 ,n587);
    xnor g1473(n967 ,n2444 ,n11[36]);
    xor g1474(n2101 ,n9[58] ,n2095);
    nand g1475(n559 ,n394 ,n558);
    xnor g1476(n2143 ,n554 ,n451);
    nand g1477(n1484 ,n2167 ,n1289);
    or g1478(n1222 ,n7[26] ,n1198);
    nand g1479(n1826 ,n1411 ,n1626);
    nand g1480(n1473 ,n2149 ,n1289);
    xnor g1481(n2448 ,n2074 ,n2449);
    nor g1482(n683 ,n2[3] ,n2[67]);
    xnor g1483(n2311 ,n2078 ,n2[3]);
    nand g1484(n1746 ,n1340 ,n1487);
    xnor g1485(n5[9] ,n2111 ,n6[9]);
    nor g1486(n768 ,n741 ,n767);
    xnor g1487(n2531 ,n722 ,n847);
    or g1488(n1203 ,n7[42] ,n1198);
    xnor g1489(n2197 ,n2[81] ,n2073);
    nand g1490(n1733 ,n1323 ,n1493);
    xnor g1491(n405 ,n11[42] ,n2205);
    xnor g1492(n947 ,n11[44] ,n2492);
    nand g1493(n519 ,n444 ,n518);
    dff g1494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1846), .Q(n7[21]));
    nor g1495(n1172 ,n9[57] ,n1155);
    nor g1496(n891 ,n2502 ,n11[33]);
    xnor g1497(n2395 ,n1004 ,n1046);
    nand g1498(n80 ,n2359 ,n11[35]);
    nand g1499(n1633 ,n1273 ,n1497);
    nand g1500(n596 ,n373 ,n595);
    nor g1501(n924 ,n2444 ,n11[36]);
    nand g1502(n332 ,n2203 ,n11[40]);
    or g1503(n1311 ,n6[43] ,n1186);
    xnor g1504(n2255 ,n179 ,n212);
    xnor g1505(n709 ,n2[56] ,n2[120]);
    xnor g1506(n2209 ,n2[93] ,n2075);
    nand g1507(n573 ,n436 ,n572);
    nor g1508(n761 ,n686 ,n760);
    nand g1509(n1455 ,n2250 ,n1289);
    nand g1510(n1772 ,n1353 ,n1488);
    nand g1511(n518 ,n346 ,n517);
    nand g1512(n258 ,n131 ,n257);
    xnor g1513(n969 ,n11[35] ,n2506);
    nand g1514(n1988 ,n1590 ,n1786);
    nor g1515(n931 ,n2480 ,n11[38]);
    or g1516(n38 ,n2344 ,n11[36]);
    or g1517(n60 ,n2324 ,n11[32]);
    dff g1518(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1836), .Q(n7[29]));
    nand g1519(n1463 ,n2434 ,n1289);
    nor g1520(n863 ,n629 ,n862);
    xnor g1521(n2401 ,n947 ,n1058);
    or g1522(n1368 ,n7[56] ,n1195);
    not g1523(n957 ,n956);
    nand g1524(n521 ,n446 ,n520);
    nand g1525(n1655 ,n1241 ,n1493);
    not g1526(n484 ,n483);
    nand g1527(n1881 ,n1614 ,n1678);
    nor g1528(n680 ,n2[11] ,n2[75]);
    or g1529(n47 ,n2325 ,n11[33]);
    nor g1530(n1161 ,n9[51] ,n1155);
    nand g1531(n1886 ,n1483 ,n1686);
    nand g1532(n1834 ,n1508 ,n1633);
    nand g1533(n1537 ,n2404 ,n1289);
    nand g1534(n1718 ,n1230 ,n1496);
    nand g1535(n1821 ,n1405 ,n1620);
    nand g1536(n1127 ,n12[1] ,n12[0]);
    nand g1537(n1775 ,n1356 ,n1495);
    nor g1538(n910 ,n2466 ,n11[31]);
    nand g1539(n318 ,n2208 ,n11[45]);
    dff g1540(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1981), .Q(n8[0]));
    or g1541(n1259 ,n7[1] ,n1190);
    nor g1542(n803 ,n656 ,n802);
    xnor g1543(n2483 ,n702 ,n799);
    or g1544(n1384 ,n7[45] ,n1188);
    nand g1545(n1708 ,n1281 ,n1489);
    nand g1546(n104 ,n2358 ,n11[34]);
    nor g1547(n1048 ,n931 ,n1047);
    nor g1548(n823 ,n666 ,n822);
    xnor g1549(n2486 ,n2077 ,n2487);
    nor g1550(n826 ,n727 ,n825);
    xnor g1551(n2451 ,n741 ,n767);
    xnor g1552(n2333 ,n2071 ,n2[25]);
    nand g1553(n1659 ,n1245 ,n1501);
    not g1554(n2071 ,n9[57]);
    nand g1555(n554 ,n326 ,n553);
    xnor g1556(n172 ,n11[38] ,n2362);
    nand g1557(n1931 ,n1536 ,n1729);
    nand g1558(n1758 ,n1315 ,n1497);
    nand g1559(n121 ,n2309 ,n11[33]);
    xnor g1560(n2438 ,n2439 ,n2068);
    nor g1561(n915 ,n2512 ,n11[38]);
    nand g1562(n94 ,n2312 ,n11[36]);
    xnor g1563(n2315 ,n2074 ,n2[7]);
    xnor g1564(n386 ,n11[38] ,n2217);
    nand g1565(n1816 ,n1518 ,n1711);
    xnor g1566(n3[53] ,n2102 ,n7[53]);
    nand g1567(n1778 ,n1357 ,n1491);
    nor g1568(n1192 ,n1139 ,n1155);
    xnor g1569(n4[33] ,n2114 ,n8[33]);
    nand g1570(n2050 ,n2016 ,n2034);
    xnor g1571(n2422 ,n962 ,n1100);
    xnor g1572(n740 ,n2[17] ,n2[81]);
    xnor g1573(n2178 ,n624 ,n483);
    xnor g1574(n2211 ,n2[95] ,n2072);
    nand g1575(n103 ,n2342 ,n11[34]);
    nand g1576(n281 ,n50 ,n280);
    xnor g1577(n2231 ,n2[115] ,n2078);
    nand g1578(n2026 ,n9[51] ,n1914);
    nor g1579(n627 ,n2[47] ,n2[111]);
    xnor g1580(n5[59] ,n2105 ,n6[59]);
    dff g1581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1865), .Q(n7[5]));
    nand g1582(n289 ,n23 ,n288);
    nand g1583(n1840 ,n1425 ,n1634);
    xnor g1584(n2158 ,n584 ,n475);
    nand g1585(n1851 ,n1439 ,n1652);
    dff g1586(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[10]), .Q(n9[58]));
    or g1587(n1202 ,n6[13] ,n1188);
    xnor g1588(n453 ,n11[45] ,n2192);
    dff g1589(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1910), .Q(n6[38]));
    nor g1590(n1292 ,n1155 ,n1184);
    nand g1591(n2030 ,n9[56] ,n1914);
    nand g1592(n1916 ,n1435 ,n1648);
    nor g1593(n1059 ,n947 ,n1058);
    nor g1594(n1022 ,n904 ,n1021);
    nand g1595(n1526 ,n2408 ,n1289);
    nand g1596(n215 ,n54 ,n214);
    dff g1597(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1828), .Q(n7[35]));
    dff g1598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1939), .Q(n8[28]));
    nand g1599(n257 ,n15 ,n256);
    xnor g1600(n157 ,n11[38] ,n2346);
    or g1601(n1298 ,n8[56] ,n1195);
    dff g1602(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1909), .Q(n8[49]));
    nand g1603(n1467 ,n2431 ,n1289);
    nand g1604(n353 ,n2218 ,n11[39]);
    or g1605(n1224 ,n7[22] ,n1197);
    nor g1606(n630 ,n2[23] ,n2[87]);
    dff g1607(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[9]), .Q(n9[57]));
    nand g1608(n1927 ,n1533 ,n1727);
    nand g1609(n1879 ,n1469 ,n1685);
    xnor g1610(n2519 ,n747 ,n835);
    nand g1611(n1448 ,n2254 ,n1289);
    nand g1612(n254 ,n117 ,n253);
    nand g1613(n1472 ,n12[0] ,n1295);
    xnor g1614(n2276 ,n136 ,n254);
    nand g1615(n1773 ,n1354 ,n1492);
    nand g1616(n11[41] ,n2077 ,n2070);
    xnor g1617(n483 ,n2242 ,n9[62]);
    xnor g1618(n2368 ,n2[60] ,n2079);
    nand g1619(n566 ,n347 ,n565);
    xnor g1620(n3[9] ,n2111 ,n7[9]);
    nand g1621(n1757 ,n1314 ,n1493);
    nor g1622(n1199 ,n1140 ,n1155);
    xnor g1623(n2212 ,n2[96] ,n2067);
    xnor g1624(n2471 ,n743 ,n787);
    xnor g1625(n5[45] ,n2103 ,n6[45]);
    not g1626(n1142 ,n10[15]);
    nor g1627(n854 ,n733 ,n853);
    nand g1628(n1679 ,n1392 ,n1494);
    nor g1629(n1095 ,n954 ,n1094);
    xnor g1630(n2533 ,n714 ,n849);
    not g1631(n1145 ,n13[2]);
    nand g1632(n579 ,n456 ,n578);
    nor g1633(n885 ,n2548 ,n11[40]);
    or g1634(n1201 ,n1183 ,n1174);
    xnor g1635(n718 ,n2[34] ,n2[98]);
    xor g1636(n2116 ,n11[33] ,n2180);
    xnor g1637(n2216 ,n2[100] ,n2065);
    nand g1638(n551 ,n406 ,n550);
    nand g1639(n342 ,n2216 ,n11[37]);
    dff g1640(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1834), .Q(n7[30]));
    xnor g1641(n2420 ,n949 ,n1096);
    nand g1642(n689 ,n2[0] ,n2[64]);
    nand g1643(n1405 ,n2284 ,n1289);
    or g1644(n1654 ,n1292 ,n1400);
    xnor g1645(n5[35] ,n2112 ,n6[35]);
    nand g1646(n1974 ,n1578 ,n1770);
    xnor g1647(n2474 ,n2065 ,n2475);
    nor g1648(n69 ,n2309 ,n11[33]);
    nand g1649(n1870 ,n1461 ,n1670);
    nand g1650(n1584 ,n2143 ,n1289);
    nand g1651(n565 ,n408 ,n564);
    dff g1652(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1944), .Q(n8[25]));
    nand g1653(n1590 ,n2304 ,n1289);
    xnor g1654(n3[37] ,n2102 ,n7[37]);
    nor g1655(n1084 ,n916 ,n1083);
    or g1656(n1233 ,n8[60] ,n1187);
    nor g1657(n1069 ,n961 ,n1068);
    dff g1658(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2053), .Q(n10[10]));
    nand g1659(n603 ,n410 ,n602);
    xnor g1660(n2195 ,n2[79] ,n2072);
    xnor g1661(n2343 ,n2078 ,n2[35]);
    xnor g1662(n723 ,n2[7] ,n2[71]);
    nor g1663(n1093 ,n965 ,n1092);
    xnor g1664(n152 ,n11[35] ,n2343);
    nand g1665(n1695 ,n1310 ,n1496);
    xnor g1666(n4[29] ,n2103 ,n8[29]);
    xnor g1667(n2138 ,n544 ,n497);
    xnor g1668(n5[41] ,n2111 ,n6[41]);
    xnor g1669(n2441 ,n715 ,n757);
    nor g1670(n791 ,n663 ,n790);
    nor g1671(n927 ,n2478 ,n11[37]);
    nand g1672(n1961 ,n1564 ,n1758);
    xnor g1673(n2478 ,n2069 ,n2479);
    nand g1674(n1766 ,n1348 ,n1486);
    nor g1675(n1086 ,n920 ,n1085);
    xnor g1676(n5[44] ,n2109 ,n6[44]);
    xnor g1677(n2288 ,n138 ,n278);
    nand g1678(n567 ,n420 ,n566);
    not g1679(n442 ,n441);
    dff g1680(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1876), .Q(n6[58]));
    xnor g1681(n3[48] ,n2107 ,n7[48]);
    nand g1682(n1737 ,n1379 ,n1498);
    xnor g1683(n2322 ,n2064 ,n2[14]);
    nand g1684(n1874 ,n1466 ,n1674);
    or g1685(n1256 ,n7[3] ,n1199);
    or g1686(n1255 ,n7[4] ,n1196);
    nor g1687(n777 ,n647 ,n776);
    dff g1688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1975), .Q(n8[5]));
    nand g1689(n1459 ,n2246 ,n1289);
    xnor g1690(n2524 ,n2075 ,n2525);
    nor g1691(n635 ,n2[33] ,n2[97]);
    xor g1692(n2106 ,n9[55] ,n2090);
    nor g1693(n1121 ,n944 ,n1120);
    xnor g1694(n2370 ,n2[62] ,n2064);
    nand g1695(n277 ,n53 ,n276);
    nor g1696(n860 ,n701 ,n859);
    xnor g1697(n703 ,n2[25] ,n2[89]);
    xnor g1698(n2452 ,n2071 ,n2453);
    xnor g1699(n751 ,n2[43] ,n2[107]);
    nand g1700(n1803 ,n1381 ,n1496);
    xnor g1701(n2384 ,n1024 ,n984);
    xnor g1702(n5[60] ,n2109 ,n6[60]);
    or g1703(n1236 ,n7[19] ,n1199);
    dff g1704(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1918), .Q(n8[42]));
    dff g1705(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1873), .Q(n6[61]));
    not g1706(n470 ,n469);
    nor g1707(n934 ,n2486 ,n11[41]);
    xnor g1708(n2357 ,n2073 ,n2[49]);
    nor g1709(n916 ,n2516 ,n11[40]);
    nor g1710(n1123 ,n968 ,n1122);
    nand g1711(n323 ,n2239 ,n11[44]);
    xnor g1712(n382 ,n11[41] ,n2188);
    not g1713(n2079 ,n9[60]);
    nand g1714(n1434 ,n2263 ,n1289);
    nand g1715(n557 ,n398 ,n556);
    xnor g1716(n5[13] ,n2103 ,n6[13]);
    nand g1717(n1888 ,n1550 ,n1688);
    nand g1718(n560 ,n324 ,n559);
    xnor g1719(n2191 ,n2[75] ,n2076);
    nor g1720(n1099 ,n943 ,n1098);
    nand g1721(n376 ,n2201 ,n11[38]);
    not g1722(n468 ,n467);
    nor g1723(n1078 ,n883 ,n1077);
    nand g1724(n124 ,n2364 ,n11[40]);
    dff g1725(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1893), .Q(n8[60]));
    nand g1726(n326 ,n2206 ,n11[43]);
    dff g1727(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1863), .Q(n7[7]));
    nand g1728(n1183 ,n1149 ,n1153);
    nand g1729(n250 ,n114 ,n249);
    xnor g1730(n2297 ,n169 ,n296);
    xnor g1731(n2201 ,n2[85] ,n2066);
    or g1732(n1248 ,n7[10] ,n1198);
    not g1733(n460 ,n459);
    xnor g1734(n2535 ,n725 ,n851);
    xnor g1735(n5[43] ,n2105 ,n6[43]);
    nand g1736(n1903 ,n1511 ,n1702);
    xnor g1737(n5[62] ,n2113 ,n6[62]);
    xnor g1738(n2449 ,n723 ,n765);
    nand g1739(n1574 ,n2391 ,n1289);
    dff g1740(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2054), .Q(n10[9]));
    nand g1741(n1618 ,n1203 ,n1496);
    xnor g1742(n491 ,n11[38] ,n2201);
    xnor g1743(n2219 ,n2[103] ,n2074);
    nand g1744(n1600 ,n2298 ,n1289);
    nor g1745(n769 ,n641 ,n768);
    xnor g1746(n2291 ,n143 ,n284);
    nand g1747(n1721 ,n1226 ,n1495);
    nand g1748(n1764 ,n1471 ,n1481);
    xnor g1749(n142 ,n11[46] ,n2354);
    xnor g1750(n2500 ,n2073 ,n2501);
    xnor g1751(n962 ,n11[33] ,n2534);
    xnor g1752(n2491 ,n693 ,n807);
    nor g1753(n1061 ,n945 ,n1060);
    nand g1754(n2097 ,n10[3] ,n11[35]);
    dff g1755(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2059), .Q(n10[0]));
    xnor g1756(n2127 ,n522 ,n449);
    nor g1757(n763 ,n638 ,n762);
    not g1758(n389 ,n388);
    or g1759(n1296 ,n6[9] ,n1185);
    xnor g1760(n2458 ,n2459 ,n2079);
    nand g1761(n344 ,n2242 ,n9[62]);
    not g1762(n424 ,n423);
    nor g1763(n652 ,n2[51] ,n2[115]);
    dff g1764(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1899), .Q(n8[55]));
    nand g1765(n1980 ,n1442 ,n1779);
    xnor g1766(n2270 ,n191 ,n242);
    xnor g1767(n2431 ,n1002 ,n1118);
    nand g1768(n328 ,n2207 ,n11[44]);
    dff g1769(.RN(1'b1), .SN(n2567), .CK(n0), .D(n9[48]), .Q(n14[2]));
    xnor g1770(n4[4] ,n2100 ,n8[4]);
    nand g1771(n532 ,n363 ,n531);
    xnor g1772(n2140 ,n548 ,n411);
    xnor g1773(n713 ,n2[33] ,n2[97]);
    nor g1774(n1087 ,n998 ,n1086);
    nand g1775(n1999 ,n1603 ,n1796);
    nand g1776(n1579 ,n2121 ,n1289);
    not g1777(n474 ,n473);
    nor g1778(n1159 ,n9[50] ,n1155);
    nand g1779(n234 ,n91 ,n233);
    or g1780(n1206 ,n7[40] ,n1195);
    nand g1781(n1820 ,n1404 ,n1619);
    or g1782(n1383 ,n7[46] ,n1192);
    xnor g1783(n2404 ,n952 ,n1064);
    nand g1784(n1892 ,n1505 ,n1696);
    or g1785(n1210 ,n6[7] ,n1189);
    xnor g1786(n4[37] ,n2102 ,n8[37]);
    nand g1787(n1761 ,n1342 ,n1488);
    xor g1788(n2115 ,n2089 ,n9[47]);
    nand g1789(n1933 ,n1473 ,n1730);
    xnor g1790(n158 ,n11[39] ,n2347);
    nand g1791(n1729 ,n1270 ,n1491);
    not g1792(n432 ,n431);
    nand g1793(n205 ,n20 ,n204);
    dff g1794(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1904), .Q(n8[52]));
    or g1795(n68 ,n2362 ,n11[38]);
    nor g1796(n1058 ,n884 ,n1057);
    nand g1797(n1952 ,n1557 ,n1752);
    nand g1798(n1571 ,n2126 ,n1289);
    nand g1799(n1970 ,n1572 ,n1766);
    xnor g1800(n2196 ,n2[80] ,n2067);
    xnor g1801(n5[0] ,n2098 ,n6[0]);
    nor g1802(n821 ,n637 ,n820);
    nand g1803(n92 ,n2351 ,n11[43]);
    nor g1804(n807 ,n679 ,n806);
    or g1805(n46 ,n2332 ,n11[40]);
    not g1806(n448 ,n447);
    nor g1807(n827 ,n646 ,n826);
    nor g1808(n1053 ,n951 ,n1052);
    nor g1809(n873 ,n681 ,n872);
    xnor g1810(n707 ,n2[1] ,n2[65]);
    nand g1811(n1976 ,n1581 ,n1774);
    nand g1812(n1765 ,n1346 ,n1496);
    dff g1813(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1923), .Q(n6[35]));
    nand g1814(n592 ,n317 ,n591);
    or g1815(n64 ,n2335 ,n11[43]);
    nand g1816(n1662 ,n1250 ,n1489);
    or g1817(n1370 ,n6[30] ,n1192);
    nand g1818(n1632 ,n1287 ,n1488);
    nand g1819(n11[37] ,n2069 ,n2065);
    not g1820(n476 ,n475);
    dff g1821(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1819), .Q(n7[42]));
    xnor g1822(n744 ,n2[53] ,n2[117]);
    dff g1823(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1818), .Q(n6[9]));
    nand g1824(n303 ,n62 ,n302);
    nand g1825(n1962 ,n1523 ,n1809);
    nor g1826(n1085 ,n995 ,n1084);
    xnor g1827(n2561 ,n690 ,n877);
    or g1828(n1231 ,n6[2] ,n1193);
    nand g1829(n2083 ,n10[9] ,n11[41]);
    xnor g1830(n3[11] ,n2105 ,n7[11]);
    nand g1831(n295 ,n21 ,n294);
    nand g1832(n365 ,n2196 ,n11[33]);
    or g1833(n58 ,n2316 ,n11[40]);
    xnor g1834(n380 ,n11[35] ,n2230);
    nor g1835(n851 ,n640 ,n850);
    xnor g1836(n2206 ,n2[90] ,n2077);
    nand g1837(n1674 ,n1266 ,n1499);
    dff g1838(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1949), .Q(n8[22]));
    or g1839(n1205 ,n8[37] ,n1191);
    dff g1840(.RN(n2567), .SN(1'b1), .CK(n0), .D(n9[53]), .Q(n9[54]));
    dff g1841(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[11]), .Q(n9[59]));
    nand g1842(n297 ,n73 ,n296);
    not g1843(n456 ,n455);
    xnor g1844(n2299 ,n173 ,n300);
    xnor g1845(n421 ,n11[34] ,n2181);
    nand g1846(n1649 ,n1236 ,n1495);
    nor g1847(n839 ,n675 ,n838);
    nor g1848(n1027 ,n985 ,n1026);
    xnor g1849(n5[54] ,n2104 ,n6[54]);
    or g1850(n1242 ,n7[14] ,n1192);
    xnor g1851(n3[18] ,n2110 ,n7[18]);
    nand g1852(n1509 ,n2127 ,n1289);
    nand g1853(n1875 ,n1467 ,n1675);
    xnor g1854(n2129 ,n526 ,n457);
    not g1855(n708 ,n707);
    xnor g1856(n5[52] ,n2100 ,n6[52]);
    xnor g1857(n2222 ,n2[106] ,n2077);
    nand g1858(n540 ,n371 ,n539);
    dff g1859(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1810), .Q(n12[0]));
    or g1860(n1399 ,n7[48] ,n1292);
    dff g1861(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2007), .Q(n7[45]));
    not g1862(n416 ,n415);
    xnor g1863(n2306 ,n2370 ,n314);
    not g1864(n2067 ,n9[48]);
    xnor g1865(n5[39] ,n2106 ,n6[39]);
    nand g1866(n1511 ,n2169 ,n1289);
    dff g1867(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1940), .Q(n8[27]));
    or g1868(n1397 ,n6[16] ,n1292);
    not g1869(n466 ,n465);
    or g1870(n1268 ,n6[58] ,n1198);
    nand g1871(n1979 ,n1583 ,n1778);
    xnor g1872(n497 ,n11[39] ,n2202);
    nand g1873(n556 ,n328 ,n555);
    nand g1874(n370 ,n2233 ,n11[38]);
    nand g1875(n325 ,n2241 ,n11[46]);
    nand g1876(n584 ,n366 ,n583);
    xnor g1877(n2247 ,n180 ,n196);
    xnor g1878(n3[29] ,n2103 ,n7[29]);
    xor g1879(n2117 ,n421 ,n348);
    nand g1880(n2003 ,n1606 ,n1800);
    nand g1881(n2047 ,n10[5] ,n2031);
    xnor g1882(n2365 ,n2071 ,n2[57]);
    xnor g1883(n2492 ,n2075 ,n2493);
    not g1884(n2078 ,n9[51]);
    nand g1885(n599 ,n414 ,n598);
    xnor g1886(n700 ,n2[44] ,n2[108]);
    xnor g1887(n2386 ,n1028 ,n988);
    not g1888(n420 ,n419);
    nand g1889(n2094 ,n10[5] ,n11[37]);
    nand g1890(n1780 ,n1398 ,n1494);
    nand g1891(n2017 ,n9[60] ,n1914);
    xnor g1892(n2453 ,n726 ,n769);
    nor g1893(n1293 ,n1 ,n1176);
    nand g1894(n2000 ,n1604 ,n1798);
    nand g1895(n1983 ,n1587 ,n1782);
    dff g1896(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1817), .Q(n7[43]));
    nand g1897(n317 ,n2225 ,n11[46]);
    dff g1898(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1930), .Q(n6[33]));
    xnor g1899(n5[51] ,n2112 ,n6[51]);
    nand g1900(n2055 ,n2017 ,n2035);
    xnor g1901(n943 ,n11[32] ,n2532);
    not g1902(n462 ,n461);
    nor g1903(n1026 ,n909 ,n1025);
    or g1904(n1382 ,n7[29] ,n1188);
    nand g1905(n1538 ,n2403 ,n1289);
    xnor g1906(n2485 ,n703 ,n801);
    or g1907(n1204 ,n7[58] ,n1198);
    xnor g1908(n2416 ,n1003 ,n1088);
    nand g1909(n1977 ,n1456 ,n1775);
    nand g1910(n235 ,n59 ,n234);
    nand g1911(n1902 ,n1521 ,n1701);
    dff g1912(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1993), .Q(n7[55]));
    xnor g1913(n3[44] ,n2109 ,n7[44]);
    nor g1914(n795 ,n670 ,n794);
    nand g1915(n1923 ,n1527 ,n1721);
    nor g1916(n758 ,n715 ,n757);
    xnor g1917(n2390 ,n1036 ,n996);
    nor g1918(n1125 ,n946 ,n1124);
    xnor g1919(n2548 ,n2071 ,n2549);
    dff g1920(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[5]), .Q(n9[53]));
    nand g1921(n1450 ,n2252 ,n1289);
    or g1922(n52 ,n2352 ,n11[44]);
    or g1923(n1339 ,n6[23] ,n1189);
    xnor g1924(n2260 ,n137 ,n222);
    nand g1925(n225 ,n47 ,n224);
    nand g1926(n1446 ,n2372 ,n1289);
    nand g1927(n1779 ,n1239 ,n1492);
    xnor g1928(n160 ,n11[41] ,n2349);
    nand g1929(n314 ,n2369 ,n313);
    nand g1930(n1441 ,n2259 ,n1289);
    nor g1931(n878 ,n2468 ,n11[32]);
    nand g1932(n1920 ,n1526 ,n1717);
    not g1933(n446 ,n445);
    xnor g1934(n395 ,n11[31] ,n2210);
    nand g1935(n1901 ,n1510 ,n1703);
    dff g1936(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1823), .Q(n7[38]));
    nand g1937(n514 ,n349 ,n513);
    xnor g1938(n2508 ,n2066 ,n2509);
    nand g1939(n1503 ,n2418 ,n1289);
    nor g1940(n802 ,n703 ,n801);
    nor g1941(n923 ,n2520 ,n11[42]);
    nand g1942(n1713 ,n1261 ,n1497);
    nand g1943(n1860 ,n1449 ,n1661);
    nand g1944(n89 ,n2313 ,n11[37]);
    nand g1945(n618 ,n375 ,n617);
    xnor g1946(n2556 ,n2557 ,n2075);
    nand g1947(n1641 ,n1228 ,n1489);
    or g1948(n1221 ,n7[27] ,n1186);
    nand g1949(n528 ,n357 ,n527);
    nand g1950(n1951 ,n1555 ,n1750);
    not g1951(n1133 ,n10[10]);
    or g1952(n24 ,n2338 ,n11[46]);
    xnor g1953(n2511 ,n732 ,n827);
    nand g1954(n610 ,n321 ,n609);
    nand g1955(n1728 ,n1251 ,n1495);
    nor g1956(n760 ,n717 ,n759);
    xnor g1957(n2362 ,n2069 ,n2[54]);
    nand g1958(n1936 ,n1599 ,n1735);
    not g1959(n383 ,n382);
    nand g1960(n1630 ,n1389 ,n1494);
    or g1961(n1365 ,n7[49] ,n1190);
    nand g1962(n1968 ,n1571 ,n1765);
    xnor g1963(n750 ,n2[22] ,n2[86]);
    or g1964(n1227 ,n6[36] ,n1196);
    nor g1965(n1116 ,n885 ,n1115);
    nand g1966(n1623 ,n1313 ,n1487);
    xnor g1967(n2383 ,n981 ,n1022);
    xor g1968(n2118 ,n392 ,n504);
    nand g1969(n1652 ,n1238 ,n1492);
    xnor g1970(n2371 ,n2[63] ,n2072);
    dff g1971(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1897), .Q(n8[57]));
    or g1972(n1502 ,n12[0] ,n1294);
    nand g1973(n307 ,n42 ,n306);
    nor g1974(n814 ,n699 ,n813);
    nand g1975(n2001 ,n1605 ,n1799);
    nand g1976(n240 ,n98 ,n239);
    not g1977(n391 ,n390);
    xnor g1978(n705 ,n2[35] ,n2[99]);
    nand g1979(n1717 ,n1227 ,n1490);
    nand g1980(n583 ,n468 ,n582);
    nor g1981(n1106 ,n906 ,n1105);
    xnor g1982(n3[46] ,n2113 ,n7[46]);
    nand g1983(n2005 ,n1611 ,n1802);
    xnor g1984(n2341 ,n2073 ,n2[33]);
    nand g1985(n1809 ,n1308 ,n1499);
    xnor g1986(n180 ,n11[35] ,n2311);
    nand g1987(n1475 ,n12[2] ,n1295);
    nor g1988(n1074 ,n897 ,n1073);
    nand g1989(n11[32] ,n2072 ,n2073);
    xnor g1990(n2522 ,n2079 ,n2523);
    nand g1991(n1966 ,n1570 ,n1761);
    nor g1992(n1651 ,n9[48] ,n1446);
    xnor g1993(n959 ,n11[42] ,n2488);
    nand g1994(n1981 ,n1586 ,n1780);
    nand g1995(n582 ,n360 ,n581);
    or g1996(n1394 ,n6[48] ,n1292);
    xnor g1997(n2287 ,n162 ,n276);
    nand g1998(n1895 ,n1506 ,n1695);
    nand g1999(n1518 ,n2411 ,n1289);
    nand g2000(n586 ,n369 ,n585);
    nand g2001(n246 ,n107 ,n245);
    dff g2002(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1871), .Q(n6[63]));
    nor g2003(n1036 ,n878 ,n1035);
    xnor g2004(n4[30] ,n2113 ,n8[30]);
    nor g2005(n645 ,n2[10] ,n2[74]);
    xnor g2006(n2326 ,n2068 ,n2[18]);
    dff g2007(.RN(n2567), .SN(1'b1), .CK(n0), .D(n9[48]), .Q(n9[49]));
    nand g2008(n1715 ,n1387 ,n1501);
    nand g2009(n516 ,n345 ,n515);
    nand g2010(n2049 ,n2015 ,n2033);
    xnor g2011(n2318 ,n2077 ,n2[10]);
    nor g2012(n866 ,n721 ,n865);
    nor g2013(n856 ,n739 ,n855);
    xnor g2014(n4[28] ,n2109 ,n8[28]);
    nand g2015(n86 ,n2350 ,n11[42]);
    nand g2016(n1474 ,n2562 ,n1293);
    nor g2017(n855 ,n652 ,n854);
    nor g2018(n818 ,n713 ,n817);
    xnor g2019(n5[32] ,n2107 ,n6[32]);
    nand g2020(n1731 ,n1395 ,n1494);
    nor g2021(n677 ,n2[14] ,n2[78]);
    dff g2022(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1835), .Q(n6[5]));
    or g2023(n1274 ,n6[49] ,n1190);
    xnor g2024(n2167 ,n602 ,n409);
    xnor g2025(n725 ,n2[50] ,n2[114]);
    nand g2026(n1829 ,n1414 ,n1628);
    dff g2027(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1983), .Q(n7[63]));
    xnor g2028(n2501 ,n713 ,n817);
    not g2029(n385 ,n384);
    nand g2030(n228 ,n84 ,n227);
    nand g2031(n537 ,n480 ,n536);
    xnor g2032(n2308 ,n2[0] ,n2067);
    nand g2033(n197 ,n65 ,n196);
    nand g2034(n1530 ,n2154 ,n1289);
    xnor g2035(n2280 ,n153 ,n262);
    xnor g2036(n2521 ,n751 ,n837);
    nor g2037(n779 ,n650 ,n778);
    nor g2038(n766 ,n723 ,n765);
    nand g2039(n1534 ,n2405 ,n1289);
    xnor g2040(n4[2] ,n2110 ,n8[2]);
    dff g2041(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1856), .Q(n7[12]));
    xnor g2042(n159 ,n11[40] ,n2348);
    xnor g2043(n411 ,n11[41] ,n2204);
    nand g2044(n1622 ,n1210 ,n1500);
    xnor g2045(n3[36] ,n2100 ,n7[36]);
    nand g2046(n1542 ,n2402 ,n1289);
    nand g2047(n115 ,n2367 ,n11[43]);
    nand g2048(n1997 ,n1601 ,n1795);
    dff g2049(.RN(1'b1), .SN(n2567), .CK(n0), .D(n9[60]), .Q(n14[14]));
    xnor g2050(n2303 ,n175 ,n308);
    or g2051(n42 ,n2366 ,n11[42]);
    nor g2052(n648 ,n2[54] ,n2[118]);
    nand g2053(n757 ,n688 ,n756);
    nor g2054(n665 ,n2[28] ,n2[92]);
    nand g2055(n569 ,n424 ,n568);
    nand g2056(n1637 ,n1221 ,n1501);
    nand g2057(n1805 ,n1384 ,n1498);
    nor g2058(n838 ,n751 ,n837);
    not g2059(n418 ,n417);
    nor g2060(n1110 ,n930 ,n1109);
    nand g2061(n260 ,n103 ,n259);
    xnor g2062(n5[15] ,n2115 ,n6[15]);
    nand g2063(n1531 ,n2406 ,n1289);
    nand g2064(n1403 ,n2286 ,n1289);
    nand g2065(n1660 ,n1248 ,n1496);
    nand g2066(n126 ,n2344 ,n11[36]);
    nand g2067(n1525 ,n2158 ,n1289);
    nand g2068(n1605 ,n2294 ,n1289);
    nand g2069(n1421 ,n2157 ,n1289);
    xnor g2070(n3[45] ,n2103 ,n7[45]);
    nand g2071(n553 ,n478 ,n552);
    xnor g2072(n184 ,n11[33] ,n2325);
    dff g2073(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1848), .Q(n7[20]));
    nand g2074(n1422 ,n2273 ,n1289);
    dff g2075(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1977), .Q(n8[3]));
    not g2076(n498 ,n497);
    nand g2077(n1598 ,n2299 ,n1289);
    xnor g2078(n5[48] ,n2107 ,n6[48]);
    xnor g2079(n4[25] ,n2111 ,n8[25]);
    nand g2080(n272 ,n78 ,n271);
    nand g2081(n2035 ,n10[12] ,n2031);
    nor g2082(n850 ,n714 ,n849);
    nand g2083(n1942 ,n1549 ,n1740);
    xor g2084(n2372 ,n2[0] ,n2[64]);
    xnor g2085(n2434 ,n946 ,n1124);
    xnor g2086(n5[53] ,n2102 ,n6[53]);
    nand g2087(n11[31] ,n2064 ,n2067);
    nand g2088(n291 ,n28 ,n290);
    nand g2089(n1791 ,n1202 ,n1498);
    nand g2090(n294 ,n80 ,n293);
    or g2091(n32 ,n2346 ,n11[38]);
    nand g2092(n1559 ,n2288 ,n1289);
    xnor g2093(n2281 ,n155 ,n264);
    nand g2094(n1885 ,n1591 ,n1683);
    or g2095(n73 ,n2361 ,n11[37]);
    nor g2096(n1103 ,n970 ,n1102);
    not g2097(n398 ,n397);
    nor g2098(n1153 ,n10[10] ,n10[11]);
    xor g2099(n2437 ,n707 ,n689);
    nand g2100(n1946 ,n1562 ,n1745);
    nand g2101(n1734 ,n1271 ,n1493);
    nand g2102(n570 ,n330 ,n569);
    nand g2103(n327 ,n2210 ,n11[31]);
    nand g2104(n1954 ,n1556 ,n1749);
    xnor g2105(n4[45] ,n2103 ,n8[45]);
    nand g2106(n1714 ,n1247 ,n1498);
    xnor g2107(n3[23] ,n2106 ,n7[23]);
    nand g2108(n201 ,n35 ,n200);
    nor g2109(n1042 ,n908 ,n1041);
    nand g2110(n1789 ,n1366 ,n1486);
    nor g2111(n1088 ,n923 ,n1087);
    nand g2112(n90 ,n2314 ,n11[38]);
    nor g2113(n1111 ,n960 ,n1110);
    xnor g2114(n419 ,n11[34] ,n2213);
    nand g2115(n1184 ,n10[0] ,n1157);
    xnor g2116(n493 ,n11[31] ,n2226);
    xnor g2117(n710 ,n2[60] ,n2[124]);
    nor g2118(n841 ,n669 ,n840);
    nand g2119(n98 ,n2332 ,n11[40]);
    xnor g2120(n467 ,n11[42] ,n2221);
    nand g2121(n1477 ,n2424 ,n1289);
    nand g2122(n204 ,n90 ,n203);
    xnor g2123(n2442 ,n2443 ,n2065);
    nand g2124(n1971 ,n1573 ,n1813);
    nand g2125(n1934 ,n1540 ,n1731);
    xnor g2126(n2139 ,n546 ,n429);
    nand g2127(n347 ,n2212 ,n11[33]);
    nor g2128(n898 ,n2446 ,n11[37]);
    not g2129(n1129 ,n1);
    nor g2130(n897 ,n2506 ,n11[35]);
    xnor g2131(n968 ,n11[44] ,n2556);
    dff g2132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1954), .Q(n6[25]));
    xnor g2133(n2455 ,n728 ,n771);
    or g2134(n1318 ,n6[54] ,n1197);
    xnor g2135(n185 ,n11[37] ,n2313);
    xnor g2136(n2336 ,n2079 ,n2[28]);
    nand g2137(n267 ,n32 ,n266);
    nand g2138(n1428 ,n2375 ,n1289);
    or g2139(n67 ,n2333 ,n11[41]);
    xnor g2140(n151 ,n11[34] ,n2342);
    nand g2141(n351 ,n2237 ,n11[42]);
    nor g2142(n864 ,n709 ,n863);
    nand g2143(n111 ,n2340 ,n11[32]);
    or g2144(n1359 ,n6[15] ,n1194);
    or g2145(n1324 ,n6[8] ,n1195);
    xnor g2146(n2160 ,n588 ,n495);
    nor g2147(n629 ,n2[55] ,n2[119]);
    nor g2148(n793 ,n667 ,n792);
    nand g2149(n1412 ,n2279 ,n1289);
    dff g2150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1868), .Q(n7[2]));
    xor g2151(n2107 ,n2088 ,n9[48]);
    xnor g2152(n4[59] ,n2105 ,n8[59]);
    xnor g2153(n3[51] ,n2112 ,n7[51]);
    nor g2154(n892 ,n2500 ,n11[32]);
    nor g2155(n933 ,n2452 ,n11[40]);
    xnor g2156(n940 ,n2560 ,n11[46]);
    xnor g2157(n4[11] ,n2105 ,n8[11]);
    xnor g2158(n170 ,n11[40] ,n2316);
    xnor g2159(n5[42] ,n2101 ,n6[42]);
    nand g2160(n507 ,n426 ,n506);
    nand g2161(n1727 ,n1282 ,n1490);
    nand g2162(n1550 ,n2179 ,n1289);
    nand g2163(n1461 ,n2244 ,n1289);
    nand g2164(n1880 ,n1470 ,n1682);
    dff g2165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1820), .Q(n7[41]));
    nor g2166(n895 ,n2504 ,n11[34]);
    nand g2167(n2048 ,n2014 ,n2032);
    nand g2168(n1794 ,n1372 ,n1487);
    or g2169(n61 ,n2365 ,n11[41]);
    nand g2170(n1704 ,n1283 ,n1486);
    nor g2171(n789 ,n661 ,n788);
    nand g2172(n1436 ,n2262 ,n1289);
    nand g2173(n2054 ,n2020 ,n2038);
    nand g2174(n1597 ,n2385 ,n1289);
    xnor g2175(n2361 ,n2066 ,n2[53]);
    nand g2176(n261 ,n55 ,n260);
    xnor g2177(n2319 ,n2076 ,n2[11]);
    nand g2178(n1560 ,n2133 ,n1289);
    xnor g2179(n153 ,n11[36] ,n2344);
    xnor g2180(n2152 ,n572 ,n435);
    nand g2181(n1588 ,n2306 ,n1289);
    dff g2182(.RN(n2567), .SN(1'b1), .CK(n0), .D(n9[60]), .Q(n9[61]));
    xnor g2183(n995 ,n11[41] ,n2518);
    nand g2184(n1589 ,n2305 ,n1289);
    xnor g2185(n950 ,n11[43] ,n2490);
    xnor g2186(n2166 ,n600 ,n380);
    nand g2187(n238 ,n96 ,n237);
    not g2188(n396 ,n395);
    nand g2189(n1861 ,n1450 ,n1662);
    nor g2190(n1170 ,n9[59] ,n1155);
    nand g2191(n1720 ,n1312 ,n1489);
    nand g2192(n1719 ,n1218 ,n1486);
    nor g2193(n899 ,n2530 ,n11[31]);
    nand g2194(n1786 ,n1362 ,n1499);
    nand g2195(n1558 ,n2134 ,n1289);
    dff g2196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1842), .Q(n7[24]));
    xnor g2197(n4[21] ,n2102 ,n8[21]);
    nand g2198(n1700 ,n1299 ,n1500);
    dff g2199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1894), .Q(n8[59]));
    nand g2200(n1949 ,n1580 ,n1746);
    not g2201(n1131 ,n10[5]);
    xnor g2202(n2427 ,n960 ,n1110);
    nand g2203(n1782 ,n1358 ,n1493);
    nor g2204(n1913 ,n1178 ,n1814);
    nor g2205(n1490 ,n1162 ,n1291);
    nand g2206(n1978 ,n1582 ,n1773);
    nand g2207(n1561 ,n2395 ,n1289);
    nand g2208(n1943 ,n1547 ,n1741);
    xnor g2209(n717 ,n2[4] ,n2[68]);
    nand g2210(n1918 ,n1525 ,n1718);
    nor g2211(n764 ,n752 ,n763);
    nand g2212(n616 ,n351 ,n615);
    or g2213(n1240 ,n6[37] ,n1191);
    nor g2214(n1044 ,n922 ,n1043);
    nor g2215(n815 ,n684 ,n814);
    nand g2216(n333 ,n2205 ,n11[42]);
    nor g2217(n801 ,n655 ,n800);
    xnor g2218(n4[47] ,n2115 ,n8[47]);
    nand g2219(n1972 ,n1485 ,n1767);
    nand g2220(n96 ,n2331 ,n11[39]);
    nand g2221(n1689 ,n1332 ,n1493);
    dff g2222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2013), .Q(n6[0]));
    dff g2223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1832), .Q(n7[32]));
    or g2224(n1258 ,n7[28] ,n1187);
    nand g2225(n1426 ,n2270 ,n1289);
    or g2226(n1254 ,n7[5] ,n1191);
    nand g2227(n209 ,n33 ,n208);
    xnor g2228(n2351 ,n2076 ,n2[43]);
    xnor g2229(n2430 ,n983 ,n1116);
    nand g2230(n1827 ,n1410 ,n1622);
    nand g2231(n275 ,n39 ,n274);
    not g2232(n1135 ,n10[7]);
    nor g2233(n1864 ,n1651 ,n1815);
    xnor g2234(n2295 ,n167 ,n292);
    nand g2235(n1882 ,n1476 ,n1680);
    nand g2236(n1570 ,n2393 ,n1289);
    nor g2237(n875 ,n653 ,n874);
    xnor g2238(n714 ,n2[49] ,n2[113]);
    nand g2239(n1174 ,n1146 ,n1152);
    nand g2240(n547 ,n430 ,n546);
    xnor g2241(n2520 ,n2076 ,n2521);
    nand g2242(n1706 ,n1280 ,n1495);
    nand g2243(n531 ,n466 ,n530);
    xnor g2244(n2389 ,n1034 ,n993);
    xnor g2245(n2440 ,n2078 ,n2441);
    nor g2246(n1122 ,n896 ,n1121);
    dff g2247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1957), .Q(n8[16]));
    nand g2248(n1648 ,n1309 ,n1501);
    nand g2249(n231 ,n57 ,n230);
    nor g2250(n1101 ,n962 ,n1100);
    dff g2251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1936), .Q(n8[30]));
    xor g2252(n2373 ,n2436 ,n9[49]);
    or g2253(n1245 ,n7[11] ,n1186);
    nor g2254(n825 ,n651 ,n824);
    or g2255(n1291 ,n1 ,n1179);
    or g2256(n1257 ,n7[2] ,n1193);
    xnor g2257(n2396 ,n958 ,n1048);
    xnor g2258(n2174 ,n616 ,n471);
    xnor g2259(n2369 ,n2[61] ,n2075);
    nor g2260(n903 ,n2496 ,n11[46]);
    xnor g2261(n4[53] ,n2102 ,n8[53]);
    xnor g2262(n2406 ,n961 ,n1068);
    dff g2263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1853), .Q(n7[15]));
    xnor g2264(n963 ,n11[34] ,n2440);
    xnor g2265(n972 ,n11[40] ,n2484);
    nor g2266(n816 ,n704 ,n815);
    nand g2267(n1900 ,n1515 ,n1699);
    dff g2268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1890), .Q(n6[46]));
    nand g2269(n1897 ,n1507 ,n1697);
    xnor g2270(n3[62] ,n2113 ,n7[62]);
    nor g2271(n920 ,n2518 ,n11[41]);
    xnor g2272(n4[56] ,n2108 ,n8[56]);
    or g2273(n1218 ,n8[41] ,n1185);
    xnor g2274(n2400 ,n950 ,n1056);
    xnor g2275(n2543 ,n701 ,n859);
    nand g2276(n211 ,n16 ,n210);
    nand g2277(n606 ,n364 ,n605);
    dff g2278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1859), .Q(n7[10]));
    dff g2279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1932), .Q(n6[31]));
    nand g2280(n245 ,n64 ,n244);
    nand g2281(n255 ,n70 ,n254);
    nand g2282(n1740 ,n1369 ,n1499);
    xnor g2283(n2164 ,n596 ,n401);
    or g2284(n63 ,n2348 ,n11[40]);
    xnor g2285(n2159 ,n586 ,n489);
    not g2286(n440 ,n439);
    xnor g2287(n2382 ,n980 ,n1020);
    xnor g2288(n2242 ,n2[126] ,n2064);
    xnor g2289(n2313 ,n2066 ,n2[5]);
    or g2290(n1230 ,n8[42] ,n1198);
    or g2291(n1264 ,n6[61] ,n1188);
    xnor g2292(n5[11] ,n2105 ,n6[11]);
    nand g2293(n368 ,n2198 ,n11[35]);
    xnor g2294(n2349 ,n2071 ,n2[41]);
    xnor g2295(n954 ,n11[46] ,n2528);
    nor g2296(n888 ,n2472 ,n11[34]);
    dff g2297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1866), .Q(n7[4]));
    nand g2298(n1449 ,n2253 ,n1289);
    xnor g2299(n2316 ,n2070 ,n2[8]);
    nand g2300(n2058 ,n2023 ,n2041);
    xnor g2301(n2236 ,n2[120] ,n2070);
    nor g2302(n1295 ,n1 ,n1175);
    or g2303(n1262 ,n6[63] ,n1194);
    xnor g2304(n413 ,n11[34] ,n2229);
    nand g2305(n1842 ,n1432 ,n1641);
    nand g2306(n526 ,n356 ,n525);
    xnor g2307(n712 ,n2[2] ,n2[66]);
    nand g2308(n1811 ,n6[0] ,n1494);
    xnor g2309(n4[44] ,n2109 ,n8[44]);
    dff g2310(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1881), .Q(n6[54]));
    nor g2311(n922 ,n2476 ,n11[36]);
    xnor g2312(n948 ,n11[46] ,n2496);
    xnor g2313(n735 ,n2[14] ,n2[78]);
    xnor g2314(n4[6] ,n2104 ,n8[6]);
    nand g2315(n1481 ,n2563 ,n1293);
    nor g2316(n869 ,n668 ,n868);
    xor g2317(n2375 ,n963 ,n1006);
    nand g2318(n1856 ,n1445 ,n1658);
    nor g2319(n784 ,n719 ,n783);
    xnor g2320(n2215 ,n2[99] ,n2078);
    nor g2321(n639 ,n2[6] ,n2[70]);
    nand g2322(n1804 ,n1383 ,n1497);
    nor g2323(n870 ,n716 ,n869);
    nand g2324(n2082 ,n10[14] ,n11[46]);
    nand g2325(n754 ,n689 ,n708);
    xnor g2326(n2332 ,n2070 ,n2[24]);
    xnor g2327(n941 ,n11[33] ,n2438);
    nand g2328(n1562 ,n2139 ,n1289);
    nand g2329(n2089 ,n10[15] ,n11[31]);
    xnor g2330(n980 ,n11[41] ,n2454);
    xnor g2331(n2513 ,n736 ,n829);
    nand g2332(n2043 ,n10[2] ,n2031);
    dff g2333(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2061), .Q(n10[2]));
    nor g2334(n1185 ,n1130 ,n1155);
    not g2335(n422 ,n421);
    xnor g2336(n2403 ,n948 ,n1062);
    nor g2337(n809 ,n665 ,n808);
    xnor g2338(n168 ,n11[36] ,n2360);
    or g2339(n1287 ,n6[5] ,n1191);
    nand g2340(n2029 ,n9[50] ,n1914);
    nand g2341(n1671 ,n1262 ,n1493);
    nand g2342(n1688 ,n1336 ,n1493);
    nor g2343(n651 ,n2[36] ,n2[100]);
    nor g2344(n780 ,n735 ,n779);
    nand g2345(n1181 ,n1147 ,n1148);
    nand g2346(n120 ,n2347 ,n11[39]);
    nand g2347(n249 ,n41 ,n248);
    nor g2348(n1092 ,n932 ,n1091);
    xnor g2349(n192 ,n11[43] ,n2335);
    or g2350(n1356 ,n8[3] ,n1199);
    nor g2351(n670 ,n2[21] ,n2[85]);
    nand g2352(n1433 ,n2264 ,n1289);
    xnor g2353(n5[38] ,n2104 ,n6[38]);
    or g2354(n1238 ,n7[17] ,n1190);
    xnor g2355(n2154 ,n576 ,n447);
    nand g2356(n1896 ,n1504 ,n1693);
    nand g2357(n91 ,n2329 ,n11[37]);
    nand g2358(n545 ,n498 ,n544);
    xnor g2359(n985 ,n2460 ,n11[44]);
    xnor g2360(n2348 ,n2070 ,n2[40]);
    nand g2361(n1528 ,n2132 ,n1289);
    or g2362(n1276 ,n6[51] ,n1199);
    nor g2363(n1047 ,n1004 ,n1046);
    nor g2364(n834 ,n742 ,n833);
    nor g2365(n1057 ,n950 ,n1056);
    xnor g2366(n465 ,n11[32] ,n2195);
    nand g2367(n1567 ,n2420 ,n1289);
    xor g2368(n2114 ,n9[49] ,n2086);
    xnor g2369(n384 ,n11[32] ,n2227);
    nand g2370(n2027 ,n9[49] ,n1914);
    not g2371(n2066 ,n9[53]);
    xnor g2372(n2490 ,n2079 ,n2491);
    nor g2373(n846 ,n697 ,n845);
    xnor g2374(n3[12] ,n2109 ,n7[12]);
    xnor g2375(n2339 ,n2072 ,n2[31]);
    xnor g2376(n953 ,n11[40] ,n2548);
    nand g2377(n1527 ,n2407 ,n1289);
    dff g2378(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1874), .Q(n6[60]));
    not g2379(n472 ,n471);
    dff g2380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1972), .Q(n8[8]));
    or g2381(n1336 ,n8[63] ,n1194);
    nand g2382(n1831 ,n1415 ,n1629);
    nand g2383(n1471 ,n12[1] ,n1295);
    nand g2384(n1643 ,n1229 ,n1500);
    nand g2385(n1819 ,n1403 ,n1618);
    or g2386(n20 ,n2315 ,n11[39]);
    xnor g2387(n2279 ,n152 ,n260);
    nor g2388(n865 ,n682 ,n864);
    not g2389(n2077 ,n9[58]);
    nand g2390(n122 ,n2363 ,n11[39]);
    dff g2391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1821), .Q(n7[40]));
    nand g2392(n226 ,n81 ,n225);
    xnor g2393(n743 ,n2[18] ,n2[82]);
    nand g2394(n217 ,n22 ,n216);
    xnor g2395(n2146 ,n560 ,n395);
    nor g2396(n1064 ,n903 ,n1063);
    nand g2397(n278 ,n92 ,n277);
    nand g2398(n1958 ,n1563 ,n1757);
    or g2399(n50 ,n2353 ,n11[45]);
    or g2400(n1369 ,n6[28] ,n1187);
    nand g2401(n1817 ,n1546 ,n1715);
    xnor g2402(n2121 ,n510 ,n433);
    nand g2403(n1887 ,n1402 ,n1689);
    xnor g2404(n960 ,n11[38] ,n2544);
    or g2405(n23 ,n2357 ,n11[33]);
    nand g2406(n1973 ,n1576 ,n1768);
    nor g2407(n845 ,n672 ,n844);
    nand g2408(n1522 ,n2410 ,n1289);
    nor g2409(n912 ,n2460 ,n11[44]);
    nand g2410(n1941 ,n1544 ,n1739);
    nor g2411(n867 ,n649 ,n866);
    nand g2412(n2080 ,n9[49] ,n10[0]);
    or g2413(n53 ,n2351 ,n11[43]);
    dff g2414(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1947), .Q(n6[27]));
    nor g2415(n1814 ,n13[0] ,n1401);
    xnor g2416(n2144 ,n556 ,n397);
    xnor g2417(n2150 ,n568 ,n423);
    nand g2418(n127 ,n2357 ,n11[33]);
    xnor g2419(n2099 ,n2072 ,n2081);
    nor g2420(n1191 ,n1131 ,n1155);
    xnor g2421(n2134 ,n536 ,n479);
    xnor g2422(n5[3] ,n2112 ,n6[3]);
    nand g2423(n1784 ,n1363 ,n1497);
    nor g2424(n668 ,n2[58] ,n2[122]);
    nand g2425(n1769 ,n1388 ,n1495);
    dff g2426(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1948), .Q(n6[26]));
    or g2427(n1362 ,n7[60] ,n1187);
    xnor g2428(n2363 ,n2074 ,n2[55]);
    xnor g2429(n5[6] ,n2104 ,n6[6]);
    xnor g2430(n2495 ,n696 ,n811);
    nor g2431(n1496 ,n1171 ,n1291);
    xnor g2432(n2544 ,n2545 ,n2074);
    nand g2433(n210 ,n79 ,n209);
    xor g2434(n2112 ,n9[51] ,n2097);
    nand g2435(n1577 ,n2177 ,n1289);
    nand g2436(n2016 ,n9[61] ,n1914);
    nor g2437(n781 ,n677 ,n780);
    nand g2438(n595 ,n385 ,n594);
    nor g2439(n1173 ,n9[56] ,n1155);
    xnor g2440(n417 ,n11[46] ,n2225);
    buf g2441(n1289 ,n1290);
    nand g2442(n44 ,n2319 ,n11[43]);
    xnor g2443(n2185 ,n2[69] ,n2066);
    xnor g2444(n135 ,n11[31] ,n2339);
    nor g2445(n1150 ,n10[6] ,n10[7]);
    nand g2446(n2096 ,n10[4] ,n11[36]);
    nor g2447(n884 ,n2490 ,n11[43]);
    xnor g2448(n5[36] ,n2100 ,n6[36]);
    dff g2449(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1895), .Q(n8[58]));
    xnor g2450(n2445 ,n720 ,n761);
    nor g2451(n1096 ,n889 ,n1095);
    nand g2452(n1846 ,n1431 ,n1646);
    xnor g2453(n501 ,n11[39] ,n2234);
    xnor g2454(n958 ,n11[39] ,n2482);
    dff g2455(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1962), .Q(n8[44]));
    nor g2456(n908 ,n2474 ,n11[35]);
    nand g2457(n1661 ,n1249 ,n1486);
    xnor g2458(n726 ,n2[9] ,n2[73]);
    xnor g2459(n2131 ,n530 ,n465);
    dff g2460(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1869), .Q(n7[1]));
    xnor g2461(n696 ,n2[30] ,n2[94]);
    xnor g2462(n4[42] ,n2101 ,n8[42]);
    xnor g2463(n2550 ,n2077 ,n2551);
    nand g2464(n1557 ,n2135 ,n1289);
    dff g2465(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1854), .Q(n7[14]));
    nand g2466(n1785 ,n1360 ,n1498);
    nand g2467(n2032 ,n10[15] ,n2031);
    nand g2468(n1796 ,n1375 ,n1490);
    xnor g2469(n473 ,n11[34] ,n2197);
    nand g2470(n1417 ,n2156 ,n1289);
    nand g2471(n296 ,n95 ,n295);
    nand g2472(n1614 ,n2426 ,n1289);
    nand g2473(n1965 ,n1509 ,n1763);
    nand g2474(n1444 ,n2257 ,n1289);
    nand g2475(n350 ,n2189 ,n11[42]);
    xnor g2476(n3[33] ,n2114 ,n7[33]);
    or g2477(n1387 ,n7[43] ,n1186);
    xnor g2478(n2346 ,n2069 ,n2[38]);
    nand g2479(n611 ,n416 ,n610);
    nand g2480(n2009 ,n1451 ,n1714);
    xnor g2481(n2238 ,n2[122] ,n2077);
    xnor g2482(n2436 ,n2073 ,n2437);
    dff g2483(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1999), .Q(n7[52]));
    xnor g2484(n4[1] ,n2114 ,n8[1]);
    nand g2485(n11[45] ,n2064 ,n2079);
    nand g2486(n1532 ,n2153 ,n1289);
    xnor g2487(n4[55] ,n2106 ,n8[55]);
    nor g2488(n835 ,n662 ,n834);
    xnor g2489(n451 ,n11[44] ,n2207);
    or g2490(n1391 ,n7[0] ,n1292);
    xnor g2491(n2253 ,n165 ,n208);
    xnor g2492(n2380 ,n976 ,n1016);
    nand g2493(n529 ,n464 ,n528);
    or g2494(n1200 ,n1181 ,n1182);
    nand g2495(n1872 ,n1463 ,n1672);
    nand g2496(n1963 ,n1566 ,n1759);
    xnor g2497(n2426 ,n1000 ,n1108);
    dff g2498(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1992), .Q(n7[56]));
    nand g2499(n1697 ,n1307 ,n1486);
    xnor g2500(n3[25] ,n2111 ,n7[25]);
    xnor g2501(n2293 ,n164 ,n288);
    xnor g2502(n2275 ,n135 ,n252);
    nand g2503(n1653 ,n1390 ,n1494);
    nand g2504(n324 ,n2209 ,n11[46]);
    nand g2505(n361 ,n2182 ,n11[35]);
    nor g2506(n667 ,n2[20] ,n2[84]);
    nor g2507(n664 ,n2[62] ,n2[126]);
    xnor g2508(n2335 ,n2076 ,n2[27]);
    nand g2509(n1628 ,n1214 ,n1491);
    nand g2510(n1774 ,n1355 ,n1490);
    dff g2511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1844), .Q(n7[22]));
    xnor g2512(n2564 ,n14[10] ,n14[12]);
    or g2513(n1330 ,n8[24] ,n1195);
    or g2514(n1314 ,n8[15] ,n1194);
    xnor g2515(n2122 ,n512 ,n390);
    xnor g2516(n2460 ,n2075 ,n2461);
    nand g2517(n590 ,n378 ,n589);
    xnor g2518(n2186 ,n2[70] ,n2069);
    xnor g2519(n2263 ,n189 ,n228);
    nor g2520(n654 ,n2[39] ,n2[103]);
    nand g2521(n305 ,n61 ,n304);
    nand g2522(n558 ,n318 ,n557);
    not g2523(n1176 ,n1175);
    nor g2524(n686 ,n2[4] ,n2[68]);
    xor g2525(n2179 ,n2243 ,n626);
    not g2526(n464 ,n463);
    xnor g2527(n2364 ,n2070 ,n2[56]);
    xnor g2528(n2482 ,n2483 ,n2070);
    nor g2529(n1163 ,n9[55] ,n1155);
    xnor g2530(n2165 ,n598 ,n413);
    nor g2531(n901 ,n2550 ,n11[41]);
    dff g2532(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2011), .Q(n8[13]));
    nor g2533(n1046 ,n927 ,n1045);
    xnor g2534(n3[60] ,n2109 ,n7[60]);
    nand g2535(n1955 ,n1615 ,n1751);
    nand g2536(n1989 ,n1592 ,n1787);
    xnor g2537(n2182 ,n2[66] ,n2068);
    nand g2538(n232 ,n88 ,n231);
    nand g2539(n2018 ,n9[59] ,n1914);
    nand g2540(n1799 ,n1377 ,n1491);
    dff g2541(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1994), .Q(n6[13]));
    nand g2542(n271 ,n63 ,n270);
    nand g2543(n99 ,n2352 ,n11[44]);
    xnor g2544(n431 ,n11[45] ,n2240);
    nand g2545(n1596 ,n2145 ,n1289);
    dff g2546(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2055), .Q(n10[12]));
    nand g2547(n1790 ,n1368 ,n1489);
    xnor g2548(n2450 ,n2451 ,n2070);
    xnor g2549(n2130 ,n528 ,n463);
    xnor g2550(n2187 ,n2[71] ,n2074);
    dff g2551(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1857), .Q(n6[1]));
    xnor g2552(n3[55] ,n2106 ,n7[55]);
    nor g2553(n796 ,n750 ,n795);
    xnor g2554(n403 ,n11[44] ,n2239);
    nand g2555(n625 ,n484 ,n624);
    nor g2556(n1060 ,n882 ,n1059);
    nor g2557(n832 ,n711 ,n831);
    nand g2558(n1549 ,n2400 ,n1289);
    dff g2559(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[14]), .Q(n9[62]));
    xnor g2560(n455 ,n11[40] ,n2219);
    xnor g2561(n2289 ,n140 ,n280);
    nor g2562(n676 ,n2[26] ,n2[90]);
    nor g2563(n1033 ,n992 ,n1032);
    nand g2564(n555 ,n452 ,n554);
    nand g2565(n1666 ,n1255 ,n1490);
    nand g2566(n1476 ,n2425 ,n1289);
    xnor g2567(n738 ,n2[58] ,n2[122]);
    nand g2568(n1891 ,n1577 ,n1692);
    not g2569(n1136 ,n10[13]);
    or g2570(n1341 ,n8[13] ,n1188);
    nand g2571(n2060 ,n2026 ,n2045);
    or g2572(n1266 ,n6[60] ,n1187);
    nor g2573(n774 ,n730 ,n773);
    nand g2574(n1507 ,n2173 ,n1289);
    not g2575(n2074 ,n9[55]);
    xnor g2576(n4[41] ,n2111 ,n8[41]);
    nor g2577(n787 ,n657 ,n786);
    nand g2578(n1670 ,n1391 ,n1494);
    nand g2579(n1016 ,n937 ,n1015);
    nand g2580(n589 ,n496 ,n588);
    nand g2581(n107 ,n2335 ,n11[43]);
    xnor g2582(n2421 ,n943 ,n1098);
    xnor g2583(n2477 ,n748 ,n793);
    xnor g2584(n2243 ,n2[127] ,n2072);
    nand g2585(n1878 ,n9[48] ,n1654);
    dff g2586(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1886), .Q(n6[49]));
    nand g2587(n352 ,n2190 ,n11[43]);
    nor g2588(n669 ,n2[44] ,n2[108]);
    xnor g2589(n2202 ,n2[86] ,n2069);
    nand g2590(n1442 ,n2117 ,n1289);
    nor g2591(n1010 ,n935 ,n1009);
    dff g2592(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[7]), .Q(n9[55]));
    xnor g2593(n148 ,n11[45] ,n2337);
    xnor g2594(n1004 ,n11[38] ,n2480);
    nor g2595(n1073 ,n969 ,n1072);
    nand g2596(n549 ,n412 ,n548);
    nand g2597(n1893 ,n1535 ,n1732);
    nor g2598(n1175 ,n13[1] ,n1151);
    xnor g2599(n2137 ,n542 ,n491);
    xnor g2600(n2307 ,n2371 ,n316);
    nor g2601(n1028 ,n912 ,n1027);
    nand g2602(n1987 ,n1593 ,n1784);
    nand g2603(n242 ,n100 ,n241);
    xnor g2604(n4[3] ,n2112 ,n8[3]);
    nor g2605(n914 ,n2456 ,n11[42]);
    dff g2606(.RN(n2567), .SN(1'b1), .CK(n0), .D(n14[0]), .Q(n9[48]));
    dff g2607(.RN(n2567), .SN(1'b1), .CK(n0), .D(n9[55]), .Q(n9[56]));
    xnor g2608(n2546 ,n2070 ,n2547);
    nand g2609(n1523 ,n2160 ,n1289);
    nand g2610(n1991 ,n1595 ,n1789);
    nand g2611(n571 ,n428 ,n570);
    xnor g2612(n2330 ,n2069 ,n2[22]);
    or g2613(n1385 ,n7[55] ,n1189);
    nand g2614(n1553 ,n2398 ,n1289);
    nand g2615(n1470 ,n2427 ,n1289);
    xnor g2616(n2218 ,n2[102] ,n2069);
    xnor g2617(n3[24] ,n2108 ,n7[24]);
    xnor g2618(n3[59] ,n2105 ,n7[59]);
    nand g2619(n1644 ,n1235 ,n1492);
    nand g2620(n266 ,n123 ,n265);
    xnor g2621(n2345 ,n2066 ,n2[37]);
    nand g2622(n1408 ,n2282 ,n1289);
    xnor g2623(n2514 ,n2070 ,n2515);
    xnor g2624(n2151 ,n570 ,n427);
    nand g2625(n1889 ,n1543 ,n1690);
    nand g2626(n1768 ,n1350 ,n1500);
    or g2627(n1381 ,n6[10] ,n1198);
    nand g2628(n2088 ,n10[0] ,n11[32]);
    xnor g2629(n999 ,n11[35] ,n2474);
    nand g2630(n2013 ,n1878 ,n1864);
    nand g2631(n1783 ,n1220 ,n1497);
    nand g2632(n1838 ,n1424 ,n1637);
    nand g2633(n1602 ,n2384 ,n1289);
    nand g2634(n131 ,n2341 ,n11[33]);
    xnor g2635(n4[52] ,n2100 ,n8[52]);
    or g2636(n25 ,n2367 ,n11[43]);
    or g2637(n1272 ,n6[53] ,n1191);
    nand g2638(n593 ,n494 ,n592);
    nand g2639(n1546 ,n2287 ,n1289);
    nand g2640(n523 ,n450 ,n522);
    nor g2641(n799 ,n630 ,n798);
    nand g2642(n1760 ,n1341 ,n1498);
    xnor g2643(n2553 ,n716 ,n869);
    xnor g2644(n4[7] ,n2106 ,n8[7]);
    nand g2645(n1646 ,n1232 ,n1488);
    xnor g2646(n2177 ,n622 ,n499);
    xnor g2647(n2205 ,n2[89] ,n2071);
    nor g2648(n833 ,n636 ,n832);
    not g2649(n315 ,n314);
    or g2650(n1353 ,n8[5] ,n1191);
    xnor g2651(n2227 ,n2[111] ,n2072);
    dff g2652(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2008), .Q(n7[44]));
    xnor g2653(n3[10] ,n2101 ,n7[10]);
    xnor g2654(n2402 ,n945 ,n1060);
    xnor g2655(n2257 ,n146 ,n216);
    xnor g2656(n2269 ,n190 ,n240);
    xnor g2657(n489 ,n11[44] ,n2223);
    or g2658(n1378 ,n6[11] ,n1186);
    nand g2659(n2038 ,n10[9] ,n2031);
    not g2660(n478 ,n477);
    nand g2661(n542 ,n374 ,n541);
    nand g2662(n1635 ,n1382 ,n1498);
    xnor g2663(n945 ,n11[45] ,n2494);
    dff g2664(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1833), .Q(n7[31]));
    xnor g2665(n2225 ,n2[109] ,n2075);
    dff g2666(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1976), .Q(n8[4]));
    nand g2667(n2042 ,n10[0] ,n2031);
    nand g2668(n84 ,n2326 ,n11[34]);
    dff g2669(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2049), .Q(n10[14]));
    nand g2670(n1506 ,n2174 ,n1289);
    or g2671(n1360 ,n7[61] ,n1188);
    dff g2672(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2051), .Q(n10[8]));
    not g2673(n2567 ,n1);
    nand g2674(n1912 ,n1519 ,n1712);
    nand g2675(n536 ,n367 ,n535);
    xnor g2676(n2277 ,n149 ,n256);
    dff g2677(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1959), .Q(n6[23]));
    nand g2678(n525 ,n454 ,n524);
    dff g2679(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1837), .Q(n7[28]));
    xnor g2680(n2505 ,n705 ,n821);
    dff g2681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1849), .Q(n7[19]));
    nand g2682(n2040 ,n10[7] ,n2031);
    nand g2683(n1410 ,n2379 ,n1289);
    nand g2684(n1513 ,n2413 ,n1289);
    nand g2685(n1692 ,n1337 ,n1498);
    nand g2686(n1984 ,n1588 ,n1783);
    or g2687(n59 ,n2330 ,n11[38]);
    nand g2688(n1684 ,n1279 ,n1491);
    dff g2689(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1965), .Q(n8[11]));
    or g2690(n17 ,n2314 ,n11[38]);
    nor g2691(n1198 ,n1133 ,n1155);
    nand g2692(n1529 ,n2175 ,n1289);
    nand g2693(n112 ,n2362 ,n11[38]);
    or g2694(n31 ,n2356 ,n11[32]);
    nand g2695(n1609 ,n2292 ,n1289);
    xnor g2696(n5[8] ,n2108 ,n6[8]);
    xnor g2697(n2399 ,n959 ,n1054);
    xnor g2698(n2515 ,n711 ,n831);
    or g2699(n193 ,n133 ,n69);
    xnor g2700(n3[28] ,n2109 ,n7[28]);
    xnor g2701(n2433 ,n968 ,n1122);
    xnor g2702(n2317 ,n2071 ,n2[9]);
    nor g2703(n636 ,n2[40] ,n2[104]);
    nor g2704(n1186 ,n1134 ,n1155);
    nand g2705(n594 ,n379 ,n593);
    nor g2706(n1041 ,n999 ,n1040);
    xnor g2707(n189 ,n11[35] ,n2327);
    nand g2708(n1848 ,n1433 ,n1647);
    nand g2709(n1479 ,n2422 ,n1289);
    xnor g2710(n2286 ,n161 ,n274);
    nand g2711(n1969 ,n1575 ,n1771);
    not g2712(n1144 ,n10[6]);
    xnor g2713(n2230 ,n2[114] ,n2068);
    xnor g2714(n2358 ,n2068 ,n2[50]);
    or g2715(n1342 ,n6[21] ,n1191);
    nor g2716(n1032 ,n879 ,n1031);
    xnor g2717(n976 ,n11[39] ,n2450);
    dff g2718(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1901), .Q(n6[42]));
    nand g2719(n320 ,n2229 ,n11[34]);
    nand g2720(n11[44] ,n2075 ,n2076);
    xnor g2721(n2147 ,n562 ,n399);
    xnor g2722(n5[22] ,n2104 ,n6[22]);
    or g2723(n1398 ,n8[0] ,n1292);
    xnor g2724(n698 ,n2[26] ,n2[90]);
    xnor g2725(n2285 ,n160 ,n272);
    xnor g2726(n2302 ,n181 ,n306);
    or g2727(n1308 ,n8[44] ,n1187);
    xnor g2728(n3[49] ,n2114 ,n7[49]);
    dff g2729(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2004), .Q(n7[48]));
    nor g2730(n790 ,n745 ,n789);
    xnor g2731(n459 ,n11[37] ,n2232);
    xnor g2732(n2342 ,n2068 ,n2[34]);
    nand g2733(n1667 ,n1256 ,n1495);
    nand g2734(n563 ,n400 ,n562);
    nand g2735(n319 ,n2228 ,n11[33]);
    nor g2736(n1499 ,n1167 ,n1291);
    xor g2737(n2111 ,n9[57] ,n2083);
    nand g2738(n304 ,n124 ,n303);
    xnor g2739(n2557 ,n729 ,n873);
    nand g2740(n580 ,n336 ,n579);
    nand g2741(n1938 ,n1596 ,n1737);
    dff g2742(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1960), .Q(n6[48]));
    nand g2743(n527 ,n458 ,n526);
    xnor g2744(n2217 ,n2[101] ,n2066);
    nand g2745(n1806 ,n1386 ,n1499);
    xnor g2746(n179 ,n11[43] ,n2319);
    xnor g2747(n4[18] ,n2110 ,n8[18]);
    nor g2748(n877 ,n664 ,n876);
    nand g2749(n1793 ,n1385 ,n1500);
    nor g2750(n853 ,n644 ,n852);
    nand g2751(n1921 ,n1417 ,n1720);
    nand g2752(n1629 ,n1215 ,n1492);
    not g2753(n502 ,n501);
    xnor g2754(n2214 ,n2[98] ,n2068);
    xnor g2755(n4[54] ,n2104 ,n8[54]);
    xnor g2756(n1003 ,n11[43] ,n2522);
    xnor g2757(n2532 ,n2073 ,n2533);
    xnor g2758(n2258 ,n145 ,n218);
    dff g2759(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1974), .Q(n8[6]));
    nor g2760(n902 ,n2558 ,n11[45]);
    xnor g2761(n165 ,n11[41] ,n2317);
    nand g2762(n614 ,n337 ,n613);
    or g2763(n1252 ,n7[7] ,n1189);
    nand g2764(n1928 ,n1537 ,n1679);
    or g2765(n631 ,n2[1] ,n2[65]);
    nor g2766(n844 ,n692 ,n843);
    dff g2767(.RN(1'b1), .SN(n2567), .CK(n0), .D(n9[51]), .Q(n14[5]));
    nand g2768(n688 ,n2[2] ,n2[66]);
    xnor g2769(n2228 ,n2[112] ,n2067);
    xnor g2770(n175 ,n11[43] ,n2367);
    nand g2771(n1837 ,n1423 ,n1636);
    xnor g2772(n993 ,n2468 ,n11[32]);
    dff g2773(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1985), .Q(n6[15]));
    xor g2774(n2108 ,n9[56] ,n2087);
    or g2775(n1243 ,n7[13] ,n1188);
    nand g2776(n550 ,n322 ,n549);
    nand g2777(n1431 ,n2265 ,n1289);
    nor g2778(n874 ,n729 ,n873);
    xnor g2779(n3[22] ,n2104 ,n7[22]);
    nand g2780(n1580 ,n2138 ,n1289);
    nand g2781(n269 ,n36 ,n268);
    nand g2782(n1690 ,n1367 ,n1497);
    nand g2783(n1849 ,n1434 ,n1649);
    nand g2784(n1544 ,n2401 ,n1289);
    nor g2785(n1070 ,n891 ,n1069);
    xnor g2786(n3[2] ,n2110 ,n7[2]);
    xnor g2787(n4[13] ,n2103 ,n8[13]);
    xnor g2788(n965 ,n11[45] ,n2526);
    xnor g2789(n2469 ,n740 ,n785);
    nand g2790(n1930 ,n1534 ,n1726);
    or g2791(n1325 ,n6[46] ,n1192);
    nor g2792(n1025 ,n984 ,n1024);
    nand g2793(n1996 ,n1607 ,n1797);
    nand g2794(n196 ,n101 ,n195);
    xnor g2795(n2529 ,n697 ,n845);
    nand g2796(n274 ,n83 ,n273);
    not g2797(n410 ,n409);
    nand g2798(n2008 ,n1559 ,n1806);
    nand g2799(n125 ,n2315 ,n11[39]);
    or g2800(n1241 ,n7[15] ,n1194);
    nand g2801(n371 ,n2199 ,n11[36]);
    nand g2802(n362 ,n2235 ,n11[40]);
    nand g2803(n2053 ,n2019 ,n2037);
    nor g2804(n1063 ,n948 ,n1062);
    or g2805(n1207 ,n7[39] ,n1189);
    nor g2806(n836 ,n747 ,n835);
    nand g2807(n1457 ,n2248 ,n1289);
    xnor g2808(n5[29] ,n2103 ,n6[29]);
    xnor g2809(n164 ,n11[33] ,n2357);
    xnor g2810(n2203 ,n2[87] ,n2074);
    nor g2811(n1056 ,n880 ,n1055);
    nand g2812(n375 ,n2238 ,n11[43]);
    dff g2813(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1922), .Q(n8[39]));
    nand g2814(n1611 ,n2291 ,n1289);
    dff g2815(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1935), .Q(n8[31]));
    xnor g2816(n3[31] ,n2115 ,n7[31]);
    nand g2817(n237 ,n18 ,n236);
    or g2818(n1269 ,n6[56] ,n1195);
    nand g2819(n93 ,n2330 ,n11[38]);
    xnor g2820(n2153 ,n574 ,n386);
    dff g2821(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1928), .Q(n6[32]));
    nor g2822(n1100 ,n887 ,n1099);
    xnor g2823(n2235 ,n2[119] ,n2074);
    nor g2824(n1038 ,n919 ,n1037);
    or g2825(n27 ,n2363 ,n11[39]);
    nand g2826(n601 ,n381 ,n600);
    nor g2827(n685 ,n2[30] ,n2[94]);
    dff g2828(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1931), .Q(n8[34]));
    xnor g2829(n2305 ,n2369 ,n312);
    xnor g2830(n475 ,n11[43] ,n2222);
    xnor g2831(n720 ,n2[5] ,n2[69]);
    nand g2832(n1904 ,n1512 ,n1705);
    or g2833(n1354 ,n6[17] ,n1190);
    xnor g2834(n2200 ,n2[84] ,n2065);
    xnor g2835(n445 ,n11[43] ,n2190);
    xnor g2836(n2472 ,n2078 ,n2473);
    nor g2837(n909 ,n2458 ,n11[43]);
    nand g2838(n1823 ,n1408 ,n1623);
    nand g2839(n1411 ,n2280 ,n1289);
    nand g2840(n334 ,n2213 ,n11[34]);
    xnor g2841(n2148 ,n564 ,n407);
    nand g2842(n1466 ,n2432 ,n1289);
    or g2843(n1364 ,n7[59] ,n1186);
    xnor g2844(n952 ,n2498 ,n11[31]);
    or g2845(n1393 ,n8[48] ,n1292);
    nand g2846(n524 ,n355 ,n523);
    or g2847(n1220 ,n7[62] ,n1192);
    nand g2848(n2025 ,n9[52] ,n1914);
    xnor g2849(n2418 ,n965 ,n1092);
    xnor g2850(n2467 ,n719 ,n783);
    xnor g2851(n745 ,n2[19] ,n2[83]);
    nand g2852(n503 ,n348 ,n422);
    xnor g2853(n163 ,n11[42] ,n2318);
    xnor g2854(n425 ,n11[36] ,n2183);
    nand g2855(n113 ,n2354 ,n11[46]);
    xnor g2856(n2447 ,n752 ,n763);
    nand g2857(n1750 ,n1334 ,n1490);
    nand g2858(n1415 ,n2277 ,n1289);
    dff g2859(.RN(1'b1), .SN(n2567), .CK(n0), .D(n14[10]), .Q(n14[11]));
    nand g2860(n1853 ,n1441 ,n1655);
    nand g2861(n1691 ,n1325 ,n1497);
    xnor g2862(n2169 ,n606 ,n481);
    nand g2863(n321 ,n2234 ,n11[39]);
    dff g2864(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1984), .Q(n7[62]));
    nor g2865(n1193 ,n1137 ,n1155);
    dff g2866(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1882), .Q(n6[53]));
    nand g2867(n346 ,n2188 ,n11[41]);
    xnor g2868(n2398 ,n951 ,n1052);
    xnor g2869(n2547 ,n709 ,n863);
    nand g2870(n1959 ,n1561 ,n1756);
    xnor g2871(n2542 ,n2069 ,n2543);
    nand g2872(n1583 ,n2118 ,n1289);
    or g2873(n1331 ,n6[25] ,n1185);
    nor g2874(n824 ,n724 ,n823);
    or g2875(n1229 ,n7[23] ,n1189);
    nor g2876(n1076 ,n900 ,n1075);
    nand g2877(n1566 ,n2394 ,n1289);
    nand g2878(n1940 ,n1584 ,n1777);
    not g2879(n1178 ,n1177);
    nand g2880(n360 ,n2220 ,n11[41]);
    xnor g2881(n2265 ,n187 ,n232);
    nor g2882(n868 ,n738 ,n867);
    xnor g2883(n2254 ,n163 ,n210);
    xnor g2884(n4[16] ,n2107 ,n8[16]);
    nand g2885(n1939 ,n1545 ,n1738);
    nand g2886(n276 ,n86 ,n275);
    dff g2887(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1919), .Q(n8[41]));
    nand g2888(n1767 ,n1349 ,n1489);
    or g2889(n30 ,n2334 ,n11[42]);
    xnor g2890(n2481 ,n753 ,n797);
    nand g2891(n76 ,n2322 ,n11[46]);
    dff g2892(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1888), .Q(n8[63]));
    xnor g2893(n2199 ,n2[83] ,n2078);
    nand g2894(n2081 ,n9[62] ,n10[15]);
    nand g2895(n1800 ,n1365 ,n1492);
    xnor g2896(n730 ,n2[11] ,n2[75]);
    or g2897(n1237 ,n7[18] ,n1193);
    nand g2898(n2063 ,n2025 ,n2046);
    not g2899(n430 ,n429);
    nand g2900(n359 ,n2194 ,n11[31]);
    xnor g2901(n3[27] ,n2105 ,n7[27]);
    nor g2902(n872 ,n710 ,n871);
    dff g2903(.RN(1'b1), .SN(n2567), .CK(n0), .D(n14[11]), .Q(n14[12]));
    nand g2904(n1413 ,n2155 ,n1289);
    or g2905(n1348 ,n8[9] ,n1185);
    nand g2906(n236 ,n93 ,n235);
    nor g2907(n1089 ,n1003 ,n1088);
    or g2908(n1323 ,n8[31] ,n1194);
    dff g2909(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1812), .Q(n12[2]));
    xnor g2910(n2340 ,n2067 ,n2[32]);
    xnor g2911(n2549 ,n721 ,n865);
    nand g2912(n374 ,n2200 ,n11[37]);
    dff g2913(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1997), .Q(n7[53]));
    nand g2914(n1610 ,n2429 ,n1289);
    xnor g2915(n2462 ,n2064 ,n2463);
    nand g2916(n345 ,n2187 ,n11[40]);
    xnor g2917(n4[23] ,n2106 ,n8[23]);
    nand g2918(n1710 ,n1393 ,n1494);
    nor g2919(n928 ,n2534 ,n11[33]);
    or g2920(n33 ,n2317 ,n11[41]);
    nand g2921(n2085 ,n10[12] ,n11[44]);
    nand g2922(n1017 ,n977 ,n1016);
    nand g2923(n605 ,n460 ,n604);
    or g2924(n34 ,n2323 ,n11[31]);
    xnor g2925(n169 ,n11[37] ,n2361);
    nor g2926(n1171 ,n9[58] ,n1155);
    not g2927(n404 ,n403);
    nand g2928(n1843 ,n1429 ,n1643);
    xnor g2929(n4[63] ,n2099 ,n8[63]);
    dff g2930(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1877), .Q(n6[57]));
    xnor g2931(n702 ,n2[24] ,n2[88]);
    nand g2932(n256 ,n111 ,n255);
    nor g2933(n1124 ,n925 ,n1123);
    or g2934(n1396 ,n8[16] ,n1292);
    or g2935(n48 ,n2349 ,n11[41]);
    nor g2936(n837 ,n643 ,n836);
    nor g2937(n660 ,n2[52] ,n2[116]);
    or g2938(n1208 ,n8[38] ,n1197);
    nor g2939(n792 ,n746 ,n791);
    nor g2940(n911 ,n2514 ,n11[39]);
    or g2941(n1212 ,n7[35] ,n1199);
    nand g2942(n132 ,n2321 ,n11[45]);
    xnor g2943(n3[19] ,n2112 ,n7[19]);
    nor g2944(n1501 ,n1170 ,n1291);
    nand g2945(n331 ,n2217 ,n11[38]);
    nand g2946(n1739 ,n1217 ,n1498);
    nor g2947(n1118 ,n901 ,n1117);
    or g2948(n1358 ,n7[63] ,n1194);
    or g2949(n1260 ,n8[47] ,n1194);
    xnor g2950(n4[14] ,n2113 ,n8[14]);
    xnor g2951(n3[34] ,n2110 ,n7[34]);
    xnor g2952(n711 ,n2[40] ,n2[104]);
    xnor g2953(n2504 ,n2078 ,n2505);
    nand g2954(n118 ,n2355 ,n11[31]);
    xnor g2955(n1002 ,n11[42] ,n2552);
    nor g2956(n808 ,n693 ,n807);
    xnor g2957(n4[35] ,n2112 ,n8[35]);
    dff g2958(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1880), .Q(n6[55]));
    or g2959(n1347 ,n6[20] ,n1196);
    nand g2960(n1625 ,n1213 ,n1487);
    xnor g2961(n5[57] ,n2111 ,n6[57]);
    nor g2962(n907 ,n2546 ,n11[39]);
    xnor g2963(n5[49] ,n2114 ,n6[49]);
    or g2964(n36 ,n2347 ,n11[39]);
    dff g2965(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1971), .Q(n6[20]));
    nor g2966(n311 ,n2368 ,n310);
    xnor g2967(n2493 ,n691 ,n809);
    nand g2968(n1742 ,n1328 ,n1486);
    dff g2969(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2000), .Q(n7[51]));
    nor g2970(n1105 ,n994 ,n1104);
    nand g2971(n2090 ,n10[7] ,n11[39]);
    nor g2972(n887 ,n2532 ,n11[32]);
    or g2973(n1374 ,n7[53] ,n1191);
    xnor g2974(n2359 ,n2078 ,n2[51]);
    xnor g2975(n477 ,n11[43] ,n2206);
    xnor g2976(n423 ,n11[35] ,n2214);
    nand g2977(n1855 ,n1444 ,n1657);
    xnor g2978(n2262 ,n186 ,n226);
    dff g2979(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1929), .Q(n8[35]));
    nor g2980(n775 ,n680 ,n774);
    or g2981(n71 ,n2359 ,n11[35]);
    dff g2982(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1825), .Q(n7[37]));
    or g2983(n1351 ,n6[18] ,n1193);
    nand g2984(n1460 ,n2245 ,n1289);
    xnor g2985(n3[32] ,n2107 ,n7[32]);
    xnor g2986(n2124 ,n516 ,n382);
    dff g2987(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1964), .Q(n8[12]));
    nand g2988(n1883 ,n1479 ,n1684);
    nand g2989(n212 ,n130 ,n211);
    nand g2990(n620 ,n323 ,n619);
    nand g2991(n2019 ,n9[58] ,n1914);
    xnor g2992(n5[55] ,n2106 ,n6[55]);
    nor g2993(n1051 ,n972 ,n1050);
    nand g2994(n1754 ,n1319 ,n1492);
    or g2995(n1244 ,n7[12] ,n1187);
    xnor g2996(n2264 ,n154 ,n230);
    nand g2997(n615 ,n440 ,n614);
    dff g2998(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1912), .Q(n8[47]));
    xnor g2999(n3[42] ,n2101 ,n7[42]);
    nand g3000(n617 ,n472 ,n616);
    or g3001(n1285 ,n6[33] ,n1190);
endmodule
