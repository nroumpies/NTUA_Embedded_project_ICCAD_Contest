module top (n0, n1, n2, n3);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3;
    wire [63:0] n4;
    wire [15:0] n5;
    wire [7:0] n6;
    wire [7:0] n7;
    wire [7:0] n8;
    wire [3:0] n9;
    wire [15:0] n10;
    wire [3:0] n11;
    wire [31:0] n12;
    wire [3:0] n13;
    wire [7:0] n14;
    wire [15:0] n15;
    wire [63:0] n16;
    wire [19:0] n17;
    wire n18, n19, n20, n21, n22, n23, n24, n25;
    wire n26, n27, n28, n29, n30, n31, n32, n33;
    wire n34, n35, n36, n37, n38, n39, n40, n41;
    wire n42, n43, n44, n45, n46, n47, n48, n49;
    wire n50, n51, n52, n53, n54, n55, n56, n57;
    wire n58, n59, n60, n61, n62, n63, n64, n65;
    wire n66, n67, n68, n69, n70, n71, n72, n73;
    wire n74, n75, n76, n77, n78, n79, n80, n81;
    wire n82, n83, n84, n85, n86, n87, n88, n89;
    wire n90, n91, n92, n93, n94, n95, n96, n97;
    wire n98, n99, n100, n101, n102, n103, n104, n105;
    wire n106, n107, n108, n109, n110, n111, n112, n113;
    wire n114, n115, n116, n117, n118, n119, n120, n121;
    wire n122, n123, n124, n125, n126, n127, n128, n129;
    wire n130, n131, n132, n133, n134, n135, n136, n137;
    wire n138, n139, n140, n141, n142, n143, n144, n145;
    wire n146, n147, n148, n149, n150, n151, n152, n153;
    wire n154, n155, n156, n157, n158, n159, n160, n161;
    wire n162, n163, n164, n165, n166, n167, n168, n169;
    wire n170, n171, n172, n173, n174, n175, n176, n177;
    wire n178, n179, n180, n181, n182, n183, n184, n185;
    wire n186, n187, n188, n189, n190, n191, n192, n193;
    wire n194, n195, n196, n197, n198, n199, n200, n201;
    wire n202, n203, n204, n205, n206, n207, n208, n209;
    wire n210, n211, n212, n213, n214, n215, n216, n217;
    wire n218, n219, n220, n221, n222, n223, n224, n225;
    wire n226, n227, n228, n229, n230, n231, n232, n233;
    wire n234, n235, n236, n237, n238, n239, n240, n241;
    wire n242, n243, n244, n245, n246, n247, n248, n249;
    wire n250, n251, n252, n253, n254, n255, n256, n257;
    wire n258, n259, n260, n261, n262, n263, n264, n265;
    wire n266, n267, n268, n269, n270, n271, n272, n273;
    wire n274, n275, n276, n277, n278, n279, n280, n281;
    wire n282, n283, n284, n285, n286, n287, n288, n289;
    wire n290, n291, n292, n293, n294, n295, n296, n297;
    wire n298, n299, n300, n301, n302, n303, n304, n305;
    wire n306, n307, n308, n309, n310, n311, n312, n313;
    wire n314, n315, n316, n317, n318, n319, n320, n321;
    wire n322, n323, n324, n325, n326, n327, n328, n329;
    wire n330, n331, n332, n333, n334, n335, n336, n337;
    wire n338, n339, n340, n341, n342, n343, n344, n345;
    wire n346, n347, n348, n349, n350, n351, n352, n353;
    wire n354, n355, n356, n357, n358, n359, n360, n361;
    wire n362, n363, n364, n365, n366, n367, n368, n369;
    wire n370, n371, n372, n373, n374, n375, n376, n377;
    wire n378, n379, n380, n381, n382, n383, n384, n385;
    wire n386, n387, n388, n389, n390, n391, n392, n393;
    wire n394, n395, n396, n397, n398, n399, n400, n401;
    wire n402, n403, n404, n405, n406, n407, n408, n409;
    wire n410, n411, n412, n413, n414, n415, n416, n417;
    wire n418, n419, n420, n421, n422, n423, n424, n425;
    wire n426, n427, n428, n429, n430, n431, n432, n433;
    wire n434, n435, n436, n437, n438, n439, n440, n441;
    dff g0(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n217), .Q(n10[2]));
    dff g1(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n419), .Q(n17[17]));
    buf g2(n3[26], n3[31]);
    nand g3(n181 ,n8[0] ,n381);
    nand g4(n225 ,n1 ,n165);
    not g5(n144 ,n11[2]);
    buf g6(n3[10], n3[15]);
    nor g7(n115 ,n10[13] ,n114);
    buf g8(n3[6], n3[7]);
    buf g9(n3[51], n3[55]);
    not g10(n145 ,n15[0]);
    or g11(n415 ,n17[5] ,n1);
    nand g12(n324 ,n16[15] ,n310);
    nor g13(n426 ,n408 ,n1);
    nand g14(n53 ,n15[1] ,n15[0]);
    dff g15(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n304), .Q(n9[2]));
    dff g16(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n335), .Q(n4[48]));
    dff g17(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n209), .Q(n10[11]));
    nor g18(n42 ,n33 ,n40);
    dff g19(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n263), .Q(n15[1]));
    nand g20(n54 ,n15[5] ,n15[4]);
    nand g21(n76 ,n15[6] ,n75);
    not g22(n65 ,n15[12]);
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n338), .Q(n4[16]));
    not g24(n82 ,n81);
    buf g25(n3[62], n3[63]);
    buf g26(n3[46], n3[47]);
    dff g27(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n417), .Q(n17[0]));
    nor g28(n306 ,n11[3] ,n297);
    nor g29(n52 ,n15[11] ,n15[10]);
    buf g30(n3[19], n3[23]);
    nor g31(n40 ,n10[1] ,n37);
    or g32(n412 ,n17[8] ,n1);
    nor g33(n47 ,n41 ,n46);
    nor g34(n206 ,n125 ,n162);
    nor g35(n184 ,n149 ,n123);
    xnor g36(n391 ,n15[7] ,n76);
    not g37(n404 ,n17[18]);
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n215), .Q(n10[5]));
    nor g39(n19 ,n15[15] ,n15[14]);
    xor g40(n434 ,n2[5] ,n17[5]);
    or g41(n416 ,n17[16] ,n1);
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n303), .Q(n9[1]));
    nor g43(n439 ,n437 ,n436);
    not g44(n408 ,n17[19]);
    not g45(n314 ,n313);
    or g46(n43 ,n10[4] ,n42);
    or g47(n280 ,n9[0] ,n272);
    nand g48(n285 ,n380 ,n273);
    nor g49(n337 ,n312 ,n325);
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n266), .Q(n15[14]));
    buf g51(n3[12], n3[15]);
    xnor g52(n388 ,n15[10] ,n81);
    nor g53(n34 ,n10[13] ,n10[12]);
    or g54(n159 ,n8[0] ,n361);
    not g55(n407 ,n17[10]);
    not g56(n117 ,n116);
    nor g57(n251 ,n168 ,n225);
    xor g58(n431 ,n2[0] ,n17[0]);
    not g59(n400 ,n17[2]);
    buf g60(n3[38], n3[39]);
    or g61(n195 ,n183 ,n159);
    not g62(n129 ,n370);
    nor g63(n208 ,n129 ,n162);
    nand g64(n441 ,n438 ,n440);
    xnor g65(n356 ,n359 ,n354);
    nor g66(n66 ,n15[1] ,n15[0]);
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n434), .Q(n16[47]));
    nor g68(n36 ,n10[15] ,n10[14]);
    or g69(n321 ,n16[23] ,n309);
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n411), .Q(n17[8]));
    nand g71(n242 ,n144 ,n178);
    nand g72(n295 ,n9[1] ,n288);
    nor g73(n221 ,n135 ,n162);
    nor g74(n310 ,n123 ,n306);
    nand g75(n237 ,n390 ,n164);
    or g76(n256 ,n180 ,n193);
    nor g77(n190 ,n10[0] ,n162);
    nand g78(n57 ,n48 ,n53);
    buf g79(n3[14], n3[15]);
    nor g80(n155 ,n142 ,n377);
    nand g81(n327 ,n16[55] ,n310);
    nand g82(n283 ,n378 ,n273);
    nor g83(n107 ,n92 ,n106);
    xnor g84(n350 ,n347 ,n8[0]);
    nand g85(n336 ,n326 ,n323);
    buf g86(n3[1], n3[7]);
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n275), .Q(n15[6]));
    nand g88(n192 ,n145 ,n164);
    xnor g89(n345 ,n13[0] ,n14[0]);
    or g90(n413 ,n17[12] ,n1);
    nand g91(n239 ,n392 ,n164);
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n205), .Q(n10[14]));
    not g93(n131 ,n368);
    not g94(n357 ,n382);
    xnor g95(n437 ,n17[11] ,n17[15]);
    buf g96(n3[3], n3[7]);
    not g97(n128 ,n363);
    or g98(n18 ,n15[1] ,n15[0]);
    nand g99(n56 ,n50 ,n52);
    nor g100(n420 ,n405 ,n1);
    nor g101(n211 ,n132 ,n162);
    not g102(n151 ,n6[3]);
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n340), .Q(n4[8]));
    or g104(n411 ,n17[9] ,n1);
    nand g105(n248 ,n15[9] ,n163);
    xor g106(n430 ,n2[1] ,n17[1]);
    nand g107(n102 ,n10[5] ,n100);
    nor g108(n197 ,n8[2] ,n166);
    buf g109(n3[41], n3[47]);
    nand g110(n180 ,n9[2] ,n9[3]);
    nand g111(n382 ,n21 ,n32);
    nor g112(n425 ,n401 ,n1);
    buf g113(n3[8], n3[15]);
    nand g114(n290 ,n9[0] ,n288);
    nand g115(n162 ,n1 ,n2[0]);
    nor g116(n87 ,n15[13] ,n86);
    nand g117(n55 ,n49 ,n51);
    nor g118(n374 ,n115 ,n117);
    nand g119(n185 ,n2[2] ,n2[1]);
    nand g120(n338 ,n331 ,n321);
    xnor g121(n386 ,n15[12] ,n85);
    nand g122(n293 ,n9[3] ,n288);
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n316), .Q(n8[2]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n341), .Q(n4[24]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n431), .Q(n16[7]));
    or g126(n317 ,n16[55] ,n309);
    not g127(n405 ,n17[14]);
    nand g128(n360 ,n377 ,n355);
    buf g129(n3[58], n3[63]);
    nand g130(n265 ,n222 ,n231);
    nand g131(n28 ,n15[6] ,n27);
    nor g132(n73 ,n15[5] ,n72);
    nand g133(n299 ,n256 ,n291);
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n252), .Q(n13[0]));
    nand g135(n99 ,n10[3] ,n98);
    nand g136(n67 ,n15[1] ,n15[0]);
    nand g137(n200 ,n15[0] ,n163);
    nor g138(n301 ,n8[2] ,n289);
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n416), .Q(n17[15]));
    nor g140(n23 ,n15[11] ,n15[10]);
    not g141(n92 ,n10[8]);
    xnor g142(n354 ,n351 ,n350);
    nor g143(n294 ,n148 ,n279);
    nor g144(n173 ,n150 ,n123);
    nor g145(n282 ,n157 ,n254);
    nor g146(n273 ,n123 ,n201);
    nand g147(n120 ,n9[1] ,n9[0]);
    not g148(n226 ,n225);
    nor g149(n342 ,n226 ,n337);
    nor g150(n355 ,n344 ,n353);
    nor g151(n154 ,n141 ,n123);
    not g152(n170 ,n169);
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n412), .Q(n17[7]));
    or g154(n344 ,n7[2] ,n6[4]);
    nand g155(n106 ,n10[7] ,n105);
    nor g156(n289 ,n281 ,n259);
    nand g157(n39 ,n10[8] ,n10[5]);
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n430), .Q(n16[15]));
    xnor g159(n368 ,n10[7] ,n104);
    not g160(n147 ,n6[5]);
    xor g161(n429 ,n2[2] ,n17[2]);
    not g162(n103 ,n102);
    nand g163(n230 ,n185 ,n167);
    nand g164(n236 ,n389 ,n164);
    buf g165(n3[0], n3[7]);
    not g166(n148 ,n11[1]);
    nor g167(n176 ,n152 ,n123);
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n267), .Q(n15[13]));
    nor g169(n343 ,n332 ,n342);
    nand g170(n259 ,n194 ,n230);
    not g171(n121 ,n120);
    nand g172(n361 ,n6[3] ,n7[1]);
    xnor g173(n363 ,n10[2] ,n95);
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n161), .Q(n7[0]));
    nor g175(n352 ,n7[0] ,n349);
    buf g176(n3[27], n3[31]);
    not g177(n48 ,n15[3]);
    not g178(n403 ,n17[11]);
    nor g179(n308 ,n169 ,n306);
    nor g180(n422 ,n406 ,n1);
    nor g181(n252 ,n123 ,n224);
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n206), .Q(n10[13]));
    nand g183(n381 ,n36 ,n47);
    nand g184(n258 ,n200 ,n192);
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n265), .Q(n15[15]));
    not g186(n132 ,n369);
    not g187(n29 ,n28);
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n414), .Q(n17[16]));
    not g189(n75 ,n74);
    not g190(n84 ,n83);
    buf g191(n3[53], n3[55]);
    not g192(n130 ,n371);
    xnor g193(n373 ,n10[12] ,n113);
    nand g194(n296 ,n9[2] ,n288);
    nand g195(n213 ,n15[5] ,n163);
    or g196(n417 ,n17[1] ,n1);
    nor g197(n397 ,n68 ,n66);
    nand g198(n88 ,n15[13] ,n86);
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n292), .Q(n11[2]));
    xnor g200(n375 ,n10[14] ,n116);
    nand g201(n313 ,n8[0] ,n307);
    or g202(n414 ,n17[17] ,n1);
    nand g203(n97 ,n10[2] ,n96);
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n421), .Q(n17[9]));
    buf g205(n3[49], n3[55]);
    xnor g206(n390 ,n15[8] ,n78);
    buf g207(n3[45], n3[47]);
    nand g208(n284 ,n379 ,n273);
    xnor g209(n3[23] ,n356 ,n4[16]);
    or g210(n22 ,n15[13] ,n15[12]);
    nand g211(n183 ,n7[0] ,n7[2]);
    xnor g212(n392 ,n15[6] ,n74);
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n212), .Q(n10[7]));
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n203), .Q(n10[15]));
    buf g215(n3[17], n3[23]);
    xor g216(n428 ,n2[3] ,n17[3]);
    nand g217(n309 ,n1 ,n306);
    nand g218(n266 ,n219 ,n232);
    nor g219(n35 ,n10[11] ,n10[10]);
    nand g220(n232 ,n384 ,n164);
    xnor g221(n369 ,n10[8] ,n106);
    nor g222(n101 ,n10[5] ,n100);
    not g223(n398 ,n355);
    nand g224(n85 ,n15[11] ,n84);
    nor g225(n316 ,n301 ,n311);
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n424), .Q(n17[1]));
    buf g227(n3[35], n3[39]);
    nand g228(n222 ,n15[15] ,n163);
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n210), .Q(n10[10]));
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n432), .Q(n16[39]));
    nor g231(n380 ,n121 ,n119);
    or g232(n315 ,n16[15] ,n309);
    buf g233(n3[60], n3[63]);
    xor g234(n435 ,n2[6] ,n17[6]);
    nand g235(n83 ,n15[10] ,n82);
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n278), .Q(n15[8]));
    nor g237(n50 ,n15[13] ,n15[12]);
    xnor g238(n224 ,n13[0] ,n16[7]);
    xnor g239(n396 ,n15[2] ,n67);
    nor g240(n167 ,n140 ,n8[1]);
    not g241(n137 ,n376);
    buf g242(n3[59], n3[63]);
    xnor g243(n347 ,n9[0] ,n10[0]);
    nand g244(n262 ,n198 ,n228);
    nand g245(n201 ,n8[2] ,n166);
    nand g246(n249 ,n15[10] ,n163);
    nor g247(n80 ,n15[9] ,n79);
    nand g248(n169 ,n1 ,n16[7]);
    not g249(n64 ,n15[8]);
    not g250(n77 ,n76);
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n221), .Q(n10[3]));
    not g252(n402 ,n17[15]);
    nor g253(n203 ,n137 ,n162);
    xnor g254(n3[63] ,n356 ,n4[56]);
    nor g255(n86 ,n65 ,n85);
    buf g256(n3[2], n3[7]);
    nand g257(n267 ,n202 ,n234);
    nor g258(n281 ,n188 ,n257);
    not g259(n149 ,n6[6]);
    not g260(n188 ,n181);
    nor g261(n421 ,n407 ,n1);
    nand g262(n229 ,n397 ,n164);
    not g263(n93 ,n10[12]);
    dff g264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n218), .Q(n10[1]));
    buf g265(n3[20], n3[23]);
    nor g266(n94 ,n10[1] ,n10[0]);
    dff g267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n174), .Q(n6[4]));
    nor g268(n157 ,n144 ,n7[0]);
    nand g269(n254 ,n148 ,n242);
    xnor g270(n359 ,n5[0] ,n360);
    xnor g271(n394 ,n15[4] ,n71);
    nand g272(n109 ,n10[9] ,n107);
    buf g273(n3[32], n3[39]);
    nor g274(n191 ,n165 ,n185);
    nand g275(n233 ,n387 ,n164);
    nand g276(n41 ,n34 ,n35);
    buf g277(n3[4], n3[7]);
    dff g278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n277), .Q(n15[4]));
    not g279(n187 ,n179);
    buf g280(n3[56], n3[63]);
    nand g281(n270 ,n249 ,n250);
    buf g282(n3[30], n3[31]);
    nor g283(n393 ,n73 ,n75);
    xnor g284(n346 ,n11[0] ,n12[0]);
    nor g285(n214 ,n134 ,n162);
    nand g286(n193 ,n187 ,n167);
    nor g287(n424 ,n400 ,n1);
    nand g288(n268 ,n196 ,n235);
    dff g289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n429), .Q(n16[23]));
    xnor g290(n372 ,n10[11] ,n111);
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n270), .Q(n15[10]));
    nand g292(n330 ,n16[31] ,n310);
    dff g293(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n261), .Q(n15[3]));
    nand g294(n260 ,n248 ,n236);
    dff g295(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n190), .Q(n10[0]));
    buf g296(n3[44], n3[47]);
    nor g297(n205 ,n133 ,n162);
    nand g298(n241 ,n394 ,n164);
    or g299(n189 ,n8[0] ,n155);
    not g300(n134 ,n367);
    dff g301(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n433), .Q(n16[63]));
    not g302(n186 ,n171);
    or g303(n45 ,n39 ,n44);
    nand g304(n261 ,n204 ,n227);
    buf g305(n3[50], n3[55]);
    nor g306(n332 ,n8[1] ,n314);
    nand g307(n113 ,n10[11] ,n112);
    nand g308(n199 ,n15[1] ,n163);
    dff g309(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n339), .Q(n4[32]));
    nor g310(n175 ,n146 ,n123);
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n258), .Q(n15[0]));
    nand g312(n30 ,n15[5] ,n29);
    nor g313(n218 ,n139 ,n162);
    nor g314(n423 ,n403 ,n1);
    dff g315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n177), .Q(n7[1]));
    buf g316(n3[43], n3[47]);
    nor g317(n20 ,n15[4] ,n15[3]);
    dff g318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n333), .Q(n4[0]));
    nor g319(n46 ,n38 ,n45);
    nor g320(n389 ,n80 ,n82);
    nand g321(n179 ,n9[0] ,n9[1]);
    nand g322(n204 ,n15[3] ,n163);
    not g323(n136 ,n372);
    not g324(n125 ,n374);
    nand g325(n171 ,n10[0] ,n11[0]);
    buf g326(n3[5], n3[7]);
    not g327(n110 ,n109);
    dff g328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n211), .Q(n10[8]));
    nand g329(n276 ,n213 ,n240);
    nand g330(n228 ,n396 ,n164);
    nor g331(n348 ,n6[6] ,n361);
    xor g332(n436 ,n17[7] ,n17[0]);
    dff g333(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n172), .Q(n6[6]));
    nand g334(n95 ,n10[1] ,n10[0]);
    nor g335(n212 ,n131 ,n162);
    nand g336(n69 ,n15[2] ,n68);
    not g337(n89 ,n88);
    dff g338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n182), .Q(n5[0]));
    nand g339(n353 ,n6[5] ,n352);
    nor g340(n427 ,n402 ,n1);
    buf g341(n3[37], n3[39]);
    not g342(n98 ,n97);
    nand g343(n111 ,n10[10] ,n110);
    nand g344(n240 ,n393 ,n164);
    not g345(n406 ,n17[3]);
    buf g346(n3[21], n3[23]);
    nor g347(n215 ,n126 ,n162);
    nor g348(n100 ,n91 ,n99);
    nand g349(n377 ,n59 ,n62);
    not g350(n139 ,n362);
    nor g351(n177 ,n143 ,n123);
    nand g352(n104 ,n10[6] ,n103);
    nor g353(n79 ,n64 ,n78);
    dff g354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n334), .Q(n4[40]));
    nor g355(n311 ,n292 ,n305);
    dff g356(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n176), .Q(n7[2]));
    nor g357(n164 ,n123 ,n398);
    nor g358(n322 ,n16[7] ,n309);
    nand g359(n27 ,n20 ,n25);
    nand g360(n264 ,n2[0] ,n191);
    dff g361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n207), .Q(n10[12]));
    or g362(n318 ,n16[47] ,n309);
    dff g363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n413), .Q(n17[11]));
    dff g364(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n435), .Q(n16[55]));
    not g365(n123 ,n1);
    xnor g366(n384 ,n15[14] ,n88);
    nor g367(n418 ,n399 ,n1);
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n441), .Q(n17[19]));
    buf g369(n3[52], n3[55]);
    nand g370(n219 ,n15[14] ,n163);
    not g371(n401 ,n17[6]);
    not g372(n140 ,n8[0]);
    xnor g373(n3[47] ,n356 ,n4[40]);
    nand g374(n238 ,n391 ,n164);
    nor g375(n62 ,n15[14] ,n61);
    dff g376(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n343), .Q(n8[1]));
    nor g377(n305 ,n123 ,n299);
    not g378(n126 ,n366);
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n216), .Q(n10[4]));
    dff g380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n274), .Q(n15[7]));
    xnor g381(n365 ,n10[4] ,n99);
    nor g382(n182 ,n123 ,n358);
    nand g383(n24 ,n19 ,n23);
    nand g384(n234 ,n385 ,n164);
    not g385(n141 ,n11[0]);
    not g386(n300 ,n299);
    not g387(n33 ,n10[3]);
    buf g388(n3[34], n3[39]);
    buf g389(n3[29], n3[31]);
    nor g390(n217 ,n128 ,n162);
    xor g391(n433 ,n2[7] ,n17[7]);
    buf g392(n3[28], n3[31]);
    not g393(n124 ,n398);
    not g394(n161 ,n162);
    buf g395(n3[24], n3[31]);
    xnor g396(n3[31] ,n356 ,n4[24]);
    buf g397(n3[25], n3[31]);
    dff g398(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n153), .Q(n11[0]));
    nand g399(n278 ,n247 ,n237);
    buf g400(n3[61], n3[63]);
    dff g401(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n422), .Q(n17[2]));
    nor g402(n59 ,n15[15] ,n56);
    buf g403(n3[40], n3[47]);
    not g404(n287 ,n288);
    dff g405(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n208), .Q(n10[9]));
    nor g406(n32 ,n15[7] ,n31);
    not g407(n105 ,n104);
    xnor g408(n383 ,n90 ,n15[15]);
    nor g409(n174 ,n151 ,n123);
    not g410(n70 ,n69);
    nor g411(n114 ,n93 ,n113);
    not g412(n112 ,n111);
    buf g413(n3[54], n3[55]);
    dff g414(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n418), .Q(n17[6]));
    nor g415(n210 ,n130 ,n162);
    xnor g416(n395 ,n15[3] ,n69);
    nand g417(n257 ,n8[1] ,n195);
    not g418(n358 ,n359);
    dff g419(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n175), .Q(n6[3]));
    dff g420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n423), .Q(n17[10]));
    dff g421(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n184), .Q(n6[7]));
    dff g422(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n268), .Q(n15[12]));
    or g423(n333 ,n308 ,n322);
    nor g424(n163 ,n123 ,n124);
    nor g425(n26 ,n22 ,n24);
    nand g426(n44 ,n10[9] ,n43);
    nand g427(n286 ,n8[2] ,n264);
    nand g428(n341 ,n330 ,n320);
    nand g429(n340 ,n324 ,n315);
    nand g430(n78 ,n15[7] ,n77);
    xnor g431(n3[7] ,n356 ,n4[0]);
    nand g432(n245 ,n15[6] ,n163);
    nor g433(n312 ,n8[0] ,n307);
    buf g434(n3[18], n3[23]);
    not g435(n152 ,n7[1]);
    nor g436(n119 ,n9[1] ,n9[0]);
    dff g437(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n337), .Q(n8[0]));
    buf g438(n3[16], n3[23]);
    nor g439(n419 ,n404 ,n1);
    nand g440(n90 ,n15[14] ,n89);
    nand g441(n326 ,n16[63] ,n310);
    nand g442(n339 ,n329 ,n319);
    dff g443(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n260), .Q(n15[9]));
    nand g444(n194 ,n357 ,n168);
    nand g445(n231 ,n383 ,n164);
    buf g446(n3[57], n3[63]);
    nand g447(n196 ,n15[12] ,n163);
    dff g448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n302), .Q(n9[3]));
    xnor g449(n379 ,n9[2] ,n120);
    or g450(n37 ,n10[2] ,n10[0]);
    nand g451(n220 ,n15[4] ,n163);
    xnor g452(n364 ,n10[3] ,n97);
    nand g453(n328 ,n16[47] ,n310);
    nand g454(n335 ,n327 ,n317);
    nor g455(n216 ,n138 ,n162);
    nor g456(n160 ,n141 ,n9[0]);
    nor g457(n209 ,n136 ,n162);
    nor g458(n51 ,n15[7] ,n15[6]);
    not g459(n91 ,n10[4]);
    nor g460(n307 ,n301 ,n300);
    not g461(n63 ,n15[4]);
    nor g462(n440 ,n1 ,n439);
    buf g463(n3[42], n3[47]);
    or g464(n410 ,n17[4] ,n1);
    xnor g465(n376 ,n118 ,n10[15]);
    not g466(n142 ,n8[1]);
    dff g467(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n273), .Q(n11[3]));
    nand g468(n122 ,n9[2] ,n121);
    buf g469(n3[48], n3[55]);
    nand g470(n274 ,n243 ,n238);
    nand g471(n269 ,n223 ,n233);
    dff g472(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n415), .Q(n17[4]));
    not g473(n143 ,n7[0]);
    nand g474(n334 ,n328 ,n318);
    xor g475(n432 ,n2[4] ,n17[4]);
    or g476(n409 ,n17[13] ,n1);
    nand g477(n165 ,n8[0] ,n8[1]);
    nor g478(n156 ,n11[0] ,n360);
    or g479(n320 ,n16[31] ,n309);
    nand g480(n331 ,n16[23] ,n310);
    nor g481(n207 ,n127 ,n162);
    nor g482(n168 ,n8[0] ,n8[1]);
    xnor g483(n371 ,n10[10] ,n109);
    dff g484(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n410), .Q(n17[3]));
    nor g485(n255 ,n398 ,n189);
    not g486(n96 ,n95);
    nand g487(n247 ,n15[8] ,n163);
    nand g488(n329 ,n16[39] ,n310);
    nand g489(n263 ,n199 ,n229);
    nand g490(n277 ,n220 ,n241);
    not g491(n127 ,n373);
    nand g492(n25 ,n15[2] ,n18);
    nand g493(n246 ,n11[2] ,n158);
    dff g494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n427), .Q(n17[14]));
    not g495(n138 ,n365);
    buf g496(n3[11], n3[15]);
    dff g497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n214), .Q(n10[6]));
    nand g498(n298 ,n280 ,n290);
    nor g499(n385 ,n87 ,n89);
    nor g500(n292 ,n197 ,n287);
    nand g501(n74 ,n15[5] ,n72);
    nand g502(n304 ,n284 ,n296);
    not g503(n133 ,n375);
    buf g504(n3[22], n3[23]);
    xnor g505(n351 ,n346 ,n345);
    not g506(n399 ,n17[7]);
    nand g507(n71 ,n15[3] ,n70);
    xnor g508(n3[55] ,n356 ,n4[48]);
    dff g509(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n251), .Q(n11[1]));
    nand g510(n223 ,n15[11] ,n163);
    nand g511(n38 ,n10[7] ,n10[6]);
    nand g512(n438 ,n436 ,n437);
    buf g513(n3[13], n3[15]);
    buf g514(n3[33], n3[39]);
    xnor g515(n367 ,n10[6] ,n102);
    dff g516(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n262), .Q(n15[2]));
    dff g517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n173), .Q(n6[5]));
    nor g518(n58 ,n15[2] ,n57);
    buf g519(n3[36], n3[39]);
    not g520(n166 ,n165);
    nor g521(n108 ,n10[9] ,n107);
    nor g522(n253 ,n160 ,n246);
    xnor g523(n3[39] ,n356 ,n4[32]);
    nand g524(n302 ,n283 ,n293);
    dff g525(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n420), .Q(n17[13]));
    or g526(n61 ,n55 ,n60);
    nor g527(n72 ,n63 ,n71);
    dff g528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n170), .Q(n12[0]));
    nand g529(n235 ,n386 ,n164);
    not g530(n146 ,n7[2]);
    or g531(n319 ,n16[39] ,n309);
    nand g532(n243 ,n15[7] ,n163);
    nor g533(n297 ,n282 ,n294);
    nand g534(n275 ,n245 ,n239);
    nand g535(n116 ,n10[13] ,n114);
    nor g536(n244 ,n186 ,n156);
    dff g537(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n428), .Q(n16[31]));
    nor g538(n60 ,n54 ,n58);
    nand g539(n31 ,n26 ,n30);
    or g540(n158 ,n11[0] ,n8[0]);
    nand g541(n303 ,n285 ,n295);
    nand g542(n325 ,n1 ,n313);
    dff g543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n336), .Q(n4[56]));
    nand g544(n198 ,n15[2] ,n163);
    xnor g545(n378 ,n9[3] ,n122);
    not g546(n272 ,n273);
    dff g547(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n425), .Q(n17[5]));
    nor g548(n291 ,n255 ,n286);
    nor g549(n21 ,n15[9] ,n15[8]);
    not g550(n68 ,n67);
    nand g551(n81 ,n15[9] ,n79);
    nor g552(n279 ,n271 ,n253);
    nor g553(n288 ,n123 ,n273);
    dff g554(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n154), .Q(n14[0]));
    nor g555(n362 ,n96 ,n94);
    dff g556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n298), .Q(n9[0]));
    nand g557(n202 ,n15[13] ,n163);
    xnor g558(n3[15] ,n356 ,n4[8]);
    dff g559(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n276), .Q(n15[5]));
    nor g560(n49 ,n15[9] ,n15[8]);
    nor g561(n366 ,n101 ,n103);
    or g562(n323 ,n16[63] ,n309);
    dff g563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n426), .Q(n17[18]));
    dff g564(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n269), .Q(n15[11]));
    nand g565(n250 ,n388 ,n164);
    nor g566(n153 ,n123 ,n8[0]);
    buf g567(n3[9], n3[15]);
    not g568(n135 ,n364);
    nand g569(n227 ,n395 ,n164);
    nand g570(n349 ,n6[7] ,n348);
    nor g571(n172 ,n147 ,n123);
    nand g572(n178 ,n11[0] ,n2[0]);
    xnor g573(n387 ,n15[11] ,n83);
    nand g574(n118 ,n10[14] ,n117);
    nor g575(n271 ,n11[2] ,n244);
    dff g576(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n409), .Q(n17[12]));
    not g577(n150 ,n6[4]);
    nor g578(n370 ,n108 ,n110);
endmodule
