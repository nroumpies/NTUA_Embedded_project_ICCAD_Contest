module top (n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n11);
    input [63:0] n0;
    input [31:0] n1;
    input [3:0] n2;
    input n3;
    input [1:0] n4;
    input [5:0] n5;
    output [63:0] n6;
    output [31:0] n7;
    output n8, n9, n10, n11;
    output [5:0] n12;
    output [7:0] n13;
    wire [63:0] n0;
    wire [31:0] n1;
    wire [3:0] n2;
    wire n3;
    wire [1:0] n4;
    wire [5:0] n5;
    wire [63:0] n6;
    wire [31:0] n7;
    wire n8, n9, n10, n11;
    wire [5:0] n12;
    wire [7:0] n13;
    wire n14, n15, n16, n17, n18, n19, n20, n21;
    wire n22, n23, n24, n25, n26, n27, n28, n29;
    wire n30, n31, n32, n33, n34, n35, n36, n37;
    wire n38, n39, n40, n41, n42, n43, n44, n45;
    wire n46, n47, n48, n49, n50, n51, n52, n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171, n172, n173;
    wire n174, n175, n176, n177, n178, n179, n180, n181;
    wire n182, n183, n184, n185, n186, n187, n188, n189;
    wire n190, n191, n192, n193, n194, n195, n196, n197;
    wire n198, n199, n200, n201, n202, n203, n204, n205;
    wire n206, n207, n208, n209, n210, n211, n212, n213;
    wire n214, n215, n216, n217, n218, n219, n220, n221;
    wire n222, n223, n224, n225, n226, n227, n228, n229;
    wire n230, n231, n232, n233, n234, n235, n236, n237;
    wire n238, n239, n240, n241, n242, n243, n244, n245;
    wire n246, n247, n248, n249, n250, n251, n252, n253;
    wire n254, n255, n256, n257, n258, n259, n260, n261;
    wire n262, n263, n264, n265, n266, n267, n268, n269;
    wire n270, n271, n272, n273, n274, n275, n276, n277;
    wire n278, n279, n280, n281, n282, n283, n284, n285;
    wire n286, n287, n288, n289, n290, n291, n292, n293;
    wire n294, n295, n296, n297, n298, n299, n300, n301;
    wire n302, n303, n304, n305, n306, n307, n308, n309;
    wire n310, n311, n312, n313, n314, n315, n316, n317;
    wire n318, n319, n320, n321, n322, n323, n324, n325;
    wire n326, n327, n328, n329, n330, n331, n332, n333;
    wire n334, n335, n336, n337, n338, n339, n340, n341;
    wire n342, n343, n344, n345, n346, n347, n348, n349;
    wire n350, n351, n352, n353, n354, n355, n356, n357;
    wire n358, n359, n360, n361, n362, n363, n364, n365;
    wire n366, n367, n368, n369, n370, n371, n372, n373;
    wire n374, n375, n376, n377, n378, n379, n380, n381;
    wire n382, n383, n384, n385, n386, n387, n388, n389;
    wire n390, n391, n392, n393, n394, n395, n396, n397;
    wire n398, n399, n400, n401, n402, n403, n404, n405;
    wire n406, n407, n408, n409, n410, n411, n412, n413;
    wire n414, n415, n416, n417, n418, n419, n420, n421;
    wire n422, n423, n424, n425, n426, n427, n428, n429;
    wire n430, n431, n432, n433, n434, n435, n436, n437;
    wire n438, n439, n440, n441, n442, n443, n444, n445;
    wire n446, n447, n448, n449, n450, n451, n452, n453;
    wire n454, n455, n456, n457, n458, n459, n460, n461;
    wire n462, n463, n464, n465, n466, n467, n468, n469;
    wire n470, n471, n472, n473, n474, n475, n476, n477;
    wire n478, n479, n480, n481, n482, n483, n484, n485;
    wire n486, n487, n488, n489, n490, n491, n492, n493;
    wire n494, n495, n496, n497, n498, n499, n500, n501;
    wire n502, n503, n504, n505, n506, n507, n508, n509;
    wire n510, n511, n512, n513, n514, n515, n516, n517;
    wire n518, n519, n520, n521, n522, n523, n524, n525;
    wire n526, n527, n528, n529, n530, n531, n532, n533;
    wire n534, n535, n536, n537, n538, n539, n540, n541;
    wire n542, n543, n544, n545, n546, n547, n548, n549;
    wire n550, n551, n552, n553, n554, n555, n556, n557;
    wire n558, n559, n560, n561, n562, n563, n564, n565;
    wire n566, n567, n568, n569, n570, n571, n572, n573;
    wire n574, n575, n576, n577, n578, n579, n580, n581;
    wire n582, n583, n584, n585, n586, n587, n588, n589;
    wire n590, n591, n592, n593, n594, n595, n596, n597;
    wire n598, n599, n600, n601, n602, n603, n604, n605;
    wire n606, n607, n608, n609, n610, n611, n612, n613;
    wire n614, n615, n616, n617, n618, n619, n620, n621;
    wire n622, n623, n624, n625, n626, n627, n628, n629;
    wire n630, n631, n632, n633, n634, n635, n636, n637;
    wire n638, n639, n640, n641, n642, n643, n644, n645;
    wire n646, n647, n648, n649, n650, n651, n652, n653;
    wire n654, n655, n656, n657, n658, n659, n660, n661;
    wire n662, n663, n664, n665, n666, n667, n668, n669;
    wire n670, n671, n672, n673, n674, n675, n676, n677;
    wire n678, n679, n680, n681, n682, n683, n684, n685;
    wire n686, n687, n688, n689, n690, n691, n692, n693;
    wire n694, n695, n696, n697, n698, n699, n700, n701;
    wire n702, n703, n704, n705, n706, n707, n708, n709;
    wire n710, n711, n712, n713, n714, n715, n716, n717;
    wire n718, n719, n720, n721, n722, n723, n724, n725;
    wire n726, n727, n728, n729, n730, n731, n732, n733;
    wire n734, n735, n736, n737, n738, n739, n740, n741;
    wire n742, n743, n744, n745, n746, n747, n748, n749;
    wire n750, n751, n752, n753, n754, n755, n756, n757;
    wire n758, n759, n760, n761, n762, n763, n764, n765;
    wire n766, n767, n768, n769, n770, n771, n772, n773;
    wire n774, n775, n776, n777, n778, n779, n780, n781;
    wire n782, n783, n784, n785, n786, n787, n788, n789;
    wire n790, n791, n792, n793, n794, n795, n796, n797;
    wire n798, n799, n800, n801, n802, n803, n804, n805;
    wire n806, n807, n808, n809, n810, n811, n812, n813;
    wire n814, n815, n816, n817, n818, n819, n820, n821;
    wire n822, n823, n824, n825, n826, n827, n828, n829;
    wire n830, n831, n832, n833, n834, n835, n836, n837;
    wire n838, n839, n840, n841, n842, n843, n844, n845;
    wire n846, n847, n848, n849, n850, n851, n852, n853;
    wire n854, n855, n856, n857, n858, n859, n860, n861;
    wire n862, n863, n864, n865, n866, n867, n868, n869;
    wire n870, n871, n872, n873, n874, n875, n876, n877;
    wire n878, n879, n880, n881, n882, n883, n884, n885;
    wire n886, n887, n888, n889, n890, n891, n892, n893;
    wire n894, n895, n896, n897, n898, n899, n900, n901;
    wire n902, n903, n904, n905, n906, n907, n908, n909;
    wire n910, n911, n912, n913, n914, n915, n916, n917;
    wire n918, n919, n920, n921, n922, n923, n924, n925;
    wire n926, n927, n928, n929, n930, n931, n932, n933;
    wire n934, n935, n936, n937, n938, n939, n940, n941;
    wire n942, n943, n944, n945, n946, n947, n948, n949;
    wire n950, n951, n952, n953, n954, n955, n956, n957;
    wire n958, n959, n960, n961, n962, n963, n964, n965;
    wire n966, n967, n968, n969, n970, n971, n972, n973;
    wire n974, n975, n976, n977, n978, n979, n980, n981;
    wire n982, n983, n984, n985, n986, n987, n988, n989;
    wire n990, n991, n992, n993, n994, n995, n996, n997;
    wire n998, n999, n1000, n1001, n1002, n1003, n1004, n1005;
    wire n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013;
    wire n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
    wire n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
    wire n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
    wire n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;
    wire n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053;
    wire n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061;
    wire n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069;
    wire n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077;
    wire n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085;
    wire n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093;
    wire n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101;
    wire n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109;
    wire n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117;
    wire n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125;
    wire n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133;
    wire n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141;
    wire n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149;
    wire n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157;
    wire n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165;
    wire n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173;
    wire n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181;
    wire n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189;
    wire n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197;
    wire n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205;
    wire n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
    wire n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221;
    wire n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229;
    wire n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237;
    wire n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245;
    wire n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253;
    wire n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261;
    wire n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269;
    wire n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277;
    wire n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285;
    wire n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293;
    wire n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301;
    wire n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309;
    wire n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;
    wire n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325;
    wire n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333;
    wire n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;
    wire n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349;
    wire n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;
    wire n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365;
    wire n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373;
    wire n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381;
    wire n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389;
    wire n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397;
    wire n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405;
    wire n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413;
    wire n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421;
    wire n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429;
    wire n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437;
    wire n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445;
    wire n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453;
    wire n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461;
    wire n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469;
    wire n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477;
    wire n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485;
    wire n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493;
    wire n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501;
    wire n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509;
    wire n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517;
    wire n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525;
    wire n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533;
    wire n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541;
    wire n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
    wire n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557;
    wire n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565;
    wire n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573;
    wire n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581;
    wire n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589;
    wire n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597;
    wire n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605;
    wire n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613;
    wire n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621;
    wire n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629;
    wire n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637;
    wire n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645;
    wire n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653;
    wire n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661;
    wire n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669;
    wire n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677;
    wire n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685;
    wire n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693;
    wire n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701;
    wire n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709;
    wire n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717;
    wire n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725;
    wire n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733;
    wire n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741;
    wire n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749;
    wire n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757;
    wire n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765;
    wire n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773;
    wire n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781;
    wire n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789;
    wire n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797;
    wire n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805;
    wire n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813;
    wire n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821;
    wire n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829;
    wire n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837;
    wire n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845;
    wire n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853;
    wire n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861;
    wire n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869;
    wire n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877;
    wire n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885;
    wire n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893;
    wire n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901;
    wire n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909;
    wire n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917;
    wire n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925;
    wire n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933;
    wire n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941;
    wire n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949;
    wire n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957;
    wire n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965;
    wire n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973;
    wire n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981;
    wire n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989;
    wire n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997;
    wire n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005;
    wire n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013;
    wire n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021;
    wire n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029;
    wire n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037;
    wire n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045;
    wire n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053;
    wire n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061;
    wire n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069;
    wire n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077;
    wire n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085;
    wire n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093;
    wire n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101;
    wire n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109;
    wire n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117;
    wire n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125;
    wire n2126;
    nand g0(n1527 ,n1[16] ,n1235);
    nand g1(n86 ,n0[19] ,n0[3]);
    nand g2(n652 ,n611 ,n638);
    nand g3(n1864 ,n1826 ,n1848);
    xnor g4(n6[49] ,n0[49] ,n1282);
    xnor g5(n428 ,n2068 ,n2063);
    nand g6(n1800 ,n1682 ,n1708);
    or g7(n58 ,n0[27] ,n0[11]);
    nor g8(n777 ,n738 ,n1[6]);
    nand g9(n1659 ,n1522 ,n1423);
    xnor g10(n871 ,n0[59] ,n0[35]);
    nand g11(n448 ,n2062 ,n384);
    xnor g12(n201 ,n96 ,n155);
    nand g13(n77 ,n0[59] ,n0[43]);
    xnor g14(n679 ,n657 ,n640);
    nor g15(n1815 ,n1536 ,n1754);
    nor g16(n1615 ,n1450 ,n1496);
    nor g17(n1347 ,n752 ,n1099);
    or g18(n237 ,n214 ,n201);
    nor g19(n1428 ,n1198 ,n1149);
    nand g20(n1289 ,n2023 ,n1107);
    nand g21(n414 ,n2086 ,n2050);
    nand g22(n328 ,n294 ,n316);
    xnor g23(n1244 ,n0[52] ,n930);
    xnor g24(n44 ,n1973 ,n1975);
    or g25(n2112 ,n5[2] ,n2105);
    nor g26(n1035 ,n1[5] ,n981);
    xor g27(n1226 ,n0[62] ,n909);
    nand g28(n1964 ,n2030 ,n1959);
    xnor g29(n869 ,n0[35] ,n0[34]);
    xnor g30(n109 ,n0[20] ,n0[4]);
    xnor g31(n279 ,n257 ,n250);
    not g32(n2034 ,n0[63]);
    or g33(n395 ,n2041 ,n2044);
    xnor g34(n850 ,n0[39] ,n0[23]);
    or g35(n61 ,n0[59] ,n0[43]);
    nand g36(n1078 ,n0[2] ,n998);
    nand g37(n87 ,n0[61] ,n0[45]);
    nand g38(n990 ,n2[3] ,n807);
    nand g39(n1163 ,n884 ,n1046);
    xnor g40(n696 ,n677 ,n634);
    nand g41(n611 ,n565 ,n582);
    nand g42(n213 ,n79 ,n181);
    not g43(n2094 ,n0[3]);
    nand g44(n1283 ,n2027 ,n1107);
    nand g45(n1642 ,n1[11] ,n1553);
    xnor g46(n922 ,n0[16] ,n0[15]);
    xnor g47(n988 ,n0[8] ,n0[7]);
    nand g48(n1785 ,n1475 ,n1755);
    nand g49(n836 ,n5[3] ,n771);
    nor g50(n1705 ,n1103 ,n1584);
    nand g51(n244 ,n78 ,n211);
    nor g52(n1507 ,n1168 ,n1371);
    nand g53(n75 ,n0[56] ,n0[8]);
    nor g54(n1449 ,n1047 ,n1245);
    nor g55(n1624 ,n1466 ,n1492);
    nand g56(n469 ,n410 ,n450);
    nor g57(n1860 ,n2009 ,n1831);
    or g58(n394 ,n2038 ,n2061);
    xnor g59(n6[58] ,n0[58] ,n1277);
    nor g60(n2022 ,n5[2] ,n2122);
    nand g61(n306 ,n244 ,n285);
    nand g62(n1853 ,n1745 ,n1794);
    nor g63(n2117 ,n2103 ,n2107);
    nor g64(n1605 ,n1511 ,n1519);
    xnor g65(n263 ,n242 ,n230);
    nand g66(n591 ,n541 ,n560);
    xnor g67(n597 ,n521 ,n572);
    nand g68(n235 ,n157 ,n198);
    nor g69(n1450 ,n1047 ,n1251);
    nand g70(n368 ,n357 ,n365);
    xnor g71(n892 ,n0[23] ,n0[22]);
    nand g72(n236 ,n217 ,n177);
    or g73(n618 ,n569 ,n597);
    xnor g74(n221 ,n152 ,n174);
    nand g75(n539 ,n496 ,n492);
    nand g76(n122 ,n0[51] ,n61);
    nand g77(n540 ,n518 ,n519);
    xnor g78(n436 ,n2085 ,n2054);
    xnor g79(n1567 ,n1217 ,n1221);
    xnor g80(n917 ,n0[26] ,n0[25]);
    nor g81(n1813 ,n1760 ,n1710);
    xnor g82(n284 ,n247 ,n258);
    nand g83(n157 ,n83 ,n126);
    not g84(n2052 ,n0[45]);
    or g85(n7[6] ,n1844 ,n1796);
    nand g86(n1397 ,n1994 ,n1106);
    xnor g87(n6[33] ,n0[33] ,n1279);
    nand g88(n481 ,n403 ,n447);
    xnor g89(n6[16] ,n0[16] ,n1320);
    xor g90(n1855 ,n1[9] ,n1791);
    nand g91(n1894 ,n1883 ,n1893);
    xnor g92(n656 ,n633 ,n637);
    nand g93(n584 ,n539 ,n561);
    nand g94(n196 ,n163 ,n162);
    xnor g95(n678 ,n660 ,n661);
    nand g96(n1270 ,n2026 ,n1053);
    nand g97(n826 ,n1999 ,n745);
    not g98(n1101 ,n1102);
    nand g99(n7[21] ,n1666 ,n1615);
    xnor g100(n976 ,n0[1] ,n0[0]);
    nor g101(n1722 ,n1554 ,n1574);
    xnor g102(n494 ,n438 ,n2046);
    nand g103(n455 ,n2058 ,n380);
    nand g104(n1345 ,n0[28] ,n1100);
    nor g105(n1719 ,n1554 ,n1573);
    nor g106(n1851 ,n1787 ,n1786);
    nand g107(n1057 ,n1[3] ,n984);
    nor g108(n1009 ,n1[4] ,n980);
    or g109(n1020 ,n1[26] ,n898);
    nor g110(n1887 ,n1854 ,n1882);
    or g111(n697 ,n676 ,n685);
    xnor g112(n1561 ,n1[11] ,n1247);
    nand g113(n74 ,n0[62] ,n0[46]);
    nand g114(n1645 ,n1[15] ,n1553);
    or g115(n1627 ,n1194 ,n1516);
    nand g116(n637 ,n606 ,n620);
    xnor g117(n28 ,n20 ,n2005);
    nand g118(n1843 ,n1595 ,n1790);
    xnor g119(n429 ,n2072 ,n2051);
    xnor g120(n1992 ,n322 ,n323);
    nand g121(n1756 ,n1518 ,n1662);
    xnor g122(n1119 ,n872 ,n910);
    nand g123(n783 ,n0[59] ,n742);
    or g124(n1753 ,n1629 ,n1542);
    nand g125(n1146 ,n982 ,n1105);
    nand g126(n73 ,n0[42] ,n0[10]);
    nand g127(n817 ,n1992 ,n741);
    nand g128(n514 ,n467 ,n472);
    nor g129(n1416 ,n1136 ,n1367);
    nor g130(n1024 ,n1[2] ,n985);
    nand g131(n184 ,n156 ,n149);
    not g132(n1099 ,n1100);
    nor g133(n1794 ,n1549 ,n1730);
    nand g134(n2118 ,n5[0] ,n2110);
    nand g135(n486 ,n417 ,n462);
    xnor g136(n942 ,n0[31] ,n0[7]);
    or g137(n1041 ,n1[15] ,n988);
    nand g138(n1398 ,n1995 ,n1106);
    or g139(n509 ,n469 ,n483);
    nand g140(n824 ,n1983 ,n758);
    xnor g141(n592 ,n571 ,n569);
    nor g142(n1181 ,n1074 ,n1047);
    nor g143(n1715 ,n1541 ,n1623);
    nor g144(n1690 ,n1[14] ,n1579);
    not g145(n2107 ,n2106);
    or g146(n42 ,n1973 ,n1974);
    xnor g147(n885 ,n0[15] ,n0[14]);
    nand g148(n1064 ,n1[8] ,n890);
    nand g149(n1532 ,n1[22] ,n1242);
    nor g150(n375 ,n369 ,n374);
    xnor g151(n941 ,n0[53] ,n0[5]);
    nor g152(n1698 ,n1659 ,n1661);
    nand g153(n724 ,n714 ,n715);
    nor g154(n1837 ,n2009 ,n2010);
    nor g155(n1694 ,n1368 ,n1600);
    xnor g156(n643 ,n619 ,n581);
    nor g157(n1004 ,n963 ,n954);
    nand g158(n215 ,n91 ,n183);
    nand g159(n291 ,n210 ,n264);
    nand g160(n148 ,n74 ,n123);
    nand g161(n1284 ,n2026 ,n1107);
    xnor g162(n106 ,n0[42] ,n0[10]);
    xnor g163(n897 ,n0[27] ,n752);
    not g164(n760 ,n0[7]);
    not g165(n2077 ,n0[20]);
    nand g166(n963 ,n802 ,n800);
    nand g167(n1143 ,n983 ,n1105);
    nor g168(n1435 ,n1018 ,n1190);
    or g169(n531 ,n491 ,n488);
    xnor g170(n427 ,n2037 ,n2082);
    nor g171(n1073 ,n739 ,n979);
    xnor g172(n1791 ,n1555 ,n902);
    or g173(n7[5] ,n1839 ,n1798);
    nand g174(n624 ,n598 ,n596);
    nand g175(n1373 ,n1022 ,n1096);
    xnor g176(n6[6] ,n0[6] ,n1309);
    nor g177(n1959 ,n1928 ,n1954);
    xnor g178(n6[2] ,n0[2] ,n1305);
    xnor g179(n432 ,n2070 ,n2056);
    nand g180(n541 ,n495 ,n494);
    xnor g181(n1583 ,n0[63] ,n1218);
    nand g182(n447 ,n2074 ,n396);
    nor g183(n971 ,n753 ,n837);
    xnor g184(n103 ,n0[39] ,n0[15]);
    nand g185(n839 ,n2[2] ,n770);
    xnor g186(n1577 ,n0[58] ,n1221);
    xor g187(n1250 ,n0[34] ,n873);
    not g188(n1974 ,n2015);
    nand g189(n452 ,n2077 ,n392);
    nor g190(n1409 ,n1377 ,n1381);
    nor g191(n807 ,n2[2] ,n2[1]);
    nor g192(n616 ,n598 ,n596);
    xnor g193(n161 ,n104 ,n95);
    or g194(n1599 ,n1498 ,n1539);
    nand g195(n571 ,n516 ,n547);
    xnor g196(n931 ,n0[60] ,n0[44]);
    xnor g197(n105 ,n0[56] ,n0[8]);
    nand g198(n349 ,n321 ,n342);
    xnor g199(n430 ,n2041 ,n2097);
    xnor g200(n1122 ,n870 ,n909);
    nand g201(n1643 ,n1[12] ,n1553);
    nor g202(n1431 ,n1379 ,n1370);
    nand g203(n818 ,n1984 ,n756);
    or g204(n324 ,n262 ,n320);
    not g205(n754 ,n0[1]);
    xnor g206(n104 ,n0[19] ,n0[3]);
    nand g207(n329 ,n297 ,n317);
    or g208(n7[30] ,n1343 ,n1765);
    or g209(n1870 ,n1811 ,n1862);
    xnor g210(n1112 ,n867 ,n938);
    nand g211(n458 ,n2034 ,n398);
    nand g212(n1200 ,n0[59] ,n1101);
    nor g213(n1610 ,n1547 ,n1543);
    not g214(n749 ,n0[60]);
    xnor g215(n861 ,n0[53] ,n0[52]);
    xnor g216(n266 ,n218 ,n160);
    not g217(n742 ,n1[3]);
    not g218(n772 ,n5[3]);
    nand g219(n1310 ,n2020 ,n1109);
    nand g220(n378 ,n344 ,n377);
    nand g221(n1797 ,n1465 ,n1724);
    nand g222(n404 ,n2079 ,n2078);
    nand g223(n472 ,n404 ,n460);
    or g224(n1179 ,n914 ,n1045);
    nor g225(n1790 ,n1721 ,n1717);
    nand g226(n1299 ,n2023 ,n1049);
    xnor g227(n113 ,n0[59] ,n0[51]);
    nand g228(n212 ,n176 ,n186);
    nor g229(n804 ,n739 ,n1987);
    nor g230(n369 ,n356 ,n368);
    nand g231(n786 ,n0[58] ,n741);
    xnor g232(n166 ,n106 ,n0[34]);
    nand g233(n1302 ,n2026 ,n1049);
    nand g234(n1097 ,n1[27] ,n915);
    nand g235(n216 ,n138 ,n184);
    nand g236(n1455 ,n1048 ,n1255);
    nand g237(n1060 ,n1[0] ,n976);
    not g238(n1254 ,n1253);
    nand g239(n1296 ,n2020 ,n1107);
    nand g240(n1095 ,n1[31] ,n914);
    xnor g241(n554 ,n504 ,n496);
    nand g242(n1634 ,n1[30] ,n1553);
    nand g243(n516 ,n479 ,n478);
    or g244(n1685 ,n1554 ,n1576);
    nand g245(n18 ,n2010 ,n2007);
    nand g246(n538 ,n491 ,n488);
    nand g247(n1349 ,n0[23] ,n1100);
    nor g248(n1149 ,n980 ,n1045);
    nand g249(n46 ,n43 ,n45);
    not g250(n1552 ,n1553);
    nand g251(n302 ,n266 ,n282);
    xnor g252(n1771 ,n1[8] ,n1566);
    xnor g253(n1995 ,n361 ,n372);
    or g254(n1036 ,n1[31] ,n914);
    nand g255(n1007 ,n756 ,n975);
    nor g256(n357 ,n333 ,n345);
    nand g257(n449 ,n2036 ,n393);
    nor g258(n1182 ,n0[2] ,n1098);
    or g259(n1821 ,n1707 ,n1737);
    nand g260(n1530 ,n1[18] ,n1257);
    nand g261(n713 ,n700 ,n706);
    not g262(n744 ,n0[5]);
    nand g263(n254 ,n233 ,n243);
    not g264(n762 ,n1[12]);
    nand g265(n1495 ,n1352 ,n1154);
    nand g266(n1298 ,n2022 ,n1049);
    nand g267(n1679 ,n1[29] ,n1553);
    nand g268(n1478 ,n1[9] ,n1256);
    nand g269(n1395 ,n1089 ,n1076);
    not g270(n1908 ,n4[1]);
    nand g271(n1949 ,n1936 ,n1934);
    nor g272(n1328 ,n945 ,n1091);
    nand g273(n1863 ,n1825 ,n1824);
    not g274(n761 ,n1[8]);
    nand g275(n1758 ,n1642 ,n1457);
    nand g276(n972 ,n2001 ,n823);
    xnor g277(n907 ,n0[28] ,n0[12]);
    nand g278(n226 ,n173 ,n194);
    not g279(n741 ,n1[2]);
    nor g280(n2120 ,n2108 ,n2115);
    xnor g281(n1114 ,n866 ,n940);
    xnor g282(n1570 ,n0[7] ,n1224);
    or g283(n604 ,n576 ,n578);
    nand g284(n560 ,n503 ,n532);
    nand g285(n1206 ,n1034 ,n1068);
    nand g286(n844 ,n5[4] ,n5[3]);
    nand g287(n142 ,n93 ,n136);
    nand g288(n134 ,n0[52] ,n64);
    xnor g289(n579 ,n524 ,n486);
    nor g290(n1617 ,n1452 ,n1404);
    or g291(n1789 ,n1548 ,n1743);
    xnor g292(n1555 ,n0[41] ,n1223);
    or g293(n632 ,n581 ,n619);
    nand g294(n473 ,n412 ,n454);
    nand g295(n1141 ,n979 ,n1105);
    nand g296(n1865 ,n1652 ,n1828);
    nand g297(n1671 ,n1[18] ,n1553);
    nand g298(n91 ,n0[21] ,n0[5]);
    nand g299(n814 ,n1988 ,n755);
    nand g300(n1903 ,n2018 ,n1898);
    nand g301(n583 ,n568 ,n567);
    or g302(n566 ,n477 ,n537);
    nand g303(n1744 ,n1[7] ,n1570);
    nand g304(n1533 ,n1356 ,n1365);
    nand g305(n257 ,n207 ,n225);
    xor g306(n2018 ,n39 ,n34);
    or g307(n392 ,n2094 ,n2089);
    nand g308(n1850 ,n1814 ,n1715);
    xor g309(n1257 ,n0[58] ,n855);
    nor g310(n1169 ,n915 ,n1045);
    or g311(n1962 ,n1916 ,n1957);
    nand g312(n252 ,n187 ,n231);
    or g313(n658 ,n646 ,n645);
    nor g314(n947 ,n787 ,n784);
    or g315(n989 ,n2[1] ,n839);
    xnor g316(n670 ,n643 ,n648);
    not g317(n735 ,n2012);
    not g318(n751 ,n0[29]);
    xnor g319(n847 ,n0[27] ,n0[11]);
    nand g320(n1160 ,n880 ,n1046);
    nand g321(n1272 ,n2025 ,n1108);
    xnor g322(n6[20] ,n0[20] ,n1300);
    xnor g323(n920 ,n0[30] ,n0[29]);
    xnor g324(n270 ,n223 ,n216);
    not g325(n2095 ,n0[2]);
    nand g326(n130 ,n0[63] ,n67);
    or g327(n1711 ,n1102 ,n1581);
    nand g328(n1070 ,n1[1] ,n976);
    or g329(n401 ,n2091 ,n2037);
    or g330(n1683 ,n1554 ,n1575);
    nand g331(n1490 ,n776 ,n1207);
    xnor g332(n108 ,n0[23] ,n0[7]);
    xnor g333(n598 ,n554 ,n492);
    nor g334(n1682 ,n1589 ,n1612);
    xnor g335(n601 ,n551 ,n503);
    xnor g336(n1775 ,n1[5] ,n1580);
    nand g337(n1730 ,n1632 ,n1428);
    nand g338(n319 ,n278 ,n296);
    nor g339(n951 ,n791 ,n781);
    nand g340(n208 ,n159 ,n160);
    xnor g341(n6[32] ,n0[32] ,n1281);
    nand g342(n1641 ,n1[10] ,n1553);
    nor g343(n1879 ,n1834 ,n1871);
    or g344(n1724 ,n1554 ,n1568);
    nand g345(n1266 ,n2020 ,n1051);
    not g346(n2050 ,n0[47]);
    nor g347(n1418 ,n1182 ,n1132);
    xnor g348(n496 ,n441 ,n2035);
    xnor g349(n223 ,n163 ,n161);
    xor g350(n1910 ,n0[20] ,n1[20]);
    nor g351(n1629 ,n756 ,n1552);
    nand g352(n209 ,n152 ,n167);
    nand g353(n1763 ,n1676 ,n1158);
    nand g354(n722 ,n713 ,n717);
    nand g355(n297 ,n267 ,n284);
    nand g356(n1657 ,n1529 ,n1480);
    nor g357(n1074 ,n0[37] ,n877);
    nor g358(n1422 ,n1[8] ,n1233);
    not g359(n423 ,n422);
    xnor g360(n710 ,n696 ,n682);
    xnor g361(n619 ,n573 ,n520);
    xor g362(n2014 ,n1976 ,n48);
    nor g363(n1886 ,n990 ,n1879);
    nor g364(n1655 ,n1545 ,n1456);
    nand g365(n1068 ,n1[6] ,n978);
    nand g366(n7[20] ,n1665 ,n1614);
    or g367(n138 ,n94 ,n115);
    nor g368(n1889 ,n2004 ,n1884);
    nor g369(n1510 ,n1[20] ,n1228);
    nor g370(n1689 ,n1[11] ,n1585);
    nor g371(n1152 ,n984 ,n1045);
    nor g372(n1822 ,n1102 ,n1791);
    nor g373(n1108 ,n808 ,n994);
    nand g374(n1290 ,n2025 ,n1053);
    nor g375(n1430 ,n1103 ,n1233);
    not g376(n743 ,n1[7]);
    nand g377(n49 ,n1976 ,n48);
    nor g378(n1826 ,n1775 ,n1818);
    xor g379(n1998 ,n351 ,n375);
    nand g380(n407 ,n2070 ,n2057);
    xnor g381(n203 ,n111 ,n147);
    or g382(n617 ,n594 ,n599);
    nor g383(n367 ,n356 ,n364);
    not g384(n1975 ,n2001);
    nand g385(n1390 ,n1991 ,n1106);
    nand g386(n825 ,n1991 ,n756);
    xnor g387(n667 ,n653 ,n647);
    nand g388(n1528 ,n1[23] ,n1248);
    nand g389(n703 ,n676 ,n685);
    nand g390(n1492 ,n1210 ,n1164);
    nor g391(n1697 ,n1103 ,n1586);
    nor g392(n1107 ,n844 ,n995);
    nor g393(n1867 ,n1835 ,n1836);
    nand g394(n718 ,n703 ,n712);
    nand g395(n608 ,n577 ,n584);
    xnor g396(n657 ,n611 ,n638);
    nand g397(n1680 ,n1[31] ,n1553);
    or g398(n533 ,n493 ,n498);
    nand g399(n204 ,n145 ,n178);
    not g400(n753 ,n2016);
    or g401(n1458 ,n1047 ,n1239);
    nand g402(n1278 ,n2022 ,n1108);
    nand g403(n1649 ,n1411 ,n1410);
    xnor g404(n6[31] ,n0[31] ,n1283);
    xnor g405(n705 ,n641 ,n694);
    or g406(n1426 ,n1140 ,n1180);
    or g407(n530 ,n496 ,n492);
    nand g408(n1082 ,n1[18] ,n883);
    or g409(n7[25] ,n1348 ,n1762);
    nand g410(n1804 ,n1734 ,n1691);
    nand g411(n390 ,n2038 ,n2061);
    nand g412(n1376 ,n1998 ,n1106);
    xnor g413(n187 ,n0[0] ,n105);
    nand g414(n1859 ,n1134 ,n1847);
    xnor g415(n2011 ,n1[1] ,n1572);
    not g416(n2067 ,n0[30]);
    not g417(n2079 ,n0[18]);
    xnor g418(n336 ,n308 ,n278);
    or g419(n264 ,n197 ,n253);
    or g420(n397 ,n2072 ,n2052);
    xnor g421(n96 ,n0[21] ,n0[5]);
    nand g422(n802 ,n0[61] ,n755);
    or g423(n1433 ,n1186 ,n1152);
    nor g424(n1799 ,n1733 ,n1714);
    xor g425(n945 ,n1[2] ,n1985);
    nand g426(n1545 ,n1212 ,n1380);
    nor g427(n1907 ,n3 ,n1906);
    nand g428(n354 ,n331 ,n339);
    nor g429(n1745 ,n1358 ,n1673);
    nand g430(n517 ,n482 ,n470);
    xnor g431(n107 ,n0[37] ,n0[13]);
    not g432(n740 ,n1[6]);
    nor g433(n1148 ,n976 ,n1045);
    not g434(n771 ,n5[4]);
    nand g435(n13[2] ,n1979 ,n1904);
    nand g436(n85 ,n0[30] ,n0[14]);
    nand g437(n82 ,n0[17] ,n0[1]);
    nand g438(n625 ,n569 ,n597);
    xnor g439(n900 ,n0[21] ,n0[20]);
    xnor g440(n1123 ,n885 ,n894);
    nand g441(n671 ,n649 ,n658);
    nand g442(n1342 ,n0[9] ,n1100);
    nand g443(n1664 ,n1[19] ,n1553);
    xor g444(n1990 ,n187 ,n231);
    not g445(n1256 ,n1255);
    nand g446(n37 ,n33 ,n30);
    xnor g447(n921 ,n0[24] ,n0[23]);
    not g448(n2066 ,n0[31]);
    nor g449(n1604 ,n1485 ,n1510);
    or g450(n1786 ,n1720 ,n1719);
    nor g451(n1693 ,n1650 ,n1649);
    nand g452(n544 ,n487 ,n489);
    xnor g453(n936 ,n0[40] ,n0[24]);
    xnor g454(n913 ,n0[10] ,n0[9]);
    nand g455(n1305 ,n2022 ,n1109);
    nand g456(n515 ,n481 ,n471);
    xnor g457(n647 ,n587 ,n627);
    or g458(n391 ,n2096 ,n2092);
    nand g459(n1672 ,n1531 ,n1532);
    not g460(n2097 ,n0[0]);
    xnor g461(n1260 ,n932 ,n903);
    not g462(n2072 ,n0[25]);
    nand g463(n1951 ,n1933 ,n1912);
    or g464(n65 ,n0[31] ,n0[15]);
    or g465(n384 ,n2084 ,n2035);
    or g466(n1171 ,n921 ,n1045);
    nand g467(n1488 ,n1[14] ,n1226);
    nand g468(n152 ,n85 ,n128);
    nor g469(n1360 ,n766 ,n1102);
    xnor g470(n434 ,n2038 ,n2060);
    nor g471(n1706 ,n1592 ,n1636);
    nand g472(n699 ,n682 ,n688);
    nand g473(n288 ,n240 ,n274);
    or g474(n1419 ,n1178 ,n1133);
    nor g475(n358 ,n343 ,n345);
    or g476(n63 ,n0[20] ,n0[4]);
    nand g477(n323 ,n306 ,n311);
    nor g478(n333 ,n303 ,n326);
    xnor g479(n6[57] ,n0[57] ,n1294);
    nand g480(n1211 ,n0[4] ,n1105);
    xnor g481(n280 ,n251 ,n256);
    nor g482(n950 ,n790 ,n789);
    nand g483(n317 ,n289 ,n298);
    or g484(n198 ,n159 ,n160);
    xnor g485(n1580 ,n0[5] ,n1216);
    or g486(n56 ,n0[17] ,n0[1]);
    nand g487(n141 ,n50 ,n130);
    or g488(n1462 ,n1047 ,n1257);
    nor g489(n784 ,n759 ,n1[8]);
    nor g490(n1026 ,n953 ,n955);
    nand g491(n1946 ,n1927 ,n1940);
    nor g492(n1006 ,n819 ,n966);
    nor g493(n733 ,n2017 ,n2003);
    or g494(n1187 ,n923 ,n1045);
    or g495(n1034 ,n1[19] ,n912);
    nor g496(n1626 ,n1469 ,n1503);
    nand g497(n1294 ,n2021 ,n1053);
    nor g498(n1067 ,n946 ,n957);
    nand g499(n1362 ,n1036 ,n1080);
    not g500(n642 ,n641);
    xnor g501(n168 ,n98 ,n0[28]);
    nand g502(n1389 ,n1984 ,n1054);
    xnor g503(n1914 ,n0[21] ,n1[21]);
    nor g504(n1417 ,n1330 ,n1205);
    nor g505(n1451 ,n1047 ,n1248);
    xnor g506(n426 ,n2076 ,n2079);
    nand g507(n1656 ,n1[13] ,n1553);
    nor g508(n1838 ,n1728 ,n1781);
    nand g509(n725 ,n716 ,n722);
    xnor g510(n310 ,n268 ,n281);
    or g511(n71 ,n0[22] ,n0[6]);
    nor g512(n1888 ,n1880 ,n1885);
    xnor g513(n1934 ,n0[26] ,n1[26]);
    nand g514(n1316 ,n2024 ,n1050);
    nand g515(n1151 ,n986 ,n1046);
    xnor g516(n101 ,n0[38] ,n0[14]);
    nand g517(n405 ,n2093 ,n2048);
    buf g518(n12[0], 1'b0);
    xnor g519(n1124 ,n881 ,n890);
    or g520(n1834 ,n1774 ,n1770);
    nand g521(n471 ,n414 ,n459);
    nand g522(n622 ,n594 ,n599);
    nand g523(n12[3] ,n1385 ,n1892);
    nor g524(n2108 ,n2102 ,n5[1]);
    nand g525(n547 ,n485 ,n507);
    not g526(n982 ,n981);
    nand g527(n2113 ,n2108 ,n2107);
    nor g528(n1726 ,n1559 ,n1588);
    nand g529(n641 ,n588 ,n627);
    nand g530(n17 ,n2011 ,n2005);
    or g531(n52 ,n0[24] ,n0[40]);
    nor g532(n1783 ,n1705 ,n1704);
    nand g533(n1279 ,n2021 ,n1108);
    nor g534(n1110 ,n2[3] ,n1001);
    nor g535(n13[3] ,n1899 ,n1982);
    xnor g536(n887 ,n0[17] ,n0[16]);
    nand g537(n403 ,n2090 ,n2075);
    nand g538(n1351 ,n0[21] ,n1100);
    nand g539(n638 ,n607 ,n626);
    xnor g540(n853 ,n0[57] ,n0[56]);
    or g541(n311 ,n252 ,n304);
    nand g542(n1062 ,n0[37] ,n877);
    nand g543(n832 ,n1996 ,n740);
    nand g544(n689 ,n634 ,n677);
    nand g545(n966 ,n824 ,n831);
    nand g546(n1660 ,n1403 ,n1523);
    nand g547(n1088 ,n1[19] ,n912);
    nand g548(n460 ,n2076 ,n382);
    nand g549(n50 ,n0[55] ,n0[47]);
    not g550(n775 ,n2014);
    xnor g551(n1229 ,n0[24] ,n911);
    xnor g552(n937 ,n0[24] ,n0[8]);
    xnor g553(n1793 ,n878 ,n1556);
    nand g554(n1904 ,n2003 ,n1898);
    nand g555(n2104 ,n2102 ,n2103);
    xnor g556(n925 ,n0[49] ,n0[1]);
    xnor g557(n499 ,n440 ,n2075);
    nand g558(n330 ,n300 ,n318);
    not g559(n758 ,n1[0]);
    nor g560(n809 ,n761 ,n1998);
    not g561(n2085 ,n0[12]);
    nand g562(n1370 ,n1082 ,n1063);
    nand g563(n1371 ,n1011 ,n1090);
    nor g564(n1847 ,n1601 ,n1807);
    xor g565(n1236 ,n0[2] ,n868);
    nand g566(n1535 ,n1213 ,n1338);
    xnor g567(n489 ,n429 ,n2052);
    nand g568(n808 ,n771 ,n772);
    xnor g569(n870 ,n0[54] ,n0[22]);
    xnor g570(n159 ,n97 ,n0[45]);
    xnor g571(n2005 ,n1[0] ,n1575);
    nor g572(n1596 ,n1537 ,n1402);
    nand g573(n1942 ,n1919 ,n1914);
    nand g574(n569 ,n512 ,n549);
    nand g575(n1330 ,n1007 ,n1065);
    nand g576(n609 ,n575 ,n585);
    or g577(n7[24] ,n1156 ,n1767);
    nand g578(n1676 ,n1[26] ,n1553);
    nand g579(n1764 ,n1679 ,n1184);
    nor g580(n1832 ,n1810 ,n1817);
    or g581(n38 ,n35 ,n34);
    not g582(n2083 ,n0[14]);
    or g583(n361 ,n353 ,n345);
    not g584(n886 ,n887);
    xnor g585(n6[44] ,n0[44] ,n1322);
    nor g586(n672 ,n595 ,n660);
    nand g587(n25 ,n17 ,n23);
    xnor g588(n6[37] ,n0[37] ,n1272);
    xnor g589(n115 ,n0[58] ,n0[50]);
    xnor g590(n488 ,n437 ,n444);
    nand g591(n793 ,n0[62] ,n740);
    or g592(n193 ,n154 ,n170);
    xnor g593(n634 ,n592 ,n597);
    xnor g594(n190 ,n141 ,n142);
    nand g595(n1080 ,n1[15] ,n922);
    xnor g596(n857 ,n0[33] ,n0[32]);
    not g597(n2086 ,n0[11]);
    nand g598(n1162 ,n891 ,n1046);
    nand g599(n1191 ,n1004 ,n1026);
    nand g600(n343 ,n303 ,n326);
    xnor g601(n433 ,n2095 ,n2036);
    nand g602(n1638 ,n1528 ,n1439);
    nand g603(n228 ,n174 ,n199);
    nor g604(n1018 ,n878 ,n876);
    or g605(n400 ,n2083 ,n2067);
    not g606(n879 ,n878);
    nand g607(n185 ,n51 ,n148);
    nand g608(n1531 ,n1[20] ,n1228);
    xnor g609(n251 ,n190 ,n217);
    nand g610(n273 ,n256 ,n251);
    or g611(n831 ,n755 ,n1988);
    nand g612(n408 ,n2069 ,n2059);
    nand g613(n1500 ,n1336 ,n1146);
    xnor g614(n1117 ,n874 ,n845);
    nor g615(n1819 ,n993 ,n1741);
    xnor g616(n1128 ,n869 ,n857);
    nor g617(n1852 ,n1789 ,n1788);
    xnor g618(n191 ,n143 ,n116);
    xnor g619(n890 ,n0[9] ,n0[8]);
    nand g620(n1952 ,n1939 ,n1938);
    not g621(n774 ,n4[1]);
    xnor g622(n938 ,n0[37] ,n0[36]);
    xnor g623(n6[17] ,n0[17] ,n1321);
    nand g624(n410 ,n2072 ,n2052);
    nand g625(n26 ,n18 ,n24);
    not g626(n2069 ,n0[28]);
    xnor g627(n959 ,n1[4] ,n1994);
    nand g628(n1517 ,n1[6] ,n1240);
    nor g629(n1735 ,n1663 ,n1602);
    nand g630(n1311 ,n2027 ,n1109);
    xnor g631(n929 ,n0[38] ,n0[22]);
    nand g632(n1588 ,n1471 ,n1473);
    not g633(n2062 ,n0[35]);
    nor g634(n810 ,n745 ,n1999);
    not g635(n1259 ,n1258);
    nand g636(n734 ,n2018 ,n2019);
    xor g637(n1237 ,n0[45] ,n924);
    nand g638(n12[4] ,n1386 ,n1881);
    not g639(n764 ,n0[25]);
    xnor g640(n600 ,n556 ,n488);
    xnor g641(n1987 ,n726 ,n729);
    not g642(n2093 ,n0[4]);
    nand g643(n1355 ,n1042 ,n1061);
    or g644(n506 ,n467 ,n472);
    xnor g645(n848 ,n0[33] ,n0[17]);
    or g646(n1027 ,n1[14] ,n885);
    or g647(n688 ,n634 ,n677);
    xnor g648(n527 ,n481 ,n471);
    nand g649(n822 ,n1993 ,n742);
    xnor g650(n1233 ,n937 ,n905);
    nor g651(n2012 ,n47 ,n49);
    nand g652(n256 ,n209 ,n228);
    xnor g653(n528 ,n485 ,n478);
    or g654(n1784 ,n1732 ,n1736);
    or g655(n7[28] ,n1159 ,n1768);
    xnor g656(n894 ,n0[11] ,n0[10]);
    or g657(n1103 ,n834 ,n990);
    xnor g658(n1921 ,n0[28] ,n1[28]);
    or g659(n717 ,n710 ,n711);
    nand g660(n1757 ,n1640 ,n1455);
    xnor g661(n926 ,n0[27] ,n0[3]);
    nand g662(n182 ,n63 ,n146);
    xnor g663(n1129 ,n896 ,n898);
    nor g664(n1709 ,n1657 ,n1587);
    or g665(n1190 ,n1103 ,n1023);
    nand g666(n954 ,n794 ,n783);
    xnor g667(n1996 ,n362 ,n370);
    xnor g668(n313 ,n280 ,n290);
    nand g669(n1287 ,n2027 ,n1051);
    not g670(n766 ,n0[56]);
    xnor g671(n919 ,n0[14] ,n0[13]);
    nand g672(n794 ,n0[63] ,n743);
    xnor g673(n1937 ,n0[22] ,n1[22]);
    nand g674(n33 ,n19 ,n31);
    xnor g675(n309 ,n267 ,n284);
    not g676(n2048 ,n0[49]);
    xor g677(n30 ,n26 ,n25);
    or g678(n659 ,n653 ,n647);
    or g679(n1483 ,n989 ,n1382);
    not g680(n2038 ,n0[59]);
    xnor g681(n661 ,n629 ,n596);
    nand g682(n242 ,n179 ,n204);
    or g683(n1017 ,n1[28] ,n893);
    xnor g684(n984 ,n0[4] ,n0[3]);
    xnor g685(n1985 ,n719 ,n713);
    xor g686(n1248 ,n0[47] ,n935);
    xnor g687(n1571 ,n0[1] ,n1223);
    xnor g688(n1582 ,n1127 ,n1118);
    xnor g689(n518 ,n439 ,n2094);
    xnor g690(n646 ,n613 ,n586);
    nand g691(n461 ,n2066 ,n400);
    xnor g692(n1558 ,n1[4] ,n1260);
    or g693(n1830 ,n2011 ,n2005);
    xnor g694(n437 ,n2088 ,n2087);
    nand g695(n153 ,n92 ,n137);
    nor g696(n1969 ,n1965 ,n3);
    or g697(n1059 ,n755 ,n982);
    or g698(n16 ,n2009 ,n2008);
    nand g699(n837 ,n2002 ,n2001);
    xnor g700(n1924 ,n0[10] ,n1[10]);
    nor g701(n1054 ,n835 ,n993);
    nand g702(n274 ,n237 ,n259);
    or g703(n1602 ,n1421 ,n1422);
    nor g704(n1511 ,n1[23] ,n1248);
    nor g705(n1415 ,n1363 ,n1131);
    nand g706(n1481 ,n745 ,n1255);
    or g707(n7[11] ,n1758 ,n1849);
    or g708(n64 ,n0[60] ,n0[44]);
    nand g709(n666 ,n639 ,n651);
    xor g710(n1916 ,n0[15] ,n1[15]);
    xnor g711(n1247 ,n0[11] ,n871);
    nor g712(n1198 ,n757 ,n1104);
    xnor g713(n6[30] ,n0[30] ,n1284);
    xnor g714(n846 ,n0[35] ,n0[19]);
    not g715(n2064 ,n0[33]);
    or g716(n68 ,n0[28] ,n0[12]);
    nand g717(n620 ,n591 ,n610);
    nand g718(n420 ,n2085 ,n2055);
    nand g719(n482 ,n420 ,n465);
    xnor g720(n268 ,n219 ,n170);
    nand g721(n586 ,n540 ,n563);
    nor g722(n1166 ,n1069 ,n1016);
    or g723(n974 ,n806 ,n805);
    xnor g724(n6[29] ,n0[29] ,n1286);
    nor g725(n1207 ,n1[11] ,n1029);
    or g726(n1425 ,n810 ,n1329);
    or g727(n295 ,n268 ,n281);
    nor g728(n1100 ,n835 ,n989);
    xnor g729(n1933 ,n0[2] ,n1[2]);
    nand g730(n1890 ,n1855 ,n1887);
    nand g731(n1403 ,n879 ,n1222);
    nor g732(n2105 ,n2029 ,n5[1]);
    xnor g733(n1926 ,n0[17] ,n1[17]);
    nor g734(n1484 ,n1[14] ,n1226);
    not g735(n1792 ,n2011);
    not g736(n2101 ,n5[0]);
    xnor g737(n438 ,n2039 ,n2045);
    nand g738(n828 ,n1987 ,n739);
    xnor g739(n6[36] ,n0[36] ,n1274);
    xnor g740(n1240 ,n929 ,n901);
    xor g741(n1559 ,n1[17] ,n1225);
    nand g742(n1845 ,n1166 ,n1780);
    nand g743(n1677 ,n1[27] ,n1553);
    nand g744(n7[7] ,n1681 ,n1846);
    nand g745(n970 ,n828 ,n820);
    nand g746(n147 ,n87 ,n131);
    or g747(n1445 ,n756 ,n1232);
    xnor g748(n864 ,n0[49] ,n0[48]);
    nor g749(n2098 ,n1830 ,n737);
    nand g750(n955 ,n793 ,n786);
    xnor g751(n928 ,n0[59] ,n0[58]);
    nand g752(n1303 ,n2027 ,n1049);
    not g753(n768 ,n0[31]);
    not g754(n765 ,n0[30]);
    nor g755(n1215 ,n988 ,n1104);
    not g756(n891 ,n892);
    xnor g757(n441 ,n2084 ,n2062);
    xnor g758(n299 ,n263 ,n269);
    xnor g759(n1115 ,n978 ,n985);
    xnor g760(n628 ,n594 ,n601);
    nand g761(n1520 ,n1192 ,n1200);
    nor g762(n1662 ,n1339 ,n1426);
    nand g763(n1766 ,n1680 ,n1179);
    xnor g764(n282 ,n248 ,n259);
    nor g765(n35 ,n33 ,n30);
    xnor g766(n503 ,n426 ,n2078);
    or g767(n67 ,n0[55] ,n0[47]);
    not g768(n2046 ,n0[51]);
    or g769(n1833 ,n1102 ,n1793);
    xnor g770(n1994 ,n350 ,n365);
    nand g771(n1300 ,n2024 ,n1049);
    nor g772(n1654 ,n1520 ,n1433);
    nand g773(n1470 ,n743 ,n1253);
    or g774(n275 ,n256 ,n251);
    nand g775(n1818 ,n1751 ,n1703);
    xnor g776(n845 ,n0[46] ,n0[41]);
    nor g777(n1741 ,n1028 ,n1627);
    nand g778(n1293 ,n2021 ,n1107);
    nand g779(n205 ,n139 ,n168);
    xnor g780(n1773 ,n1[1] ,n1571);
    nand g781(n145 ,n75 ,n132);
    xnor g782(n1135 ,n1[24] ,n888);
    or g783(n9 ,n2100 ,n1907);
    nand g784(n320 ,n273 ,n301);
    xnor g785(n6[38] ,n0[38] ,n1271);
    nand g786(n1439 ,n755 ,n1252);
    nand g787(n462 ,n2082 ,n401);
    nand g788(n301 ,n290 ,n275);
    nand g789(n1361 ,n0[63] ,n1101);
    nor g790(n1727 ,n1651 ,n1564);
    nand g791(n1947 ,n1926 ,n1923);
    xnor g792(n1131 ,n1[9] ,n913);
    nand g793(n1071 ,n875 ,n959);
    or g794(n399 ,n2085 ,n2055);
    xor g795(n314 ,n279 ,n270);
    nand g796(n137 ,n0[2] ,n69);
    nand g797(n1331 ,n1017 ,n1064);
    nor g798(n1723 ,n1103 ,n1569);
    nand g799(n1805 ,n1727 ,n1693);
    nand g800(n1209 ,n0[22] ,n1100);
    nor g801(n781 ,n744 ,n1[10]);
    not g802(n757 ,n0[2]);
    or g803(n15 ,n2011 ,n2005);
    nor g804(n1780 ,n1191 ,n1690);
    xnor g805(n435 ,n2071 ,n2034);
    nand g806(n370 ,n364 ,n368);
    xnor g807(n614 ,n576 ,n589);
    nand g808(n1350 ,n0[8] ,n1100);
    nor g809(n1343 ,n765 ,n1099);
    not g810(n2060 ,n0[37]);
    nand g811(n24 ,n2006 ,n14);
    xnor g812(n1563 ,n1[12] ,n1241);
    xnor g813(n2030 ,n0[0] ,n1[0]);
    nor g814(n1469 ,n1047 ,n1236);
    not g815(n2053 ,n0[44]);
    nor g816(n1878 ,n2007 ,n1869);
    xnor g817(n118 ,n0[48] ,n0[16]);
    nand g818(n321 ,n291 ,n299);
    nand g819(n1443 ,n1[4] ,n1245);
    nand g820(n1264 ,n2026 ,n1052);
    nand g821(n1668 ,n1[23] ,n1553);
    nor g822(n1486 ,n1[12] ,n1239);
    nand g823(n1153 ,n982 ,n1046);
    nand g824(n1346 ,n0[27] ,n1100);
    xnor g825(n1986 ,n727 ,n725);
    not g826(n732 ,n731);
    nand g827(n606 ,n580 ,n579);
    or g828(n1513 ,n1[19] ,n1246);
    or g829(n287 ,n271 ,n270);
    xnor g830(n1578 ,n1224 ,n1218);
    xnor g831(n867 ,n0[39] ,n0[38]);
    nand g832(n964 ,n2[0] ,n807);
    xnor g833(n6[21] ,n0[21] ,n1301);
    nand g834(n374 ,n355 ,n371);
    nand g835(n409 ,n2083 ,n2067);
    nand g836(n93 ,n0[31] ,n0[15]);
    xnor g837(n916 ,n0[22] ,n0[21]);
    nor g838(n1869 ,n2008 ,n1860);
    not g839(n1898 ,n1982);
    nor g840(n1493 ,n0[37] ,n1222);
    nand g841(n217 ,n81 ,n185);
    xnor g842(n883 ,n0[19] ,n0[18]);
    nand g843(n1630 ,n1[2] ,n1553);
    not g844(n2045 ,n0[52]);
    xnor g845(n224 ,n151 ,n166);
    nand g846(n8 ,n2099 ,n1972);
    nand g847(n13[0] ,n1980 ,n1902);
    nand g848(n1061 ,n1[7] ,n988);
    xnor g849(n1239 ,n849 ,n749);
    nand g850(n1482 ,n1201 ,n1150);
    nor g851(n1696 ,n1102 ,n1567);
    not g852(n2102 ,n5[2]);
    xnor g853(n859 ,n0[26] ,n0[10]);
    or g854(n1778 ,n1474 ,n1761);
    xnor g855(n668 ,n654 ,n655);
    nand g856(n7[9] ,n1695 ,n1858);
    xor g857(n1242 ,n0[46] ,n934);
    xnor g858(n909 ,n0[38] ,n0[14]);
    nand g859(n815 ,n1995 ,n755);
    nand g860(n411 ,n2068 ,n2064);
    nor g861(n1628 ,n740 ,n1552);
    nor g862(n1717 ,n1102 ,n1578);
    not g863(n2036 ,n0[61]);
    xnor g864(n1935 ,n0[19] ,n1[19]);
    nand g865(n1540 ,n2030 ,n1138);
    or g866(n1781 ,n1697 ,n1696);
    not g867(n769 ,n3);
    xnor g868(n445 ,n2093 ,n2047);
    xnor g869(n1127 ,n858 ,n928);
    nand g870(n1317 ,n2025 ,n1050);
    nand g871(n356 ,n346 ,n348);
    xnor g872(n1999 ,n341 ,n378);
    xnor g873(n6[59] ,n0[59] ,n1269);
    xnor g874(n6[12] ,n0[12] ,n1316);
    not g875(n2044 ,n0[53]);
    nand g876(n709 ,n690 ,n701);
    xnor g877(n1930 ,n0[18] ,n1[18]);
    or g878(n1607 ,n1444 ,n1493);
    xnor g879(n6[22] ,n0[22] ,n1302);
    nor g880(n1178 ,n998 ,n1044);
    nand g881(n255 ,n242 ,n230);
    xnor g882(n901 ,n0[54] ,n0[6]);
    or g883(n382 ,n2079 ,n2078);
    xnor g884(n599 ,n552 ,n500);
    nand g885(n412 ,n2041 ,n2044);
    nand g886(n1769 ,n1346 ,n1677);
    xnor g887(n1556 ,n0[13] ,n1216);
    or g888(n1963 ,n1931 ,n1958);
    nor g889(n1738 ,n1658 ,n1607);
    nand g890(n1640 ,n1[9] ,n1553);
    nand g891(n1502 ,n1335 ,n1187);
    nand g892(n1341 ,n0[12] ,n1100);
    or g893(n1031 ,n1[12] ,n881);
    nor g894(n798 ,n739 ,n0[60]);
    nand g895(n1212 ,n0[5] ,n1105);
    nor g896(n1829 ,n1653 ,n1819);
    xnor g897(n6[50] ,n0[50] ,n1280);
    nand g898(n730 ,n720 ,n729);
    nand g899(n1977 ,n807 ,n1110);
    nand g900(n550 ,n486 ,n508);
    nand g901(n1292 ,n2020 ,n1053);
    nand g902(n7[17] ,n1670 ,n1625);
    nand g903(n1765 ,n1634 ,n1157);
    nand g904(n973 ,n814 ,n818);
    nor g905(n2020 ,n5[0] ,n2104);
    nand g906(n1504 ,n1333 ,n1189);
    nand g907(n565 ,n477 ,n537);
    xnor g908(n6[43] ,n0[43] ,n1323);
    xnor g909(n648 ,n614 ,n578);
    nor g910(n1204 ,n1025 ,n1073);
    xnor g911(n978 ,n0[7] ,n0[6]);
    nand g912(n123 ,n0[54] ,n62);
    or g913(n55 ,n0[21] ,n0[5]);
    nand g914(n1076 ,n1[12] ,n881);
    nand g915(n327 ,n307 ,n314);
    xnor g916(n6[10] ,n0[10] ,n1314);
    xnor g917(n1581 ,n1130 ,n907);
    nor g918(n1427 ,n1206 ,n1369);
    nand g919(n1394 ,n1986 ,n1054);
    xnor g920(n1579 ,n1122 ,n908);
    or g921(n51 ,n0[23] ,n0[7]);
    nand g922(n1746 ,n1[10] ,n1577);
    nand g923(n474 ,n390 ,n446);
    not g924(n41 ,n40);
    not g925(n2091 ,n0[6]);
    nand g926(n700 ,n687 ,n686);
    or g927(n1465 ,n1047 ,n1228);
    nor g928(n1509 ,n1[21] ,n1237);
    nand g929(n1392 ,n1985 ,n1054);
    xnor g930(n500 ,n433 ,n2073);
    nand g931(n7[12] ,n1711 ,n1813);
    not g932(n975 ,n976);
    xnor g933(n1116 ,n980 ,n976);
    nor g934(n1452 ,n1047 ,n1227);
    nor g935(n1044 ,n739 ,n1000);
    nand g936(n1335 ,n0[17] ,n1100);
    or g937(n7[31] ,n1340 ,n1766);
    xnor g938(n649 ,n612 ,n580);
    xnor g939(n439 ,n2077 ,n2089);
    nand g940(n1749 ,n1[12] ,n1581);
    nand g941(n2110 ,n2028 ,n2103);
    xnor g942(n1576 ,n1114 ,n1120);
    or g943(n227 ,n213 ,n200);
    nor g944(n1137 ,n792 ,n1038);
    nand g945(n1325 ,n2024 ,n1053);
    nor g946(n952 ,n798 ,n795);
    nor g947(n1891 ,n843 ,n1888);
    xnor g948(n6[11] ,n0[11] ,n1315);
    xnor g949(n1231 ,n925 ,n764);
    nand g950(n1461 ,n1048 ,n1225);
    nor g951(n1406 ,n1366 ,n1327);
    nand g952(n80 ,n0[29] ,n0[13]);
    nand g953(n1315 ,n2023 ,n1050);
    nand g954(n1811 ,n1738 ,n1709);
    xnor g955(n114 ,n0[62] ,n0[54]);
    nand g956(n422 ,n2042 ,n2043);
    nand g957(n450 ,n2051 ,n397);
    nor g958(n1848 ,n1820 ,n1782);
    nand g959(n303 ,n276 ,n287);
    nor g960(n1109 ,n808 ,n995);
    nor g961(n59 ,n0[19] ,n0[3]);
    nand g962(n1066 ,n1[15] ,n988);
    nand g963(n1505 ,n0[37] ,n1222);
    nand g964(n1632 ,n1[4] ,n1553);
    or g965(n1168 ,n1008 ,n1014);
    not g966(n1245 ,n1244);
    nand g967(n1622 ,n1459 ,n1429);
    xnor g968(n924 ,n0[21] ,n0[1]);
    nand g969(n1288 ,n2024 ,n1107);
    nand g970(n1359 ,n0[57] ,n1101);
    nand g971(n650 ,n633 ,n637);
    or g972(n1695 ,n1103 ,n1571);
    xnor g973(n250 ,n189 ,n186);
    xnor g974(n1243 ,n927 ,n908);
    nor g975(n1025 ,n1[1] ,n996);
    xnor g976(n1249 ,n933 ,n911);
    or g977(n53 ,n0[42] ,n0[10]);
    nor g978(n2016 ,n1943 ,n1962);
    not g979(n1976 ,n2002);
    nand g980(n621 ,n590 ,n603);
    nand g981(n7[18] ,n1671 ,n1626);
    or g982(n698 ,n687 ,n686);
    xnor g983(n939 ,n0[47] ,n0[40]);
    nor g984(n1049 ,n838 ,n995);
    or g985(n1598 ,n1508 ,n1407);
    or g986(n1707 ,n1637 ,n1590);
    xnor g987(n962 ,n1[7] ,n1997);
    xnor g988(n202 ,n109 ,n146);
    nand g989(n1267 ,n2025 ,n1052);
    nand g990(n1767 ,n1208 ,n1674);
    nand g991(n365 ,n327 ,n360);
    not g992(n2087 ,n0[10]);
    nand g993(n149 ,n94 ,n115);
    xnor g994(n1586 ,n0[2] ,n1217);
    xnor g995(n493 ,n432 ,n2057);
    xnor g996(n170 ,n101 ,n0[30]);
    xnor g997(n903 ,n0[52] ,n0[36]);
    nor g998(n2021 ,n2106 ,n2104);
    xnor g999(n1993 ,n340 ,n349);
    nand g1000(n1356 ,n0[6] ,n1100);
    xnor g1001(n6[41] ,n0[41] ,n1263);
    or g1002(n1713 ,n1103 ,n1580);
    nand g1003(n1729 ,n1506 ,n1621);
    nand g1004(n958 ,n821 ,n822);
    nor g1005(n359 ,n354 ,n347);
    not g1006(n840 ,n839);
    nand g1007(n286 ,n249 ,n269);
    xnor g1008(n6[26] ,n0[26] ,n1291);
    nand g1009(n485 ,n411 ,n456);
    xnor g1010(n1241 ,n931 ,n907);
    nor g1011(n1353 ,n767 ,n1099);
    not g1012(n877 ,n876);
    nor g1013(n1413 ,n1175 ,n1331);
    nand g1014(n1760 ,n1341 ,n1643);
    nand g1015(n2024 ,n2124 ,n2125);
    nand g1016(n691 ,n655 ,n681);
    nand g1017(n1537 ,n1374 ,n1147);
    or g1018(n1836 ,n2007 ,n2008);
    nand g1019(n723 ,n705 ,n718);
    xnor g1020(n99 ,n0[60] ,n0[52]);
    or g1021(n312 ,n291 ,n299);
    nand g1022(n1321 ,n2021 ,n1049);
    xnor g1023(n169 ,n112 ,n0[1]);
    or g1024(n199 ,n152 ,n167);
    not g1025(n117 ,n116);
    nand g1026(n835 ,n2[0] ,n3);
    nand g1027(n1329 ,n1067 ,n1072);
    nor g1028(n1618 ,n1453 ,n1491);
    or g1029(n603 ,n575 ,n585);
    xnor g1030(n1927 ,n0[31] ,n1[31]);
    nand g1031(n582 ,n520 ,n566);
    or g1032(n1184 ,n920 ,n1045);
    xnor g1033(n22 ,n2009 ,n2008);
    or g1034(n396 ,n2090 ,n2075);
    or g1035(n1420 ,n1[9] ,n1234);
    xnor g1036(n613 ,n577 ,n584);
    nand g1037(n315 ,n306 ,n305);
    xor g1038(n1228 ,n0[0] ,n906);
    not g1039(n770 ,n2[3]);
    not g1040(n1965 ,n2033);
    nand g1041(n1369 ,n1085 ,n1059);
    nand g1042(n1882 ,n1856 ,n1875);
    nand g1043(n708 ,n700 ,n698);
    nand g1044(n1165 ,n882 ,n1046);
    xnor g1045(n933 ,n0[32] ,n0[16]);
    nand g1046(n1324 ,n2026 ,n1051);
    nand g1047(n1479 ,n1[8] ,n1227);
    xnor g1048(n1568 ,n1112 ,n1128);
    nor g1049(n387 ,n2088 ,n2087);
    xnor g1050(n1920 ,n0[14] ,n1[14]);
    nand g1051(n821 ,n1998 ,n761);
    xnor g1052(n645 ,n615 ,n575);
    xnor g1053(n856 ,n0[50] ,n0[18]);
    nand g1054(n719 ,n716 ,n717);
    nand g1055(n1210 ,n0[16] ,n1100);
    nand g1056(n1380 ,n2000 ,n1106);
    nand g1057(n1091 ,n829 ,n944);
    xnor g1058(n160 ,n107 ,n0[29]);
    xnor g1059(n6[52] ,n0[52] ,n1273);
    xnor g1060(n863 ,n0[37] ,n0[21]);
    nand g1061(n1086 ,n1[17] ,n923);
    xnor g1062(n529 ,n480 ,n468);
    xnor g1063(n1919 ,n0[23] ,n1[23]);
    nor g1064(n1358 ,n749 ,n1102);
    not g1065(n983 ,n984);
    xnor g1066(n269 ,n224 ,n171);
    nand g1067(n706 ,n692 ,n698);
    xnor g1068(n220 ,n169 ,n165);
    or g1069(n293 ,n265 ,n283);
    nor g1070(n790 ,n748 ,n0[7]);
    nand g1071(n1262 ,n2022 ,n1051);
    not g1072(n2047 ,n0[50]);
    nand g1073(n1295 ,n2025 ,n1051);
    xnor g1074(n593 ,n568 ,n567);
    nand g1075(n1093 ,n1[30] ,n896);
    nand g1076(n520 ,n421 ,n466);
    nor g1077(n2109 ,n2103 ,n2028);
    nand g1078(n78 ,n0[24] ,n0[40]);
    xnor g1079(n1569 ,n0[59] ,n1219);
    nor g1080(n345 ,n328 ,n336);
    xnor g1081(n1573 ,n1125 ,n1126);
    nor g1082(n2126 ,n2115 ,n2123);
    nand g1083(n402 ,n2040 ,n2081);
    nor g1084(n1856 ,n1845 ,n1772);
    nand g1085(n1374 ,n1989 ,n1054);
    nand g1086(n1195 ,n0[3] ,n1105);
    nand g1087(n1591 ,n1481 ,n1487);
    xnor g1088(n502 ,n434 ,n2061);
    not g1089(n881 ,n880);
    or g1090(n816 ,n740 ,n1996);
    nand g1091(n126 ,n0[36] ,n68);
    nand g1092(n997 ,n2013 ,n775);
    xnor g1093(n6[1] ,n0[1] ,n1304);
    nand g1094(n1399 ,n1988 ,n1054);
    nand g1095(n1639 ,n1[8] ,n1553);
    xnor g1096(n6[48] ,n0[48] ,n1285);
    nand g1097(n1874 ,n992 ,n1865);
    nand g1098(n1644 ,n1[14] ,n1553);
    or g1099(n2121 ,n2105 ,n2117);
    nand g1100(n1334 ,n0[18] ,n1100);
    nand g1101(n1593 ,n1488 ,n1438);
    nor g1102(n780 ,n740 ,n0[3]);
    nor g1103(n1056 ,n843 ,n989);
    nand g1104(n94 ,n0[57] ,n0[49]);
    nor g1105(n1405 ,n1355 ,n1326);
    nand g1106(n1612 ,n1505 ,n1513);
    nand g1107(n40 ,n37 ,n38);
    nor g1108(n1053 ,n844 ,n994);
    or g1109(n1782 ,n1701 ,n1702);
    nand g1110(n1280 ,n2022 ,n1052);
    nand g1111(n1733 ,n1644 ,n1163);
    nor g1112(n948 ,n777 ,n779);
    xnor g1113(n875 ,n1[10] ,n2000);
    nand g1114(n418 ,n2039 ,n2046);
    nand g1115(n727 ,n724 ,n721);
    nand g1116(n627 ,n583 ,n602);
    nand g1117(n13[1] ,n1978 ,n1903);
    or g1118(n192 ,n151 ,n166);
    nand g1119(n585 ,n543 ,n558);
    nor g1120(n1814 ,n1524 ,n1753);
    nand g1121(n1069 ,n943 ,n961);
    nor g1122(n1013 ,n1[20] ,n900);
    xnor g1123(n1940 ,n0[30] ,n1[30]);
    nor g1124(n1052 ,n838 ,n994);
    xnor g1125(n1255 ,n0[57] ,n854);
    xnor g1126(n553 ,n505 ,n498);
    or g1127(n176 ,n153 ,n150);
    nand g1128(n570 ,n513 ,n546);
    xnor g1129(n1223 ,n0[49] ,n848);
    nand g1130(n1319 ,n2027 ,n1050);
    xnor g1131(n865 ,n0[45] ,n0[44]);
    or g1132(n534 ,n499 ,n497);
    or g1133(n1175 ,n1012 ,n1019);
    nor g1134(n2119 ,n2109 ,n2112);
    xnor g1135(n1217 ,n0[34] ,n856);
    nor g1136(n833 ,n769 ,n2[0]);
    nand g1137(n89 ,n0[27] ,n0[11]);
    nor g1138(n1466 ,n1047 ,n1230);
    not g1139(n2040 ,n0[57]);
    nand g1140(n1646 ,n1427 ,n1405);
    or g1141(n177 ,n141 ,n142);
    nand g1142(n1372 ,n1020 ,n1097);
    nor g1143(n1519 ,n1[8] ,n1227);
    xnor g1144(n248 ,n214 ,n201);
    xnor g1145(n695 ,n674 ,n679);
    nor g1146(n1827 ,n1785 ,n1729);
    xnor g1147(n246 ,n215 ,n203);
    nand g1148(n1164 ,n886 ,n1046);
    nor g1149(n1155 ,n894 ,n1045);
    not g1150(n979 ,n980);
    nand g1151(n1087 ,n1[23] ,n921);
    nand g1152(n1157 ,n895 ,n1046);
    or g1153(n1424 ,n1103 ,n1260);
    xnor g1154(n440 ,n2074 ,n2090);
    nand g1155(n464 ,n2045 ,n389);
    nand g1156(n1385 ,n972 ,n1056);
    nand g1157(n1631 ,n1[3] ,n1553);
    nor g1158(n1186 ,n996 ,n1104);
    nor g1159(n1410 ,n1395 ,n1357);
    nand g1160(n1021 ,n763 ,n982);
    or g1161(n1189 ,n912 ,n1045);
    nor g1162(n776 ,n1[13] ,n1[12]);
    nand g1163(n1085 ,n1[16] ,n887);
    nand g1164(n453 ,n2047 ,n388);
    nand g1165(n1648 ,n1409 ,n1408);
    nor g1166(n2001 ,n1949 ,n1963);
    nand g1167(n1201 ,n0[7] ,n1100);
    not g1168(n522 ,n521);
    nand g1169(n1313 ,n2021 ,n1050);
    or g1170(n680 ,n661 ,n672);
    nand g1171(n7[23] ,n1668 ,n1619);
    nand g1172(n7[13] ,n1833 ,n1840);
    xnor g1173(n188 ,n0[32] ,n118);
    not g1174(n898 ,n897);
    nor g1175(n1840 ,n1816 ,n1756);
    not g1176(n977 ,n978);
    nand g1177(n413 ,n2071 ,n2053);
    or g1178(n1177 ,n917 ,n1045);
    xnor g1179(n999 ,n0[3] ,n755);
    not g1180(n991 ,n992);
    xnor g1181(n1912 ,n0[1] ,n1[1]);
    nand g1182(n1817 ,n1747 ,n1688);
    nand g1183(n1271 ,n2026 ,n1108);
    nand g1184(n127 ,n0[35] ,n58);
    nand g1185(n665 ,n640 ,n644);
    nand g1186(n150 ,n73 ,n135);
    nand g1187(n654 ,n622 ,n631);
    nand g1188(n1282 ,n2021 ,n1052);
    xnor g1189(n715 ,n704 ,n707);
    xnor g1190(n6[24] ,n0[24] ,n1296);
    nor g1191(n1603 ,n1509 ,n1484);
    xnor g1192(n615 ,n590 ,n585);
    not g1193(n2084 ,n0[13]);
    nand g1194(n421 ,n2088 ,n2087);
    nor g1195(n1831 ,n1792 ,n2010);
    or g1196(n1423 ,n1[14] ,n1243);
    or g1197(n957 ,n809 ,n813);
    xnor g1198(n110 ,n0[41] ,n0[9]);
    or g1199(n1961 ,n1910 ,n1960);
    or g1200(n1176 ,n1040 ,n1013);
    nand g1201(n1944 ,n1915 ,n1925);
    or g1202(n69 ,n0[26] ,n0[18]);
    not g1203(n1966 ,n2031);
    nor g1204(n1012 ,n1[17] ,n923);
    nor g1205(n961 ,n799 ,n801);
    nand g1206(n175 ,n153 ,n150);
    xnor g1207(n2007 ,n1[5] ,n1565);
    nand g1208(n1375 ,n1996 ,n1106);
    nand g1209(n1208 ,n0[24] ,n1100);
    nor g1210(n1712 ,n1[12] ,n1581);
    nor g1211(n1905 ,n1900 ,n2019);
    nand g1212(n1471 ,n1[7] ,n1254);
    nand g1213(n1587 ,n1443 ,n1442);
    nand g1214(n1681 ,n1[7] ,n1553);
    nand g1215(n1476 ,n947 ,n1137);
    nor g1216(n1444 ,n1[2] ,n1236);
    nand g1217(n261 ,n208 ,n235);
    nand g1218(n1544 ,n1195 ,n1375);
    nand g1219(n1377 ,n1095 ,n1093);
    xnor g1220(n267 ,n221 ,n167);
    xnor g1221(n677 ,n656 ,n639);
    nand g1222(n83 ,n0[28] ,n0[12]);
    nand g1223(n362 ,n354 ,n346);
    nand g1224(n1276 ,n2023 ,n1108);
    not g1225(n2057 ,n0[40]);
    nand g1226(n1291 ,n2022 ,n1107);
    nor g1227(n1895 ,n1886 ,n1894);
    xnor g1228(n6[62] ,n0[62] ,n1270);
    nor g1229(n1015 ,n1[29] ,n920);
    nand g1230(n2033 ,n734 ,n733);
    or g1231(n7[4] ,n1853 ,n1797);
    nand g1232(n1808 ,n1699 ,n1698);
    not g1233(n2073 ,n0[24]);
    or g1234(n511 ,n480 ,n468);
    nand g1235(n662 ,n632 ,n648);
    xnor g1236(n100 ,n0[63] ,n0[55]);
    or g1237(n812 ,n758 ,n1990);
    not g1238(n2074 ,n0[23]);
    or g1239(n238 ,n215 ,n203);
    not g1240(n1477 ,n1447);
    xnor g1241(n27 ,n21 ,n2007);
    or g1242(n690 ,n674 ,n679);
    nand g1243(n1379 ,n1087 ,n1083);
    nand g1244(n589 ,n544 ,n564);
    nand g1245(n542 ,n493 ,n498);
    or g1246(n788 ,n741 ,n0[58]);
    nand g1247(n1678 ,n1[28] ,n1553);
    nand g1248(n1980 ,n2014 ,n1056);
    not g1249(n1111 ,n1110);
    not g1250(n1899 ,n2017);
    xnor g1251(n1997 ,n363 ,n376);
    nor g1252(n1956 ,n1948 ,n1947);
    nor g1253(n1048 ,n835 ,n990);
    not g1254(n2082 ,n0[15]);
    xnor g1255(n1918 ,n0[13] ,n1[13]);
    nand g1256(n682 ,n663 ,n671);
    xnor g1257(n1585 ,n1220 ,n1219);
    or g1258(n1954 ,n1944 ,n1950);
    nor g1259(n792 ,n747 ,n1[12]);
    not g1260(n2096 ,n0[1]);
    nand g1261(n1661 ,n1525 ,n1420);
    nor g1262(n1702 ,n1[15] ,n1583);
    xnor g1263(n1932 ,n0[5] ,n1[5]);
    nand g1264(n7[0] ,n1683 ,n1827);
    xnor g1265(n492 ,n442 ,n2059);
    nor g1266(n813 ,n755 ,n1995);
    nand g1267(n1058 ,n1[2] ,n985);
    or g1268(n1042 ,n1[18] ,n883);
    not g1269(n1000 ,n999);
    or g1270(n1688 ,n1[15] ,n1578);
    not g1271(n756 ,n1[1]);
    nand g1272(n1075 ,n1[14] ,n885);
    nor g1273(n1842 ,n1802 ,n1784);
    or g1274(n14 ,n2010 ,n2007);
    not g1275(n2090 ,n0[7]);
    nand g1276(n800 ,n0[60] ,n739);
    xor g1277(n1928 ,n0[3] ,n1[3]);
    nand g1278(n1491 ,n1209 ,n1162);
    nor g1279(n1704 ,n1102 ,n1585);
    or g1280(n1037 ,n1[15] ,n922);
    xnor g1281(n1575 ,n1115 ,n1116);
    or g1282(n249 ,n242 ,n230);
    nand g1283(n545 ,n474 ,n506);
    nor g1284(n789 ,n762 ,n0[6]);
    xnor g1285(n523 ,n425 ,n2040);
    xnor g1286(n940 ,n0[51] ,n0[50]);
    nor g1287(n1740 ,n968 ,n1609);
    nand g1288(n736 ,n2013 ,n2014);
    or g1289(n1512 ,n1[18] ,n1257);
    or g1290(n1468 ,n1047 ,n1237);
    nand g1291(n240 ,n214 ,n201);
    nor g1292(n1885 ,n990 ,n1877);
    nand g1293(n178 ,n116 ,n144);
    nand g1294(n456 ,n2063 ,n381);
    xnor g1295(n1125 ,n892 ,n883);
    nand g1296(n726 ,n723 ,n720);
    xnor g1297(n874 ,n0[43] ,n0[42]);
    or g1298(n296 ,n266 ,n282);
    nor g1299(n1156 ,n888 ,n1045);
    nand g1300(n1674 ,n1[24] ,n1553);
    nand g1301(n241 ,n213 ,n200);
    nand g1302(n1564 ,n1414 ,n1413);
    nand g1303(n1909 ,n4[1] ,n4[0]);
    or g1304(n393 ,n2095 ,n2073);
    or g1305(n1609 ,n969 ,n1490);
    xnor g1306(n1854 ,n1[13] ,n1793);
    xnor g1307(n904 ,n0[57] ,n0[41]);
    nand g1308(n1636 ,n1470 ,n1526);
    nand g1309(n1457 ,n1048 ,n1247);
    not g1310(n338 ,n337);
    xnor g1311(n6[46] ,n0[46] ,n1324);
    nand g1312(n549 ,n484 ,n509);
    nor g1313(n830 ,n773 ,n1[0]);
    nor g1314(n1876 ,n993 ,n1868);
    nand g1315(n712 ,n697 ,n707);
    nand g1316(n1393 ,n1993 ,n1106);
    nand g1317(n7[19] ,n1664 ,n1613);
    nor g1318(n1614 ,n1449 ,n1495);
    or g1319(n1472 ,n758 ,n1229);
    or g1320(n820 ,n756 ,n1984);
    nand g1321(n965 ,n826 ,n803);
    not g1322(n2071 ,n0[26]);
    nand g1323(n590 ,n542 ,n559);
    not g1324(n759 ,n0[4]);
    or g1325(n70 ,n0[56] ,n0[8]);
    nand g1326(n146 ,n77 ,n122);
    nand g1327(n1382 ,n997 ,n1092);
    nand g1328(n1363 ,n1002 ,n1079);
    xnor g1329(n158 ,n94 ,n115);
    nand g1330(n206 ,n154 ,n170);
    xnor g1331(n580 ,n525 ,n474);
    nand g1332(n372 ,n343 ,n366);
    nand g1333(n838 ,n5[4] ,n772);
    nor g1334(n304 ,n244 ,n285);
    not g1335(n738 ,n0[3]);
    nand g1336(n1265 ,n2027 ,n1053);
    not g1337(n2070 ,n0[27]);
    nand g1338(n1312 ,n2020 ,n1050);
    nand g1339(n322 ,n321 ,n312);
    nor g1340(n806 ,n742 ,n1993);
    nor g1341(n1955 ,n1946 ,n1945);
    nand g1342(n548 ,n476 ,n510);
    nand g1343(n1354 ,n0[6] ,n1105);
    nand g1344(n1322 ,n2024 ,n1051);
    not g1345(n348 ,n347);
    or g1346(n1002 ,n1[30] ,n896);
    nand g1347(n7[3] ,n1631 ,n1852);
    xnor g1348(n525 ,n467 ,n472);
    xnor g1349(n1121 ,n893 ,n888);
    nand g1350(n1647 ,n1507 ,n1406);
    xnor g1351(n555 ,n501 ,n519);
    nand g1352(n340 ,n327 ,n325);
    nor g1353(n1475 ,n1360 ,n1148);
    nand g1354(n1751 ,n1[15] ,n1583);
    or g1355(n995 ,n5[5] ,n842);
    or g1356(n535 ,n487 ,n489);
    not g1357(n739 ,n1[4]);
    nand g1358(n278 ,n234 ,n254);
    buf g1359(n12[2], 1'b0);
    nand g1360(n463 ,n2065 ,n391);
    nand g1361(n1547 ,n1392 ,n1197);
    nand g1362(n1202 ,n0[4] ,n1100);
    or g1363(n1438 ,n740 ,n1259);
    xnor g1364(n915 ,n0[28] ,n0[27]);
    xnor g1365(n32 ,n22 ,n27);
    nand g1366(n1038 ,n949 ,n951);
    nand g1367(n1673 ,n1397 ,n1434);
    xnor g1368(n629 ,n598 ,n600);
    xnor g1369(n425 ,n2080 ,n2081);
    xnor g1370(n265 ,n222 ,n168);
    xnor g1371(n855 ,n0[42] ,n0[18]);
    xnor g1372(n888 ,n0[25] ,n0[24]);
    nand g1373(n1943 ,n1920 ,n1918);
    nand g1374(n823 ,n2002 ,n753);
    nand g1375(n1199 ,n0[58] ,n1101);
    nor g1376(n787 ,n746 ,n0[5]);
    xnor g1377(n854 ,n0[33] ,n0[9]);
    not g1378(n2123 ,n2122);
    nand g1379(n1546 ,n1388 ,n1387);
    nor g1380(n2099 ,n1891 ,n1897);
    xnor g1381(n849 ,n0[36] ,n0[12]);
    nand g1382(n1948 ,n1935 ,n1930);
    nand g1383(n379 ,n324 ,n378);
    nand g1384(n84 ,n0[33] ,n0[9]);
    nand g1385(n290 ,n241 ,n272);
    xnor g1386(n335 ,n309 ,n289);
    not g1387(n882 ,n883);
    nand g1388(n953 ,n788 ,n796);
    xnor g1389(n1770 ,n1[2] ,n1586);
    nand g1390(n1666 ,n1[21] ,n1553);
    nand g1391(n1979 ,n2012 ,n1056);
    nand g1392(n1333 ,n0[19] ,n1100);
    nand g1393(n419 ,n2095 ,n2073);
    nand g1394(n1498 ,n1342 ,n1141);
    not g1395(n2089 ,n0[8]);
    nand g1396(n1327 ,n1033 ,n1075);
    nand g1397(n1083 ,n1[22] ,n892);
    nor g1398(n799 ,n743 ,n0[63]);
    xnor g1399(n245 ,n140 ,n202);
    xnor g1400(n1923 ,n0[16] ,n1[16]);
    xnor g1401(n219 ,n154 ,n172);
    nand g1402(n693 ,n674 ,n679);
    xnor g1403(n1120 ,n861 ,n864);
    nand g1404(n543 ,n499 ,n497);
    nand g1405(n154 ,n80 ,n133);
    xnor g1406(n1925 ,n0[6] ,n1[6]);
    xnor g1407(n2006 ,n1[6] ,n1576);
    xnor g1408(n1776 ,n1[11] ,n1569);
    xnor g1409(n6[8] ,n0[8] ,n1312);
    nand g1410(n1407 ,n1172 ,n1204);
    nor g1411(n1823 ,n1805 ,n1804);
    xnor g1412(n174 ,n0[47] ,n100);
    not g1413(n2035 ,n0[62]);
    nand g1414(n316 ,n260 ,n293);
    xnor g1415(n119 ,n0[35] ,n0[11]);
    nand g1416(n243 ,n175 ,n212);
    nand g1417(n968 ,n825 ,n816);
    or g1418(n1725 ,n1554 ,n1565);
    nand g1419(n1810 ,n1749 ,n1748);
    nor g1420(n1411 ,n1372 ,n1364);
    not g1421(n1232 ,n1231);
    nor g1422(n1684 ,n1593 ,n1591);
    nor g1423(n1046 ,n834 ,n989);
    nand g1424(n1809 ,n1700 ,n1735);
    not g1425(n334 ,n333);
    nand g1426(n640 ,n609 ,n621);
    xnor g1427(n165 ,n110 ,n0[33]);
    xnor g1428(n189 ,n153 ,n150);
    or g1429(n574 ,n568 ,n567);
    not g1430(n2081 ,n0[16]);
    not g1431(n899 ,n900);
    nand g1432(n484 ,n416 ,n448);
    not g1433(n2051 ,n0[46]);
    nand g1434(n841 ,n2028 ,n774);
    nand g1435(n561 ,n504 ,n530);
    nand g1436(n1307 ,n2024 ,n1109);
    not g1437(n746 ,n1[10]);
    nand g1438(n1501 ,n1337 ,n1185);
    xnor g1439(n1133 ,n1[9] ,n980);
    nand g1440(n151 ,n84 ,n129);
    xnor g1441(n6[27] ,n0[27] ,n1289);
    or g1442(n383 ,n2070 ,n2057);
    xnor g1443(n6[9] ,n0[9] ,n1313);
    or g1444(n1835 ,n2004 ,n2006);
    nand g1445(n88 ,n0[20] ,n0[4]);
    not g1446(n2041 ,n0[56]);
    nand g1447(n214 ,n88 ,n182);
    xnor g1448(n1225 ,n0[17] ,n904);
    nor g1449(n1967 ,n2098 ,n1982);
    not g1450(n985 ,n986);
    xor g1451(n1261 ,n0[63] ,n862);
    nor g1452(n949 ,n780 ,n778);
    or g1453(n605 ,n577 ,n584);
    nand g1454(n587 ,n522 ,n572);
    xnor g1455(n1988 ,n731 ,n702);
    nand g1456(n1675 ,n1[25] ,n1553);
    nand g1457(n318 ,n288 ,n295);
    or g1458(n60 ,n0[30] ,n0[14]);
    nand g1459(n451 ,n2056 ,n383);
    nand g1460(n1473 ,n758 ,n1229);
    nand g1461(n457 ,n2080 ,n386);
    xnor g1462(n6[40] ,n0[40] ,n1266);
    nand g1463(n332 ,n262 ,n320);
    or g1464(n7[1] ,n1718 ,n1850);
    xnor g1465(n704 ,n676 ,n685);
    nand g1466(n676 ,n652 ,n665);
    nor g1467(n1613 ,n1477 ,n1504);
    xnor g1468(n497 ,n430 ,n2044);
    nor g1469(n1841 ,n1800 ,n1821);
    nor g1470(n1105 ,n834 ,n993);
    or g1471(n1065 ,n763 ,n982);
    nor g1472(n1884 ,n2006 ,n1878);
    nand g1473(n2032 ,n735 ,n736);
    nand g1474(n272 ,n227 ,n258);
    nand g1475(n1269 ,n2023 ,n1053);
    xnor g1476(n247 ,n213 ,n200);
    nand g1477(n363 ,n355 ,n348);
    nand g1478(n2028 ,n4[0] ,n1908);
    nand g1479(n1902 ,n2019 ,n1898);
    nand g1480(n1525 ,n1[14] ,n1243);
    xnor g1481(n1929 ,n0[25] ,n1[25]);
    or g1482(n720 ,n705 ,n718);
    nor g1483(n1858 ,n1806 ,n1822);
    nand g1484(n355 ,n330 ,n335);
    not g1485(n2092 ,n0[5]);
    xnor g1486(n1774 ,n1[3] ,n1584);
    nor g1487(n1801 ,n1597 ,n1731);
    xnor g1488(n6[15] ,n0[15] ,n1319);
    nand g1489(n136 ,n0[39] ,n65);
    not g1490(n491 ,n490);
    nand g1491(n1592 ,n1445 ,n1478);
    or g1492(n1982 ,n3 ,n1977);
    nand g1493(n1323 ,n2023 ,n1051);
    nand g1494(n1364 ,n1032 ,n1081);
    or g1495(n1906 ,n1977 ,n2031);
    nor g1496(n271 ,n257 ,n250);
    nor g1497(n1050 ,n836 ,n995);
    xnor g1498(n1227 ,n766 ,n910);
    nor g1499(n1883 ,n1876 ,n1857);
    nand g1500(n342 ,n323 ,n312);
    xnor g1501(n1218 ,n0[47] ,n851);
    xnor g1502(n980 ,n0[5] ,n0[4]);
    xnor g1503(n6[7] ,n0[7] ,n1311);
    not g1504(n2080 ,n0[17]);
    or g1505(n386 ,n2040 ,n2081);
    nand g1506(n729 ,n728 ,n724);
    nand g1507(n1352 ,n0[20] ,n1100);
    nand g1508(n1981 ,n2032 ,n1400);
    xnor g1509(n1911 ,n0[11] ,n1[11]);
    nand g1510(n1084 ,n1[20] ,n900);
    nor g1511(n811 ,n758 ,n1983);
    xnor g1512(n711 ,n695 ,n701);
    nand g1513(n635 ,n571 ,n618);
    xnor g1514(n998 ,n0[1] ,n1[3]);
    nand g1515(n415 ,n2096 ,n2092);
    not g1516(n162 ,n161);
    nor g1517(n778 ,n741 ,n0[1]);
    nand g1518(n702 ,n642 ,n694);
    nand g1519(n1589 ,n1437 ,n1472);
    nand g1520(n1958 ,n1929 ,n1955);
    or g1521(n1892 ,n1982 ,n1889);
    nand g1522(n2125 ,n5[0] ,n2119);
    xnor g1523(n660 ,n628 ,n599);
    nand g1524(n470 ,n405 ,n453);
    nand g1525(n1494 ,n1354 ,n1160);
    nand g1526(n563 ,n501 ,n536);
    nand g1527(n607 ,n576 ,n578);
    xnor g1528(n6[35] ,n0[35] ,n1276);
    nand g1529(n360 ,n325 ,n349);
    nand g1530(n289 ,n239 ,n277);
    xnor g1531(n669 ,n646 ,n645);
    xnor g1532(n116 ,n0[57] ,n0[49]);
    nand g1533(n1534 ,n1211 ,n1350);
    nor g1534(n1485 ,n1[15] ,n1261);
    nand g1535(n1301 ,n2025 ,n1049);
    nand g1536(n1496 ,n1351 ,n1167);
    nand g1537(n1446 ,n756 ,n1232);
    or g1538(n385 ,n2086 ,n2050);
    not g1539(n164 ,n163);
    or g1540(n7[26] ,n1347 ,n1763);
    xnor g1541(n930 ,n0[28] ,n0[4]);
    nand g1542(n714 ,n693 ,n709);
    nand g1543(n1154 ,n899 ,n1046);
    nand g1544(n1880 ,n1829 ,n1874);
    xnor g1545(n866 ,n0[55] ,n0[54]);
    xnor g1546(n1224 ,n0[55] ,n850);
    or g1547(n1608 ,n1515 ,n1514);
    xnor g1548(n6[18] ,n0[18] ,n1298);
    nand g1549(n1945 ,n1922 ,n1921);
    xnor g1550(n1939 ,n0[9] ,n1[9]);
    nand g1551(n1203 ,n0[5] ,n1100);
    xnor g1552(n912 ,n0[20] ,n0[19]);
    nand g1553(n1332 ,n0[61] ,n1101);
    or g1554(n1714 ,n1535 ,n1622);
    nand g1555(n1731 ,n1639 ,n1617);
    xnor g1556(n1572 ,n1123 ,n1124);
    nand g1557(n572 ,n517 ,n550);
    nand g1558(n179 ,n117 ,n143);
    xnor g1559(n1113 ,n865 ,n939);
    xor g1560(n1931 ,n0[24] ,n1[24]);
    nor g1561(n1606 ,n1170 ,n1500);
    nor g1562(n1755 ,n1635 ,n1546);
    not g1563(n1045 ,n1046);
    nand g1564(n376 ,n354 ,n373);
    or g1565(n681 ,n654 ,n670);
    nor g1566(n1828 ,n1071 ,n1812);
    nand g1567(n946 ,n815 ,n817);
    xnor g1568(n1251 ,n941 ,n751);
    or g1569(n66 ,n0[29] ,n0[13]);
    nand g1570(n1761 ,n1383 ,n1616);
    or g1571(n1716 ,n1102 ,n1579);
    nor g1572(n1421 ,n1[6] ,n1240);
    xnor g1573(n1134 ,n1[13] ,n977);
    nand g1574(n1526 ,n1[21] ,n1237);
    not g1575(n1104 ,n1105);
    xor g1576(n2019 ,n28 ,n32);
    xor g1577(n1246 ,n0[59] ,n860);
    nand g1578(n1441 ,n739 ,n1244);
    nand g1579(n673 ,n595 ,n660);
    or g1580(n1752 ,n1628 ,n1533);
    nand g1581(n1844 ,n1803 ,n1596);
    xnor g1582(n878 ,n0[45] ,n0[29]);
    xnor g1583(n872 ,n0[48] ,n0[16]);
    xor g1584(n1235 ,n0[16] ,n905);
    xnor g1585(n171 ,n0[2] ,n102);
    nand g1586(n707 ,n689 ,n699);
    nand g1587(n366 ,n334 ,n365);
    or g1588(n1437 ,n755 ,n1252);
    nand g1589(n1096 ,n1[29] ,n920);
    nand g1590(n1442 ,n740 ,n1259);
    xnor g1591(n573 ,n477 ,n537);
    nand g1592(n1548 ,n1394 ,n1393);
    or g1593(n803 ,n756 ,n1991);
    nand g1594(n1480 ,n1[10] ,n1250);
    nand g1595(n1214 ,n1003 ,n1058);
    nand g1596(n1192 ,n0[3] ,n1100);
    nand g1597(n1309 ,n2026 ,n1109);
    nor g1598(n1803 ,n1544 ,n1752);
    or g1599(n7[27] ,n1169 ,n1769);
    or g1600(n532 ,n495 ,n494);
    nor g1601(n1825 ,n1776 ,n1809);
    nor g1602(n791 ,n760 ,n1[14]);
    nor g1603(n337 ,n313 ,n329);
    nor g1604(n1621 ,n1460 ,n1430);
    nand g1605(n7[16] ,n1669 ,n1624);
    nor g1606(n1635 ,n758 ,n1552);
    or g1607(n1597 ,n1534 ,n1538);
    nand g1608(n225 ,n171 ,n192);
    xor g1609(n1983 ,n678 ,n595);
    xnor g1610(n1584 ,n0[3] ,n1220);
    nor g1611(n1019 ,n1[13] ,n919);
    xnor g1612(n6[13] ,n0[13] ,n1317);
    nand g1613(n131 ,n0[53] ,n54);
    xnor g1614(n687 ,n669 ,n649);
    or g1615(n389 ,n2039 ,n2046);
    nand g1616(n692 ,n673 ,n680);
    xnor g1617(n1557 ,n1[0] ,n1249);
    nor g1618(n1970 ,n1966 ,n2033);
    or g1619(n1003 ,n1[8] ,n890);
    nand g1620(n1273 ,n2024 ,n1052);
    nand g1621(n639 ,n608 ,n623);
    nand g1622(n1396 ,n1987 ,n1054);
    nand g1623(n465 ,n2054 ,n399);
    nand g1624(n1005 ,n743 ,n987);
    nand g1625(n1957 ,n1913 ,n1953);
    nor g1626(n1611 ,n1401 ,n1435);
    not g1627(n896 ,n895);
    xnor g1628(n1126 ,n900 ,n887);
    nand g1629(n1543 ,n1391 ,n1151);
    not g1630(n305 ,n304);
    nand g1631(n1205 ,n1021 ,n1070);
    or g1632(n1185 ,n922 ,n1045);
    xnor g1633(n6[54] ,n0[54] ,n1264);
    xnor g1634(n495 ,n428 ,n2064);
    not g1635(n47 ,n46);
    xnor g1636(n6[0] ,n0[0] ,n1310);
    nand g1637(n1193 ,n0[1] ,n1100);
    xnor g1638(n860 ,n0[43] ,n0[19]);
    xnor g1639(n2003 ,n40 ,n29);
    nand g1640(n1742 ,n1462 ,n1610);
    or g1641(n380 ,n2069 ,n2059);
    nand g1642(n10 ,n1981 ,n1971);
    not g1643(n889 ,n890);
    nand g1644(n11 ,n990 ,n1111);
    nand g1645(n181 ,n71 ,n147);
    nand g1646(n1667 ,n1[22] ,n1553);
    nor g1647(n1467 ,n1047 ,n1231);
    nand g1648(n1326 ,n1005 ,n1077);
    not g1649(n1400 ,n1384);
    nor g1650(n197 ,n169 ,n165);
    xnor g1651(n934 ,n0[22] ,n0[2]);
    not g1652(n144 ,n143);
    nor g1653(n1408 ,n1373 ,n1362);
    not g1654(n842 ,n841);
    not g1655(n750 ,n0[13]);
    nor g1656(n1499 ,n1353 ,n1155);
    nor g1657(n1051 ,n836 ,n994);
    nand g1658(n1508 ,n1188 ,n1173);
    nor g1659(n2100 ,n997 ,n1055);
    nand g1660(n684 ,n659 ,n675);
    nand g1661(n512 ,n469 ,n483);
    nand g1662(n1144 ,n1027 ,n1057);
    nand g1663(n468 ,n407 ,n451);
    xnor g1664(n6[3] ,n0[3] ,n1306);
    nand g1665(n129 ,n0[41] ,n72);
    nand g1666(n1522 ,n1[8] ,n1233);
    nand g1667(n1077 ,n1[1] ,n996);
    nand g1668(n1747 ,n1[14] ,n1579);
    xnor g1669(n20 ,n2011 ,n2004);
    not g1670(n1384 ,n1056);
    nand g1671(n277 ,n238 ,n261);
    nand g1672(n1378 ,n1999 ,n1106);
    not g1673(n36 ,n35);
    or g1674(n346 ,n331 ,n339);
    nand g1675(n1816 ,n1656 ,n1713);
    xnor g1676(n253 ,n191 ,n145);
    nor g1677(n1515 ,n1[22] ,n1242);
    nor g1678(n1172 ,n1010 ,n1024);
    or g1679(n194 ,n139 ,n168);
    nor g1680(n1348 ,n764 ,n1099);
    nand g1681(n1759 ,n1645 ,n1464);
    nand g1682(n31 ,n16 ,n27);
    not g1683(n1055 ,n1056);
    nor g1684(n1861 ,n1836 ,n1837);
    xnor g1685(n1565 ,n1113 ,n1117);
    xnor g1686(n556 ,n523 ,n490);
    not g1687(n2043 ,n0[54]);
    nand g1688(n1197 ,n0[2] ,n1100);
    or g1689(n536 ,n518 ,n519);
    xnor g1690(n577 ,n529 ,n475);
    nand g1691(n1812 ,n962 ,n1740);
    xnor g1692(n283 ,n245 ,n243);
    nand g1693(n373 ,n346 ,n370);
    or g1694(n510 ,n481 ,n471);
    or g1695(n1022 ,n1[10] ,n894);
    nand g1696(n664 ,n653 ,n647);
    nor g1697(n805 ,n741 ,n1992);
    nor g1698(n1691 ,n1647 ,n1646);
    or g1699(n1703 ,n1[10] ,n1577);
    nand g1700(n1669 ,n1[16] ,n1553);
    not g1701(n748 ,n1[14]);
    nand g1702(n331 ,n302 ,n319);
    nand g1703(n1286 ,n2025 ,n1107);
    xnor g1704(n2013 ,n46 ,n49);
    nand g1705(n1150 ,n987 ,n1046);
    xnor g1706(n594 ,n553 ,n493);
    xnor g1707(n444 ,n2042 ,n2043);
    or g1708(n121 ,n95 ,n59);
    or g1709(n1873 ,n1779 ,n1866);
    nor g1710(n1414 ,n1135 ,n1176);
    not g1711(n2088 ,n0[9]);
    nand g1712(n23 ,n2004 ,n15);
    xnor g1713(n442 ,n2069 ,n2058);
    nand g1714(n133 ,n0[37] ,n66);
    nand g1715(n631 ,n601 ,n617);
    nand g1716(n1506 ,n0[0] ,n1139);
    nor g1717(n1039 ,n1[3] ,n984);
    xnor g1718(n231 ,n120 ,n188);
    nand g1719(n1391 ,n1992 ,n1106);
    nor g1720(n1339 ,n750 ,n1099);
    nand g1721(n341 ,n332 ,n324);
    not g1722(n1001 ,n964);
    nand g1723(n81 ,n0[23] ,n0[7]);
    nand g1724(n7[2] ,n1630 ,n1851);
    nand g1725(n1147 ,n977 ,n1046);
    nand g1726(n7[10] ,n1641 ,n1838);
    not g1727(n2049 ,n0[48]);
    xnor g1728(n1136 ,n1[25] ,n917);
    or g1729(n630 ,n600 ,n616);
    nor g1730(n347 ,n330 ,n335);
    nand g1731(n406 ,n2094 ,n2089);
    or g1732(n610 ,n580 ,n579);
    xnor g1733(n685 ,n667 ,n675);
    xnor g1734(n1222 ,n1[13] ,n877);
    nor g1735(n1454 ,n1047 ,n1254);
    or g1736(n325 ,n307 ,n314);
    nand g1737(n483 ,n418 ,n464);
    nor g1738(n1652 ,n965 ,n1425);
    nand g1739(n1487 ,n1[15] ,n1261);
    xnor g1740(n1118 ,n852 ,n853);
    nand g1741(n1663 ,n1436 ,n1517);
    xnor g1742(n326 ,n292 ,n283);
    nor g1743(n1023 ,n879 ,n877);
    nand g1744(n513 ,n480 ,n468);
    buf g1745(n13[5], 1'b0);
    xnor g1746(n575 ,n526 ,n484);
    xnor g1747(n905 ,n0[56] ,n0[40]);
    nand g1748(n45 ,n1975 ,n42);
    nand g1749(n1337 ,n0[15] ,n1100);
    nand g1750(n1158 ,n897 ,n1046);
    nand g1751(n653 ,n625 ,n635);
    nand g1752(n19 ,n2009 ,n2008);
    nand g1753(n229 ,n172 ,n193);
    nand g1754(n1297 ,n2027 ,n1052);
    or g1755(n1167 ,n916 ,n1045);
    xnor g1756(n6[60] ,n0[60] ,n1325);
    nor g1757(n1344 ,n751 ,n1099);
    xnor g1758(n633 ,n593 ,n570);
    nand g1759(n156 ,n82 ,n125);
    xnor g1760(n6[23] ,n0[23] ,n1303);
    nand g1761(n143 ,n76 ,n124);
    nand g1762(n416 ,n2084 ,n2035);
    nor g1763(n1138 ,n782 ,n1043);
    xnor g1764(n686 ,n668 ,n670);
    nand g1765(n1386 ,n837 ,n1056);
    nand g1766(n1728 ,n1499 ,n1655);
    nand g1767(n1387 ,n1990 ,n1106);
    nand g1768(n1318 ,n2026 ,n1050);
    nor g1769(n1616 ,n1451 ,n1482);
    xnor g1770(n1772 ,n1[10] ,n1567);
    or g1771(n1028 ,n973 ,n970);
    xnor g1772(n1917 ,n0[4] ,n1[4]);
    not g1773(n755 ,n1[5]);
    nand g1774(n43 ,n1973 ,n1974);
    xnor g1775(n1220 ,n0[51] ,n846);
    or g1776(n644 ,n611 ,n638);
    nor g1777(n1625 ,n1467 ,n1502);
    nand g1778(n1016 ,n956 ,n952);
    nand g1779(n2111 ,n2029 ,n5[1]);
    not g1780(n884 ,n885);
    nor g1781(n1824 ,n1773 ,n1808);
    nand g1782(n1474 ,n1361 ,n1143);
    not g1783(n2061 ,n0[36]);
    xnor g1784(n902 ,n0[25] ,n0[9]);
    xnor g1785(n1238 ,n0[51] ,n926);
    xnor g1786(n526 ,n469 ,n483);
    nor g1787(n1402 ,n1103 ,n1243);
    nand g1788(n1277 ,n2022 ,n1053);
    nand g1789(n701 ,n683 ,n691);
    nand g1790(n478 ,n413 ,n458);
    xnor g1791(n102 ,n0[26] ,n0[18]);
    not g1792(n2114 ,n2113);
    or g1793(n7[29] ,n1344 ,n1764);
    nand g1794(n1737 ,n1561 ,n1562);
    or g1795(n1029 ,n1[14] ,n967);
    or g1796(n54 ,n0[61] ,n0[45]);
    xnor g1797(n981 ,n0[6] ,n0[5]);
    nor g1798(n1700 ,n1660 ,n1563);
    nand g1799(n1081 ,n1[13] ,n919);
    xnor g1800(n498 ,n431 ,n2050);
    xnor g1801(n6[61] ,n0[61] ,n1290);
    nand g1802(n1497 ,n1349 ,n1171);
    not g1803(n1973 ,n2016);
    nand g1804(n1539 ,n1378 ,n1174);
    nand g1805(n1941 ,n1911 ,n1924);
    xnor g1806(n6[53] ,n0[53] ,n1267);
    nand g1807(n1365 ,n0[62] ,n1101);
    nand g1808(n993 ,n2[1] ,n840);
    xnor g1809(n1915 ,n0[7] ,n1[7]);
    nor g1810(n1619 ,n1454 ,n1497);
    nor g1811(n371 ,n359 ,n367);
    nand g1812(n1862 ,n1841 ,n1842);
    nand g1813(n1658 ,n1530 ,n1489);
    nand g1814(n180 ,n141 ,n142);
    xnor g1815(n578 ,n527 ,n476);
    xnor g1816(n21 ,n2010 ,n2006);
    nand g1817(n663 ,n646 ,n645);
    nand g1818(n1306 ,n2023 ,n1109);
    not g1819(n747 ,n0[6]);
    nor g1820(n2027 ,n2102 ,n2121);
    xnor g1821(n986 ,n757 ,n0[3]);
    xnor g1822(n167 ,n103 ,n0[31]);
    xnor g1823(n98 ,n0[36] ,n0[12]);
    nor g1824(n1008 ,n1[6] ,n978);
    nand g1825(n1524 ,n1193 ,n1359);
    nand g1826(n29 ,n26 ,n25);
    nand g1827(n2000 ,n332 ,n379);
    nor g1828(n1653 ,n2032 ,n1483);
    nand g1829(n1590 ,n1479 ,n1446);
    nand g1830(n2031 ,n1905 ,n1901);
    xnor g1831(n996 ,n0[2] ,n0[1]);
    nand g1832(n475 ,n419 ,n449);
    nor g1833(n1633 ,n755 ,n1552);
    nand g1834(n1553 ,n3 ,n11);
    xnor g1835(n1219 ,n0[43] ,n847);
    nand g1836(n564 ,n502 ,n535);
    nor g1837(n1721 ,n1103 ,n1570);
    nand g1838(n1665 ,n1[20] ,n1553);
    xnor g1839(n918 ,n0[12] ,n0[11]);
    xnor g1840(n1938 ,n0[8] ,n1[8]);
    nor g1841(n1595 ,n1215 ,n1501);
    nor g1842(n1897 ,n3 ,n1896);
    nand g1843(n139 ,n89 ,n127);
    xnor g1844(n893 ,n0[29] ,n0[28]);
    nand g1845(n1560 ,n1441 ,n1440);
    or g1846(n1787 ,n1521 ,n1742);
    nand g1847(n1368 ,n1066 ,n1078);
    xnor g1848(n2010 ,n1[2] ,n1573);
    or g1849(n1806 ,n1757 ,n1599);
    nor g1850(n1140 ,n978 ,n1104);
    nand g1851(n2116 ,n2101 ,n2105);
    xnor g1852(n935 ,n0[23] ,n0[3]);
    nor g1853(n1989 ,n702 ,n732);
    nand g1854(n1381 ,n1094 ,n1088);
    not g1855(n767 ,n0[10]);
    nor g1856(n1188 ,n1035 ,n1009);
    nand g1857(n1440 ,n1[2] ,n1236);
    or g1858(n1030 ,n1[23] ,n921);
    or g1859(n1463 ,n1047 ,n1246);
    nand g1860(n1748 ,n1[15] ,n1578);
    nand g1861(n344 ,n313 ,n329);
    nand g1862(n1550 ,n1203 ,n1398);
    nand g1863(n7[8] ,n1692 ,n1801);
    nand g1864(n559 ,n505 ,n533);
    xnor g1865(n230 ,n158 ,n156);
    nand g1866(n210 ,n169 ,n165);
    nand g1867(n1161 ,n889 ,n1046);
    nand g1868(n155 ,n90 ,n134);
    xnor g1869(n880 ,n0[12] ,n750);
    xnor g1870(n120 ,n0[24] ,n0[40]);
    nand g1871(n1620 ,n1458 ,n1424);
    nor g1872(n1734 ,n1648 ,n1598);
    nand g1873(n1401 ,n1145 ,n1153);
    nand g1874(n79 ,n0[22] ,n0[6]);
    xnor g1875(n927 ,n0[62] ,n0[14]);
    or g1876(n967 ,n1[15] ,n830);
    xnor g1877(n944 ,n1[3] ,n1986);
    nand g1878(n454 ,n2097 ,n395);
    not g1879(n2029 ,n1909);
    nand g1880(n307 ,n255 ,n286);
    nor g1881(n1412 ,n1144 ,n1214);
    nor g1882(n1968 ,n1966 ,n1977);
    nor g1883(n1340 ,n768 ,n1099);
    nor g1884(n1701 ,n1[7] ,n1570);
    xnor g1885(n858 ,n0[63] ,n0[62]);
    nand g1886(n1971 ,n1969 ,n1968);
    nor g1887(n2106 ,n2028 ,n5[0]);
    or g1888(n1174 ,n913 ,n1045);
    nor g1889(n1594 ,n1486 ,n1551);
    xnor g1890(n1922 ,n0[29] ,n1[29]);
    nand g1891(n1304 ,n2021 ,n1109);
    nand g1892(n728 ,n725 ,n721);
    nor g1893(n1857 ,n989 ,n1823);
    nand g1894(n1388 ,n1983 ,n1054);
    nand g1895(n351 ,n344 ,n338);
    or g1896(n72 ,n0[33] ,n0[9]);
    nand g1897(n211 ,n52 ,n188);
    nand g1898(n843 ,n2[0] ,n769);
    nand g1899(n829 ,n1989 ,n740);
    nor g1900(n1868 ,n1419 ,n1859);
    or g1901(n298 ,n267 ,n284);
    or g1902(n1871 ,n1864 ,n1863);
    xnor g1903(n1258 ,n765 ,n901);
    xnor g1904(n111 ,n0[22] ,n0[6]);
    nand g1905(n39 ,n36 ,n37);
    nor g1906(n1040 ,n1[21] ,n916);
    nand g1907(n1600 ,n1041 ,n1417);
    xnor g1908(n339 ,n310 ,n288);
    or g1909(n1032 ,n1[27] ,n915);
    nand g1910(n827 ,n2[1] ,n770);
    nand g1911(n480 ,n402 ,n457);
    xnor g1912(n914 ,n0[32] ,n0[31]);
    not g1913(n987 ,n988);
    not g1914(n745 ,n1[9]);
    xnor g1915(n852 ,n0[61] ,n0[60]);
    nand g1916(n479 ,n409 ,n461);
    xnor g1917(n163 ,n119 ,n0[27]);
    nand g1918(n1139 ,n1104 ,n1099);
    nand g1919(n1796 ,n1448 ,n1685);
    or g1920(n1011 ,n1[16] ,n887);
    nand g1921(n1194 ,n743 ,n1006);
    nor g1922(n1456 ,n1047 ,n1250);
    or g1923(n508 ,n482 ,n470);
    xnor g1924(n612 ,n579 ,n591);
    not g1925(n2054 ,n0[43]);
    nor g1926(n797 ,n740 ,n0[62]);
    nor g1927(n1173 ,n1015 ,n1039);
    nand g1928(n1893 ,n992 ,n1890);
    nand g1929(n300 ,n268 ,n281);
    nor g1930(n2026 ,n2022 ,n2126);
    not g1931(n773 ,n1990);
    xnor g1932(n862 ,n0[39] ,n0[15]);
    nand g1933(n7[22] ,n1667 ,n1618);
    nand g1934(n1089 ,n1[21] ,n916);
    xnor g1935(n851 ,n0[31] ,n0[15]);
    or g1936(n1183 ,n996 ,n1045);
    nand g1937(n1768 ,n1345 ,n1678);
    nor g1938(n1551 ,n1[10] ,n1250);
    nand g1939(n239 ,n215 ,n203);
    nand g1940(n737 ,n1837 ,n1867);
    nand g1941(n1314 ,n2022 ,n1050);
    or g1942(n651 ,n633 ,n637);
    xnor g1943(n1566 ,n936 ,n1119);
    nor g1944(n1872 ,n1835 ,n1861);
    or g1945(n1896 ,n2[0] ,n1895);
    nand g1946(n1268 ,n2027 ,n1108);
    nand g1947(n234 ,n140 ,n202);
    nor g1948(n1846 ,n1778 ,n1777);
    nand g1949(n1798 ,n1468 ,n1725);
    xnor g1950(n876 ,n0[61] ,n0[13]);
    nand g1951(n1750 ,n1[11] ,n1585);
    nand g1952(n1637 ,n1527 ,n1512);
    xnor g1953(n6[5] ,n0[5] ,n1308);
    nand g1954(n1820 ,n1744 ,n1746);
    xnor g1955(n443 ,n2096 ,n2065);
    or g1956(n1779 ,n1712 ,n1689);
    nand g1957(n276 ,n257 ,n250);
    nor g1958(n1170 ,n918 ,n1045);
    nand g1959(n1795 ,n1739 ,n1726);
    or g1960(n381 ,n2068 ,n2064);
    nor g1961(n1460 ,n1047 ,n1235);
    nand g1962(n626 ,n589 ,n604);
    or g1963(n466 ,n387 ,n444);
    nand g1964(n1536 ,n1399 ,n1332);
    xnor g1965(n200 ,n108 ,n148);
    nand g1966(n1516 ,n960 ,n1328);
    nand g1967(n1529 ,n1[19] ,n1246);
    nor g1968(n992 ,n2[2] ,n827);
    nor g1969(n1180 ,n919 ,n1045);
    nand g1970(n183 ,n55 ,n155);
    or g1971(n2124 ,n5[0] ,n2120);
    xnor g1972(n505 ,n424 ,n2066);
    nor g1973(n782 ,n761 ,n0[4]);
    nand g1974(n207 ,n151 ,n166);
    xnor g1975(n6[42] ,n0[42] ,n1262);
    xnor g1976(n292 ,n265 ,n260);
    or g1977(n1459 ,n1047 ,n1226);
    nand g1978(n1094 ,n1[28] ,n893);
    nand g1979(n1489 ,n1[12] ,n1239);
    xnor g1980(n6[55] ,n0[55] ,n1297);
    nand g1981(n1366 ,n1030 ,n1084);
    or g1982(n233 ,n140 ,n202);
    nand g1983(n1950 ,n1932 ,n1917);
    or g1984(n57 ,n0[48] ,n0[16]);
    nor g1985(n801 ,n755 ,n0[61]);
    not g1986(n1252 ,n1251);
    xnor g1987(n943 ,n0[57] ,n1[1]);
    nor g1988(n1708 ,n1560 ,n1638);
    or g1989(n1710 ,n1494 ,n1620);
    nand g1990(n417 ,n2091 ,n2037);
    not g1991(n1901 ,n2003);
    not g1992(n763 ,n1[11]);
    nand g1993(n1866 ,n1750 ,n1832);
    nor g1994(n1687 ,n1554 ,n1582);
    or g1995(n1429 ,n1103 ,n1240);
    nand g1996(n1274 ,n2024 ,n1108);
    not g1997(n2059 ,n0[38]);
    nand g1998(n1367 ,n1031 ,n1086);
    nand g1999(n1839 ,n1815 ,n1611);
    not g2000(n2076 ,n0[21]);
    nor g2001(n1699 ,n1557 ,n1558);
    nor g2002(n779 ,n754 ,n1[2]);
    nor g2003(n2015 ,n1951 ,n1964);
    nand g2004(n683 ,n654 ,n670);
    nor g2005(n1953 ,n1941 ,n1952);
    nand g2006(n1503 ,n1334 ,n1165);
    xnor g2007(n186 ,n0[43] ,n113);
    nand g2008(n294 ,n265 ,n283);
    xnor g2009(n6[51] ,n0[51] ,n1275);
    nand g2010(n731 ,n730 ,n723);
    xnor g2011(n504 ,n2091 ,n427);
    xnor g2012(n2008 ,n1[4] ,n1568);
    nand g2013(n1623 ,n1461 ,n1432);
    nor g2014(n1014 ,n1[0] ,n976);
    or g2015(n1448 ,n1047 ,n1242);
    nand g2016(n694 ,n664 ,n684);
    xnor g2017(n1562 ,n1[3] ,n1238);
    not g2018(n2042 ,n0[55]);
    xnor g2019(n551 ,n495 ,n494);
    xor g2020(n1991 ,n315 ,n252);
    nand g2021(n459 ,n2049 ,n385);
    nand g2022(n352 ,n328 ,n336);
    nand g2023(n260 ,n196 ,n232);
    xnor g2024(n6[25] ,n0[25] ,n1293);
    not g2025(n2068 ,n0[29]);
    xnor g2026(n1936 ,n0[27] ,n1[27]);
    nand g2027(n1518 ,n1062 ,n1181);
    xnor g2028(n595 ,n555 ,n518);
    not g2029(n353 ,n352);
    not g2030(n2078 ,n0[19]);
    nor g2031(n1106 ,n835 ,n991);
    nor g2032(n1720 ,n1103 ,n1577);
    nand g2033(n1651 ,n1416 ,n1415);
    nor g2034(n1739 ,n1672 ,n1608);
    nor g2035(n1686 ,n1103 ,n1583);
    xnor g2036(n557 ,n502 ,n487);
    xnor g2037(n519 ,n445 ,n2048);
    xnor g2038(n1574 ,n1129 ,n1121);
    nand g2039(n1145 ,n986 ,n1105);
    nand g2040(n1521 ,n1196 ,n1199);
    nand g2041(n796 ,n1[0] ,n766);
    xnor g2042(n172 ,n0[46] ,n114);
    nand g2043(n1549 ,n1396 ,n1202);
    xnor g2044(n6[47] ,n0[47] ,n1287);
    not g2045(n2058 ,n0[39]);
    nand g2046(n1447 ,n1048 ,n1238);
    nand g2047(n1357 ,n1037 ,n1060);
    xnor g2048(n2004 ,n1[7] ,n1582);
    nand g2049(n92 ,n0[26] ,n0[18]);
    xnor g2050(n6[34] ,n0[34] ,n1278);
    xnor g2051(n6[4] ,n0[4] ,n1307);
    nand g2052(n1338 ,n0[14] ,n1100);
    xnor g2053(n308 ,n266 ,n282);
    or g2054(n1601 ,n1540 ,n1476);
    xnor g2055(n173 ,n0[44] ,n99);
    nand g2056(n258 ,n206 ,n229);
    nand g2057(n476 ,n408 ,n455);
    xnor g2058(n487 ,n435 ,n2053);
    nand g2059(n132 ,n0[0] ,n70);
    or g2060(n398 ,n2071 ,n2053);
    nand g2061(n135 ,n0[34] ,n53);
    nor g2062(n819 ,n740 ,n1989);
    nand g2063(n1320 ,n2020 ,n1049);
    buf g2064(n13[7], 1'b0);
    xnor g2065(n923 ,n0[18] ,n0[17]);
    nand g2066(n140 ,n86 ,n121);
    nand g2067(n124 ,n0[32] ,n57);
    nand g2068(n636 ,n581 ,n619);
    nand g2069(n2122 ,n2118 ,n2116);
    or g2070(n721 ,n714 ,n715);
    nand g2071(n1281 ,n2020 ,n1108);
    nand g2072(n125 ,n0[25] ,n56);
    nor g2073(n1718 ,n1554 ,n1572);
    not g2074(n834 ,n833);
    or g2075(n1434 ,n1103 ,n1241);
    xnor g2076(n490 ,n443 ,n2092);
    or g2077(n1788 ,n1723 ,n1722);
    nand g2078(n1762 ,n1675 ,n1177);
    xnor g2079(n868 ,n0[50] ,n0[26]);
    nand g2080(n1090 ,n1[26] ,n898);
    xnor g2081(n895 ,n0[30] ,n768);
    nand g2082(n1650 ,n1431 ,n1412);
    xnor g2083(n908 ,n0[46] ,n0[30]);
    xnor g2084(n222 ,n139 ,n173);
    nand g2085(n1802 ,n1684 ,n1706);
    or g2086(n1881 ,n1982 ,n1872);
    nand g2087(n969 ,n832 ,n812);
    xnor g2088(n911 ,n0[48] ,n0[0]);
    xnor g2089(n6[28] ,n0[28] ,n1288);
    nand g2090(n1736 ,n1604 ,n1603);
    xnor g2091(n6[19] ,n0[19] ,n1299);
    nand g2092(n568 ,n514 ,n545);
    nand g2093(n674 ,n636 ,n662);
    xnor g2094(n424 ,n2083 ,n2067);
    nor g2095(n960 ,n804 ,n811);
    not g2096(n2056 ,n0[41]);
    or g2097(n1436 ,n879 ,n1222);
    nand g2098(n602 ,n570 ,n574);
    xnor g2099(n431 ,n2086 ,n2049);
    or g2100(n2025 ,n2115 ,n2114);
    xnor g2101(n1130 ,n903 ,n906);
    nand g2102(n1285 ,n2020 ,n1052);
    xnor g2103(n910 ,n0[32] ,n0[8]);
    buf g2104(n13[4], 1'b0);
    or g2105(n1464 ,n1047 ,n1261);
    nand g2106(n1102 ,n833 ,n992);
    not g2107(n1900 ,n2018);
    nor g2108(n1875 ,n1771 ,n1873);
    xnor g2109(n112 ,n0[25] ,n0[17]);
    nor g2110(n956 ,n797 ,n785);
    xnor g2111(n1221 ,n0[42] ,n859);
    xnor g2112(n1253 ,n0[55] ,n942);
    nand g2113(n1383 ,n1997 ,n1106);
    or g2114(n1554 ,n769 ,n1977);
    xor g2115(n285 ,n220 ,n253);
    nand g2116(n76 ,n0[48] ,n0[16]);
    nand g2117(n1308 ,n2025 ,n1109);
    nand g2118(n1142 ,n975 ,n1105);
    nand g2119(n623 ,n586 ,n605);
    xnor g2120(n48 ,n1974 ,n44);
    xnor g2121(n6[56] ,n0[56] ,n1292);
    xnor g2122(n1216 ,n0[53] ,n863);
    xnor g2123(n537 ,n422 ,n473);
    nand g2124(n521 ,n423 ,n473);
    not g2125(n2065 ,n0[32]);
    nand g2126(n350 ,n343 ,n334);
    nand g2127(n1541 ,n1389 ,n1142);
    nand g2128(n655 ,n624 ,n630);
    not g2129(n1047 ,n1048);
    nor g2130(n2017 ,n29 ,n41);
    not g2131(n1230 ,n1229);
    nand g2132(n1063 ,n1[10] ,n894);
    nand g2133(n477 ,n415 ,n463);
    nand g2134(n467 ,n406 ,n452);
    nand g2135(n1972 ,n1970 ,n1967);
    xnor g2136(n1132 ,n1[7] ,n984);
    nor g2137(n364 ,n353 ,n358);
    nand g2138(n128 ,n0[38] ,n60);
    not g2139(n2075 ,n0[22]);
    nand g2140(n581 ,n531 ,n562);
    xnor g2141(n501 ,n436 ,n2055);
    nand g2142(n1043 ,n950 ,n948);
    xnor g2143(n873 ,n0[58] ,n0[10]);
    nand g2144(n259 ,n205 ,n226);
    nand g2145(n446 ,n2060 ,n394);
    not g2146(n2103 ,n5[1]);
    nand g2147(n546 ,n475 ,n511);
    nand g2148(n195 ,n164 ,n161);
    not g2149(n2037 ,n0[60]);
    nor g2150(n785 ,n742 ,n0[59]);
    nor g2151(n2023 ,n2117 ,n2112);
    xnor g2152(n6[14] ,n0[14] ,n1318);
    nand g2153(n34 ,n28 ,n32);
    xnor g2154(n281 ,n246 ,n261);
    nand g2155(n1542 ,n1390 ,n1183);
    nand g2156(n232 ,n216 ,n195);
    nor g2157(n1159 ,n893 ,n1045);
    or g2158(n377 ,n337 ,n375);
    nor g2159(n1098 ,n1[4] ,n999);
    nand g2160(n675 ,n650 ,n666);
    or g2161(n1432 ,n1103 ,n1234);
    nor g2162(n12[5] ,n1982 ,n1867);
    not g2163(n588 ,n587);
    buf g2164(n13[6], 1'b0);
    xnor g2165(n1984 ,n708 ,n692);
    nand g2166(n1263 ,n2021 ,n1051);
    nand g2167(n1092 ,n2015 ,n971);
    nand g2168(n95 ,n0[58] ,n0[50]);
    xnor g2169(n1913 ,n0[12] ,n1[12]);
    xnor g2170(n552 ,n499 ,n497);
    nand g2171(n1213 ,n0[7] ,n1105);
    nand g2172(n7[14] ,n1716 ,n1799);
    nor g2173(n1877 ,n1795 ,n1870);
    nand g2174(n558 ,n500 ,n534);
    nand g2175(n716 ,n710 ,n711);
    or g2176(n7[15] ,n1759 ,n1843);
    nor g2177(n1010 ,n1[22] ,n892);
    xnor g2178(n932 ,n0[20] ,n0[4]);
    nand g2179(n90 ,n0[60] ,n0[44]);
    or g2180(n62 ,n0[62] ,n0[46]);
    nand g2181(n1538 ,n1376 ,n1161);
    nor g2182(n1404 ,n1103 ,n1249);
    nand g2183(n1523 ,n1[9] ,n1234);
    nand g2184(n562 ,n523 ,n538);
    not g2185(n752 ,n0[26]);
    xnor g2186(n218 ,n157 ,n159);
    xnor g2187(n596 ,n557 ,n489);
    or g2188(n1754 ,n1633 ,n1550);
    nand g2189(n1732 ,n1594 ,n1605);
    nand g2190(n567 ,n515 ,n548);
    xnor g2191(n6[63] ,n0[63] ,n1265);
    or g2192(n388 ,n2093 ,n2048);
    not g2193(n2063 ,n0[34]);
    or g2194(n1692 ,n1102 ,n1566);
    nand g2195(n994 ,n5[5] ,n841);
    nor g2196(n1453 ,n1047 ,n1258);
    buf g2197(n12[1], 1'b0);
    nand g2198(n1849 ,n1606 ,n1783);
    nor g2199(n1072 ,n958 ,n974);
    nand g2200(n1079 ,n1[11] ,n918);
    nand g2201(n262 ,n180 ,n236);
    xnor g2202(n97 ,n0[61] ,n0[53]);
    nand g2203(n1807 ,n1418 ,n1694);
    or g2204(n507 ,n479 ,n478);
    xnor g2205(n6[39] ,n0[39] ,n1268);
    nand g2206(n1336 ,n0[11] ,n1100);
    or g2207(n1033 ,n1[11] ,n918);
    nand g2208(n1670 ,n1[17] ,n1553);
    not g2209(n2039 ,n0[58]);
    nor g2210(n1514 ,n1[16] ,n1235);
    xnor g2211(n576 ,n528 ,n479);
    nand g2212(n1196 ,n0[1] ,n1105);
    xnor g2213(n2009 ,n1[3] ,n1574);
    xnor g2214(n524 ,n482 ,n470);
    xnor g2215(n906 ,n0[44] ,n0[20]);
    xnor g2216(n6[45] ,n0[45] ,n1295);
    nor g2217(n2115 ,n5[2] ,n2111);
    not g2218(n2055 ,n0[42]);
    xnor g2219(n1234 ,n904 ,n902);
    nand g2220(n1978 ,n2013 ,n1056);
    nor g2221(n795 ,n766 ,n1[0]);
    nand g2222(n1275 ,n2023 ,n1052);
    nand g2223(n1960 ,n1937 ,n1956);
    nand g2224(n1743 ,n1463 ,n1654);
    or g2225(n1777 ,n1686 ,n1687);
    nor g2226(n2002 ,n1942 ,n1961);
endmodule
