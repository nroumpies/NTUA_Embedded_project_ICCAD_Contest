module top (n0, n1, n2, n3, n4, n5, n6, n7, n8);
    input n0, n1, n2;
    input [11:0] n3, n4;
    input [2:0] n5;
    output n6, n7;
    output [11:0] n8;
    wire n0, n1, n2;
    wire [11:0] n3, n4;
    wire [2:0] n5;
    wire n6, n7;
    wire [11:0] n8;
    wire [11:0] n9;
    wire [11:0] n10;
    wire [2:0] n11;
    wire [11:0] n12;
    wire [19:0] n13;
    wire [18:0] n14;
    wire [12:0] n15;
    wire [12:0] n16;
    wire [12:0] n17;
    wire [12:0] n18;
    wire [3:0] n19;
    wire n20, n21, n22, n23, n24, n25, n26, n27;
    wire n28, n29, n30, n31, n32, n33, n34, n35;
    wire n36, n37, n38, n39, n40, n41, n42, n43;
    wire n44, n45, n46, n47, n48, n49, n50, n51;
    wire n52, n53, n54, n55, n56, n57, n58, n59;
    wire n60, n61, n62, n63, n64, n65, n66, n67;
    wire n68, n69, n70, n71, n72, n73, n74, n75;
    wire n76, n77, n78, n79, n80, n81, n82, n83;
    wire n84, n85, n86, n87, n88, n89, n90, n91;
    wire n92, n93, n94, n95, n96, n97, n98, n99;
    wire n100, n101, n102, n103, n104, n105, n106, n107;
    wire n108, n109, n110, n111, n112, n113, n114, n115;
    wire n116, n117, n118, n119, n120, n121, n122, n123;
    wire n124, n125, n126, n127, n128, n129, n130, n131;
    wire n132, n133, n134, n135, n136, n137, n138, n139;
    wire n140, n141, n142, n143, n144, n145, n146, n147;
    wire n148, n149, n150, n151, n152, n153, n154, n155;
    wire n156, n157, n158, n159, n160, n161, n162, n163;
    wire n164, n165, n166, n167, n168, n169, n170, n171;
    wire n172, n173, n174, n175, n176, n177, n178, n179;
    wire n180, n181, n182, n183, n184, n185, n186, n187;
    wire n188, n189, n190, n191, n192, n193, n194, n195;
    wire n196, n197, n198, n199, n200, n201, n202, n203;
    wire n204, n205, n206, n207, n208, n209, n210, n211;
    wire n212, n213, n214, n215, n216, n217, n218, n219;
    wire n220, n221, n222, n223, n224, n225, n226, n227;
    wire n228, n229, n230, n231, n232, n233, n234, n235;
    wire n236, n237, n238, n239, n240, n241, n242, n243;
    wire n244, n245, n246, n247, n248, n249, n250, n251;
    wire n252, n253, n254, n255, n256, n257, n258, n259;
    wire n260, n261, n262, n263, n264, n265, n266, n267;
    wire n268, n269, n270, n271, n272, n273, n274, n275;
    wire n276, n277, n278, n279, n280, n281, n282, n283;
    wire n284, n285, n286, n287, n288, n289, n290, n291;
    wire n292, n293, n294, n295, n296, n297, n298, n299;
    wire n300, n301, n302, n303, n304, n305, n306, n307;
    wire n308, n309, n310, n311, n312, n313, n314, n315;
    wire n316, n317, n318, n319, n320, n321, n322, n323;
    wire n324, n325, n326, n327, n328, n329, n330, n331;
    wire n332, n333, n334, n335, n336, n337, n338, n339;
    wire n340, n341, n342, n343, n344, n345, n346, n347;
    wire n348, n349, n350, n351, n352, n353, n354, n355;
    wire n356, n357, n358, n359, n360, n361, n362, n363;
    wire n364, n365, n366, n367, n368, n369, n370, n371;
    wire n372, n373, n374, n375, n376, n377, n378, n379;
    wire n380, n381, n382, n383, n384, n385, n386, n387;
    wire n388, n389, n390, n391, n392, n393, n394, n395;
    wire n396, n397, n398, n399, n400, n401, n402, n403;
    wire n404, n405, n406, n407, n408, n409, n410, n411;
    wire n412, n413, n414, n415, n416, n417, n418, n419;
    wire n420, n421, n422, n423, n424, n425, n426, n427;
    wire n428, n429, n430, n431, n432, n433, n434, n435;
    wire n436, n437, n438, n439, n440, n441, n442, n443;
    wire n444, n445, n446, n447, n448, n449, n450, n451;
    wire n452, n453, n454, n455, n456, n457, n458, n459;
    wire n460, n461, n462, n463, n464, n465, n466, n467;
    wire n468, n469, n470, n471, n472, n473, n474, n475;
    wire n476, n477, n478, n479, n480, n481, n482, n483;
    wire n484, n485, n486, n487, n488, n489, n490, n491;
    wire n492, n493, n494, n495, n496, n497, n498, n499;
    wire n500, n501, n502, n503, n504, n505, n506, n507;
    wire n508, n509, n510, n511, n512, n513, n514, n515;
    wire n516, n517, n518, n519, n520, n521, n522, n523;
    wire n524, n525, n526, n527, n528, n529, n530, n531;
    wire n532, n533, n534, n535, n536, n537, n538, n539;
    wire n540, n541, n542, n543, n544, n545, n546, n547;
    wire n548, n549, n550, n551, n552, n553, n554, n555;
    wire n556, n557, n558, n559, n560, n561, n562, n563;
    wire n564, n565, n566, n567, n568, n569, n570, n571;
    wire n572, n573, n574, n575, n576, n577, n578, n579;
    wire n580, n581, n582, n583, n584, n585, n586, n587;
    wire n588, n589, n590, n591, n592, n593, n594, n595;
    wire n596, n597, n598, n599, n600, n601, n602, n603;
    wire n604, n605, n606, n607, n608, n609, n610, n611;
    wire n612, n613, n614, n615, n616, n617, n618, n619;
    wire n620, n621, n622, n623, n624, n625, n626, n627;
    wire n628, n629, n630, n631, n632, n633, n634, n635;
    wire n636, n637, n638, n639, n640, n641, n642, n643;
    wire n644, n645, n646, n647, n648, n649, n650, n651;
    wire n652, n653, n654, n655, n656, n657, n658, n659;
    wire n660, n661, n662, n663, n664, n665, n666, n667;
    wire n668, n669, n670, n671, n672, n673, n674, n675;
    wire n676, n677, n678, n679, n680, n681, n682, n683;
    wire n684, n685, n686, n687, n688, n689, n690, n691;
    wire n692, n693, n694, n695, n696, n697, n698, n699;
    wire n700, n701, n702, n703, n704, n705, n706, n707;
    wire n708, n709, n710, n711, n712, n713, n714, n715;
    wire n716, n717, n718, n719, n720, n721, n722, n723;
    wire n724, n725, n726, n727, n728, n729, n730, n731;
    wire n732, n733, n734, n735, n736, n737, n738, n739;
    wire n740, n741, n742, n743, n744, n745, n746, n747;
    wire n748, n749, n750, n751, n752, n753, n754, n755;
    wire n756, n757, n758, n759, n760, n761, n762, n763;
    wire n764, n765, n766, n767, n768, n769, n770, n771;
    wire n772, n773, n774, n775, n776, n777, n778, n779;
    wire n780, n781, n782, n783, n784, n785, n786, n787;
    wire n788, n789, n790, n791, n792, n793, n794, n795;
    wire n796, n797, n798, n799, n800, n801, n802, n803;
    wire n804, n805, n806, n807, n808, n809, n810, n811;
    wire n812, n813, n814, n815, n816, n817, n818, n819;
    wire n820, n821, n822, n823, n824, n825, n826, n827;
    wire n828, n829, n830, n831, n832, n833, n834, n835;
    wire n836, n837, n838, n839, n840, n841, n842, n843;
    wire n844, n845, n846, n847, n848, n849, n850, n851;
    wire n852, n853, n854, n855, n856, n857, n858, n859;
    wire n860, n861, n862, n863, n864, n865, n866, n867;
    wire n868, n869, n870, n871, n872, n873, n874, n875;
    wire n876, n877, n878, n879, n880, n881, n882, n883;
    wire n884, n885, n886, n887, n888, n889, n890, n891;
    wire n892, n893, n894, n895, n896, n897, n898, n899;
    wire n900, n901, n902, n903, n904, n905, n906, n907;
    wire n908, n909, n910, n911, n912, n913, n914, n915;
    wire n916, n917, n918, n919, n920, n921, n922, n923;
    wire n924, n925, n926, n927, n928, n929, n930, n931;
    wire n932, n933, n934, n935, n936, n937, n938, n939;
    wire n940, n941, n942, n943, n944, n945, n946, n947;
    wire n948, n949, n950, n951, n952, n953, n954, n955;
    wire n956, n957, n958, n959, n960, n961, n962, n963;
    wire n964, n965, n966, n967, n968, n969, n970, n971;
    wire n972, n973, n974, n975, n976, n977, n978, n979;
    wire n980, n981, n982, n983, n984, n985, n986, n987;
    wire n988, n989, n990, n991, n992, n993, n994, n995;
    wire n996, n997, n998, n999, n1000, n1001, n1002, n1003;
    wire n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011;
    wire n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
    wire n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
    wire n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
    wire n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
    wire n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051;
    wire n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059;
    wire n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067;
    wire n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075;
    wire n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083;
    wire n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091;
    wire n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099;
    wire n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107;
    wire n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115;
    wire n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123;
    wire n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131;
    wire n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139;
    wire n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147;
    wire n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155;
    wire n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163;
    wire n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171;
    wire n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179;
    wire n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187;
    wire n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195;
    wire n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203;
    wire n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
    wire n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219;
    wire n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227;
    wire n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235;
    wire n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243;
    wire n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251;
    wire n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259;
    wire n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267;
    wire n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275;
    wire n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;
    wire n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291;
    wire n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;
    wire n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307;
    wire n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315;
    wire n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323;
    wire n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331;
    wire n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;
    wire n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;
    wire n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;
    wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
    wire n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;
    wire n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;
    wire n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387;
    wire n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395;
    wire n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403;
    wire n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411;
    wire n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419;
    wire n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427;
    wire n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435;
    wire n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443;
    wire n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451;
    wire n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459;
    wire n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467;
    wire n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475;
    wire n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483;
    wire n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491;
    wire n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499;
    wire n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507;
    wire n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515;
    wire n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523;
    wire n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531;
    wire n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539;
    wire n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547;
    wire n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555;
    wire n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563;
    wire n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571;
    wire n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579;
    wire n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587;
    wire n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595;
    wire n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603;
    wire n1604, n1605;
    nor g0(n270 ,n70 ,n164);
    xnor g1(n49 ,n30 ,n10[2]);
    xnor g2(n574 ,n474 ,n512);
    xnor g3(n66 ,n10[3] ,n9[8]);
    nand g4(n1268 ,n1176 ,n1132);
    nor g5(n280 ,n45 ,n214);
    nand g6(n169 ,n23 ,n52);
    xnor g7(n478 ,n366 ,n351);
    not g8(n928 ,n1440);
    xnor g9(n1489 ,n868 ,n894);
    nand g10(n1163 ,n1514 ,n1093);
    not g11(n1095 ,n1094);
    dff g12(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[5]), .Q(n10[5]));
    nor g13(n282 ,n129 ,n165);
    nor g14(n269 ,n119 ,n162);
    nor g15(n703 ,n590 ,n686);
    nor g16(n252 ,n78 ,n162);
    xnor g17(n764 ,n740 ,n721);
    not g18(n1087 ,n1072);
    nand g19(n1443 ,n1427 ,n1400);
    buf g20(n10[11] ,n1388);
    nor g21(n224 ,n75 ,n162);
    nor g22(n388 ,n167 ,n363);
    or g23(n729 ,n680 ,n722);
    not g24(n1390 ,n10[11]);
    or g25(n492 ,n324 ,n442);
    nor g26(n1036 ,n13[15] ,n13[14]);
    dff g27(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[4]), .Q(n9[4]));
    nor g28(n1305 ,n1028 ,n1215);
    nand g29(n737 ,n689 ,n714);
    xnor g30(n651 ,n531 ,n616);
    nand g31(n1175 ,n1494 ,n1095);
    nand g32(n987 ,n981 ,n986);
    nand g33(n1243 ,n1438 ,n1153);
    nand g34(n1426 ,n1474 ,n9[11]);
    nor g35(n523 ,n416 ,n483);
    nand g36(n1231 ,n1464 ,n1200);
    nand g37(n1221 ,n1484 ,n1152);
    nor g38(n898 ,n861 ,n897);
    nor g39(n1114 ,n1101 ,n1089);
    xnor g40(n453 ,n353 ,n370);
    nand g41(n1110 ,n1064 ,n1102);
    nor g42(n1297 ,n1269 ,n1268);
    xnor g43(n59 ,n24 ,n9[11]);
    nand g44(n1324 ,n1140 ,n1233);
    xnor g45(n702 ,n659 ,n632);
    nand g46(n1235 ,n1461 ,n1200);
    nor g47(n1340 ,n1274 ,n1322);
    buf g48(n913 ,n912);
    nand g49(n1394 ,n1452 ,n1391);
    nor g50(n944 ,n924 ,n1469);
    dff g51(.RN(n1), .SN(1'b1), .CK(n0), .D(n2), .Q(n1605));
    nand g52(n1395 ,n10[6] ,n1393);
    xnor g53(n623 ,n300 ,n570);
    not g54(n440 ,n422);
    xnor g55(n622 ,n509 ,n564);
    xnor g56(n624 ,n543 ,n510);
    not g57(n917 ,n1444);
    nand g58(n1135 ,n1510 ,n1103);
    nand g59(n610 ,n334 ,n572);
    xnor g60(n457 ,n349 ,n357);
    xnor g61(n878 ,n1516 ,n12[2]);
    nand g62(n1184 ,n1520 ,n1093);
    nor g63(n1116 ,n1027 ,n1099);
    nor g64(n331 ,n202 ,n237);
    not g65(n1152 ,n1151);
    not g66(n981 ,n9[3]);
    xnor g67(n131 ,n10[7] ,n9[10]);
    nand g68(n1542 ,n10[6] ,n1533);
    nand g69(n1459 ,n1418 ,n1396);
    not g70(n995 ,n10[0]);
    or g71(n806 ,n9[1] ,n10[1]);
    nor g72(n355 ,n179 ,n238);
    nand g73(n211 ,n33 ,n94);
    or g74(n943 ,n920 ,n1437);
    nand g75(n888 ,n863 ,n887);
    nand g76(n1401 ,n9[4] ,n1392);
    nor g77(n950 ,n930 ,n1445);
    nand g78(n1047 ,n10[2] ,n1019);
    nand g79(n1081 ,n12[8] ,n1012);
    nand g80(n432 ,n304 ,n318);
    xnor g81(n1558 ,n9[5] ,n10[5]);
    nor g82(n264 ,n112 ,n162);
    nor g83(n884 ,n860 ,n883);
    nor g84(n1209 ,n1067 ,n1111);
    nand g85(n1160 ,n1524 ,n1093);
    nor g86(n1118 ,n13[11] ,n1097);
    nand g87(n1132 ,n9[7] ,n1096);
    nor g88(n354 ,n171 ,n281);
    nand g89(n423 ,n170 ,n369);
    not g90(n932 ,n1464);
    nor g91(n599 ,n298 ,n537);
    xnor g92(n827 ,n9[1] ,n10[1]);
    not g93(n352 ,n351);
    not g94(n800 ,n799);
    nand g95(n645 ,n563 ,n592);
    nor g96(n256 ,n68 ,n164);
    nand g97(n294 ,n24 ,n211);
    nand g98(n774 ,n707 ,n773);
    not g99(n684 ,n683);
    nor g100(n400 ,n28 ,n296);
    nand g101(n1375 ,n1046 ,n1361);
    nand g102(n833 ,n814 ,n828);
    nor g103(n152 ,n62 ,n102);
    not g104(n1021 ,n9[7]);
    nor g105(n363 ,n142 ,n220);
    nand g106(n665 ,n603 ,n635);
    xor g107(n1506 ,n815 ,n836);
    or g108(n754 ,n721 ,n740);
    nor g109(n1067 ,n1026 ,n10[5]);
    nor g110(n1003 ,n10[2] ,n1002);
    nand g111(n1196 ,n1517 ,n1093);
    nor g112(n276 ,n123 ,n165);
    nand g113(n1178 ,n1521 ,n1093);
    nor g114(n933 ,n925 ,n1465);
    xnor g115(n74 ,n10[5] ,n9[8]);
    nor g116(n149 ,n61 ,n102);
    dff g117(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[10]), .Q(n9[10]));
    xnor g118(n879 ,n1518 ,n12[4]);
    nor g119(n1085 ,n1024 ,n10[3]);
    nand g120(n771 ,n712 ,n770);
    nor g121(n158 ,n63 ,n102);
    nor g122(n184 ,n114 ,n51);
    nor g123(n957 ,n10[0] ,n956);
    xnor g124(n57 ,n24 ,n9[2]);
    nor g125(n893 ,n869 ,n892);
    xnor g126(n820 ,n9[11] ,n802);
    nand g127(n844 ,n826 ,n843);
    nor g128(n1372 ,n1210 ,n1358);
    xnor g129(n473 ,n310 ,n347);
    nand g130(n18[12] ,n1544 ,n1583);
    nand g131(n1279 ,n1441 ,n1153);
    not g132(n1025 ,n9[10]);
    nor g133(n1336 ,n1254 ,n1318);
    or g134(n666 ,n613 ,n633);
    nand g135(n1167 ,n1515 ,n1093);
    nand g136(n1072 ,n13[17] ,n13[16]);
    nor g137(n522 ,n410 ,n490);
    nand g138(n1288 ,n1197 ,n1196);
    nand g139(n39 ,n23 ,n10[10]);
    nor g140(n247 ,n66 ,n215);
    not g141(n1012 ,n1605);
    or g142(n690 ,n589 ,n670);
    or g143(n384 ,n368 ,n302);
    nor g144(n343 ,n196 ,n254);
    xnor g145(n1501 ,n1578 ,n1557);
    nand g146(n562 ,n480 ,n526);
    nand g147(n1422 ,n1472 ,n9[11]);
    nand g148(n1312 ,n1068 ,n1221);
    nor g149(n584 ,n436 ,n542);
    nor g150(n344 ,n150 ,n282);
    nand g151(n956 ,n952 ,n9[0]);
    xnor g152(n592 ,n468 ,n514);
    nor g153(n691 ,n674 ,n642);
    dff g154(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[10]), .Q(n10[10]));
    nand g155(n1245 ,n1147 ,n1123);
    xnor g156(n1509 ,n825 ,n843);
    nor g157(n507 ,n345 ,n502);
    nand g158(n1543 ,n10[3] ,n1536);
    xnor g159(n116 ,n10[3] ,n9[2]);
    xnor g160(n58 ,n24 ,n9[9]);
    nor g161(n843 ,n803 ,n842);
    nand g162(n508 ,n417 ,n481);
    or g163(n496 ,n330 ,n449);
    nor g164(n301 ,n216 ,n243);
    nor g165(n362 ,n180 ,n263);
    xnor g166(n570 ,n478 ,n328);
    nor g167(n279 ,n131 ,n164);
    nand g168(n975 ,n953 ,n974);
    nor g169(n1051 ,n1018 ,n10[1]);
    nand g170(n1418 ,n1470 ,n9[11]);
    nand g171(n1044 ,n11[0] ,n11[1]);
    or g172(n395 ,n347 ,n310);
    nand g173(n1054 ,n10[9] ,n1017);
    nand g174(n1189 ,n1486 ,n1091);
    xnor g175(n876 ,n1523 ,n12[9]);
    xnor g176(n1600 ,n1599 ,n1591);
    nor g177(n730 ,n694 ,n711);
    not g178(n166 ,n167);
    nor g179(n1100 ,n11[2] ,n1030);
    xnor g180(n119 ,n10[9] ,n9[5]);
    xnor g181(n700 ,n655 ,n521);
    nand g182(n165 ,n93 ,n100);
    xnor g183(n64 ,n10[9] ,n9[10]);
    not g184(n656 ,n655);
    nor g185(n265 ,n113 ,n165);
    nand g186(n1417 ,n1480 ,n9[11]);
    nor g187(n904 ,n855 ,n901);
    nor g188(n954 ,n918 ,n1463);
    nor g189(n490 ,n371 ,n441);
    nand g190(n1220 ,n1485 ,n1152);
    nand g191(n1319 ,n1128 ,n1228);
    not g192(n915 ,n912);
    nor g193(n673 ,n580 ,n640);
    not g194(n620 ,n608);
    nand g195(n1123 ,n9[1] ,n1096);
    nor g196(n513 ,n381 ,n484);
    nor g197(n366 ,n182 ,n264);
    xnor g198(n471 ,n341 ,n308);
    nor g199(n934 ,n923 ,n1447);
    dff g200(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[11]), .Q(n9[11]));
    xnor g201(n762 ,n742 ,n746);
    nand g202(n1405 ,n10[2] ,n1393);
    not g203(n596 ,n579);
    nand g204(n1551 ,n10[9] ,n1534);
    xnor g205(n1476 ,n9[7] ,n990);
    not g206(n837 ,n836);
    xnor g207(n576 ,n525 ,n522);
    xor g208(n13[13] ,n910 ,n14[13]);
    not g209(n1392 ,n9[11]);
    not g210(n1391 ,n1390);
    nand g211(n619 ,n392 ,n561);
    nand g212(n1583 ,n1526 ,n1582);
    nand g213(n1468 ,n1416 ,n1414);
    nand g214(n435 ,n362 ,n341);
    xnor g215(n621 ,n545 ,n520);
    nand g216(n1574 ,n1542 ,n1573);
    nand g217(n1462 ,n1424 ,n1401);
    or g218(n1030 ,n11[0] ,n11[1]);
    nor g219(n1299 ,n1273 ,n1272);
    not g220(n1535 ,n9[1]);
    xnor g221(n90 ,n23 ,n10[7]);
    nand g222(n720 ,n671 ,n679);
    xnor g223(n708 ,n654 ,n674);
    or g224(n493 ,n376 ,n443);
    not g225(n711 ,n705);
    xnor g226(n80 ,n10[1] ,n9[6]);
    nand g227(n951 ,n1442 ,n932);
    nand g228(n775 ,n731 ,n774);
    nor g229(n642 ,n563 ,n592);
    xnor g230(n13[14] ,n912 ,n14[14]);
    nor g231(n263 ,n82 ,n214);
    nand g232(n213 ,n36 ,n92);
    nand g233(n1240 ,n1488 ,n1152);
    nor g234(n1104 ,n1014 ,n1043);
    nand g235(n1576 ,n1541 ,n1575);
    dff g236(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[7]), .Q(n10[7]));
    not g237(n1090 ,n1091);
    nand g238(n887 ,n880 ,n886);
    dff g239(.RN(n1), .SN(1'b1), .CK(n0), .D(n1313), .Q(n12[2]));
    nand g240(n1434 ,n1455 ,n1391);
    nor g241(n368 ,n192 ,n287);
    nand g242(n42 ,n23 ,n10[6]);
    nor g243(n1062 ,n1021 ,n10[7]);
    xnor g244(n52 ,n29 ,n10[6]);
    nor g245(n489 ,n373 ,n440);
    nand g246(n766 ,n748 ,n755);
    nor g247(n375 ,n194 ,n259);
    nand g248(n1150 ,n9[9] ,n1096);
    xnor g249(n1450 ,n10[3] ,n1003);
    not g250(n448 ,n433);
    nor g251(n187 ,n68 ,n53);
    nand g252(n1270 ,n1179 ,n1178);
    nand g253(n1257 ,n1164 ,n1150);
    dff g254(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[1]), .Q(n11[1]));
    nand g255(n1381 ,n1271 ,n1369);
    nor g256(n988 ,n9[4] ,n987);
    xor g257(n1470 ,n9[1] ,n979);
    xor g258(n470 ,n338 ,n354);
    nand g259(n1399 ,n9[3] ,n1392);
    nand g260(n1145 ,n1516 ,n1093);
    nor g261(n1338 ,n1264 ,n1320);
    nand g262(n863 ,n1518 ,n12[4]);
    nand g263(n1330 ,n1081 ,n1239);
    xnor g264(n84 ,n10[9] ,n9[3]);
    dff g265(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[3]), .Q(n9[3]));
    not g266(n856 ,n14[13]);
    nand g267(n1048 ,n12[4] ,n1012);
    nor g268(n192 ,n84 ,n51);
    not g269(n920 ,n1459);
    nor g270(n369 ,n186 ,n271);
    nor g271(n401 ,n166 ,n364);
    xnor g272(n108 ,n10[7] ,n9[1]);
    nor g273(n616 ,n413 ,n558);
    nor g274(n254 ,n57 ,n214);
    nand g275(n760 ,n666 ,n749);
    or g276(n941 ,n931 ,n1468);
    nand g277(n1409 ,n9[5] ,n1392);
    nor g278(n479 ,n321 ,n401);
    nand g279(n1261 ,n1171 ,n1129);
    xnor g280(n474 ,n292 ,n332);
    nor g281(n312 ,n177 ,n221);
    xnor g282(n533 ,n166 ,n467);
    nand g283(n1465 ,n1431 ,n1407);
    nand g284(n1216 ,n1389 ,n1200);
    nand g285(n427 ,n347 ,n310);
    not g286(n539 ,n538);
    xnor g287(n465 ,n168 ,n307);
    nand g288(n905 ,n902 ,n901);
    nor g289(n160 ,n129 ,n100);
    nand g290(n170 ,n23 ,n101);
    nor g291(n1031 ,n13[13] ,n13[12]);
    xnor g292(n63 ,n24 ,n9[7]);
    nor g293(n1295 ,n1256 ,n1257);
    or g294(n421 ,n337 ,n323);
    nor g295(n175 ,n59 ,n102);
    nand g296(n1445 ,n1425 ,n1403);
    nand g297(n1281 ,n1191 ,n1199);
    nand g298(n796 ,n644 ,n795);
    xor g299(n1505 ,n831 ,n834);
    xnor g300(n538 ,n455 ,n376);
    nand g301(n1064 ,n10[6] ,n1023);
    xnor g302(n699 ,n589 ,n670);
    nor g303(n852 ,n821 ,n851);
    nand g304(n1078 ,n14[12] ,n14[11]);
    xnor g305(n1557 ,n9[9] ,n10[9]);
    xnor g306(n15[11] ,n1582 ,n1526);
    nor g307(n188 ,n132 ,n100);
    nor g308(n733 ,n673 ,n719);
    nand g309(n781 ,n756 ,n780);
    nand g310(n953 ,n1468 ,n931);
    nor g311(n201 ,n32 ,n87);
    nor g312(n509 ,n403 ,n485);
    nor g313(n719 ,n593 ,n683);
    not g314(n823 ,n822);
    nand g315(n780 ,n758 ,n779);
    not g316(n649 ,n639);
    nor g317(n141 ,n115 ,n51);
    nand g318(n1317 ,n1226 ,n1290);
    nand g319(n608 ,n474 ,n532);
    xnor g320(n117 ,n10[3] ,n9[11]);
    xnor g321(n1483 ,n878 ,n882);
    nand g322(n782 ,n781 ,n757);
    nor g323(n1332 ,n1242 ,n1291);
    nand g324(n749 ,n638 ,n735);
    xnor g325(n458 ,n302 ,n368);
    nand g326(n1568 ,n1543 ,n1567);
    nand g327(n1566 ,n1550 ,n1565);
    nand g328(n43 ,n23 ,n10[2]);
    nor g329(n243 ,n128 ,n163);
    nand g330(n520 ,n395 ,n487);
    nand g331(n1134 ,n9[6] ,n1096);
    nand g332(n1247 ,n1175 ,n1144);
    xnor g333(n1484 ,n877 ,n884);
    nor g334(n315 ,n155 ,n224);
    nand g335(n1308 ,n1057 ,n1217);
    xnor g336(n459 ,n342 ,n343);
    xnor g337(n83 ,n10[3] ,n9[3]);
    xnor g338(n1502 ,n1580 ,n1556);
    dff g339(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[1]), .Q(n9[1]));
    nand g340(n1570 ,n1549 ,n1569);
    nor g341(n383 ,n174 ,n336);
    nand g342(n1406 ,n10[4] ,n1393);
    xnor g343(n679 ,n623 ,n528);
    nor g344(n407 ,n292 ,n332);
    nand g345(n1403 ,n10[9] ,n1393);
    nand g346(n606 ,n551 ,n568);
    xnor g347(n468 ,n298 ,n315);
    not g348(n1528 ,n1527);
    nor g349(n138 ,n71 ,n54);
    nor g350(n859 ,n1522 ,n12[8]);
    not g351(n923 ,n1469);
    nand g352(n1149 ,n1482 ,n1091);
    xnor g353(n1560 ,n9[1] ,n10[1]);
    xnor g354(n469 ,n166 ,n363);
    nand g355(n1593 ,n1525 ,n19[0]);
    or g356(n390 ,n313 ,n314);
    nand g357(n1265 ,n1444 ,n1153);
    nor g358(n1204 ,n1045 ,n1106);
    nor g359(n960 ,n939 ,n959);
    dff g360(.RN(n1), .SN(1'b1), .CK(n0), .D(n1386), .Q(n8[8]));
    xnor g361(n725 ,n590 ,n686);
    xnor g362(n577 ,n339 ,n508);
    xnor g363(n107 ,n10[5] ,n9[11]);
    nand g364(n1376 ,n1243 ,n1364);
    xnor g365(n768 ,n755 ,n748);
    nor g366(n671 ,n601 ,n649);
    nand g367(n808 ,n9[8] ,n10[8]);
    nand g368(n993 ,n982 ,n992);
    not g369(n31 ,n23);
    nand g370(n1129 ,n9[8] ,n1096);
    dff g371(.RN(n1), .SN(1'b1), .CK(n0), .D(n1382), .Q(n8[6]));
    nand g372(n429 ,n343 ,n342);
    not g373(n1534 ,n9[9]);
    nor g374(n694 ,n521 ,n656);
    nor g375(n284 ,n120 ,n163);
    xor g376(n21 ,n568 ,n515);
    nor g377(n1053 ,n1025 ,n10[10]);
    or g378(n491 ,n325 ,n447);
    nand g379(n1442 ,n1419 ,n1395);
    nand g380(n1084 ,n12[11] ,n1012);
    xnor g381(n69 ,n24 ,n9[4]);
    nand g382(n1430 ,n1475 ,n9[11]);
    nand g383(n1010 ,n999 ,n1009);
    nor g384(n334 ,n193 ,n285);
    nor g385(n309 ,n134 ,n231);
    xnor g386(n81 ,n10[7] ,n9[7]);
    nand g387(n1547 ,n10[5] ,n1538);
    nand g388(n1327 ,n1084 ,n1236);
    dff g389(.RN(n1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n8[11]));
    xnor g390(n124 ,n10[5] ,n9[9]);
    nand g391(n745 ,n730 ,n708);
    nand g392(n866 ,n1515 ,n12[1]);
    or g393(n480 ,n301 ,n406);
    nor g394(n1360 ,n1203 ,n1350);
    xnor g395(n742 ,n701 ,n682);
    xor g396(n13[12] ,n907 ,n14[12]);
    not g397(n996 ,n995);
    nand g398(n1318 ,n1126 ,n1227);
    dff g399(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[6]), .Q(n9[6]));
    not g400(n594 ,n593);
    nor g401(n245 ,n59 ,n214);
    nand g402(n1101 ,n11[2] ,n1029);
    xnor g403(n1498 ,n1572 ,n1559);
    nand g404(n1262 ,n1172 ,n1199);
    not g405(n650 ,n645);
    nor g406(n1352 ,n977 ,n1343);
    nand g407(n1359 ,n1338 ,n1296);
    or g408(n1213 ,n1075 ,n1186);
    nor g409(n972 ,n950 ,n971);
    not g410(n931 ,n1446);
    nor g411(n153 ,n111 ,n54);
    not g412(n1536 ,n9[3]);
    xnor g413(n1555 ,n9[8] ,n10[8]);
    nor g414(n413 ,n354 ,n338);
    not g415(n927 ,n1461);
    xnor g416(n825 ,n9[6] ,n10[6]);
    xor g417(n1448 ,n10[1] ,n996);
    nand g418(n1357 ,n1341 ,n1300);
    nand g419(n426 ,n305 ,n309);
    nand g420(n1186 ,n13[15] ,n1087);
    xnor g421(n675 ,n613 ,n633);
    nor g422(n242 ,n88 ,n215);
    xnor g423(n531 ,n338 ,n451);
    nand g424(n1168 ,n1523 ,n1093);
    nor g425(n1436 ,n944 ,n976);
    nor g426(n379 ,n136 ,n226);
    nand g427(n1441 ,n1394 ,n1413);
    not g428(n1018 ,n9[1]);
    not g429(n826 ,n825);
    xnor g430(n1454 ,n10[7] ,n1007);
    nand g431(n1256 ,n1165 ,n1199);
    nor g432(n346 ,n157 ,n273);
    nor g433(n838 ,n815 ,n837);
    not g434(n830 ,n829);
    xnor g435(n657 ,n576 ,n549);
    nor g436(n221 ,n116 ,n215);
    nor g437(n179 ,n131 ,n53);
    or g438(n392 ,n315 ,n298);
    nor g439(n218 ,n69 ,n214);
    or g440(n901 ,n14[11] ,n900);
    xnor g441(n79 ,n10[7] ,n9[9]);
    nand g442(n695 ,n589 ,n670);
    xnor g443(n73 ,n10[3] ,n9[9]);
    nand g444(n514 ,n389 ,n491);
    dff g445(.RN(n1), .SN(1'b1), .CK(n0), .D(n1377), .Q(n8[0]));
    not g446(n27 ,n10[7]);
    nor g447(n524 ,n414 ,n486);
    not g448(n1393 ,n1391);
    nand g449(n40 ,n23 ,n10[8]);
    nand g450(n1156 ,n16[11] ,n1100);
    nand g451(n417 ,n338 ,n358);
    nor g452(n1206 ,n1062 ,n1109);
    nor g453(n204 ,n32 ,n77);
    not g454(n32 ,n10[0]);
    not g455(n1020 ,n9[8]);
    xnor g456(n1553 ,n9[3] ,n10[3]);
    not g457(n1215 ,n1118);
    nor g458(n858 ,n1521 ,n12[7]);
    xnor g459(n680 ,n622 ,n619);
    xor g460(n1473 ,n9[4] ,n987);
    nor g461(n200 ,n32 ,n72);
    or g462(n759 ,n737 ,n741);
    dff g463(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[7]), .Q(n9[7]));
    nand g464(n693 ,n534 ,n657);
    nor g465(n347 ,n146 ,n244);
    nand g466(n1428 ,n1450 ,n1391);
    nor g467(n1005 ,n10[4] ,n1004);
    nand g468(n1309 ,n1082 ,n1218);
    nand g469(n1329 ,n1083 ,n1238);
    nor g470(n370 ,n158 ,n278);
    nand g471(n846 ,n830 ,n845);
    nor g472(n396 ,n351 ,n367);
    dff g473(.RN(n1), .SN(1'b1), .CK(n0), .D(n1310), .Q(n12[4]));
    nor g474(n889 ,n870 ,n888);
    xor g475(n20 ,n295 ,n335);
    nor g476(n1365 ,n1202 ,n1349);
    xnor g477(n1512 ,n822 ,n849);
    not g478(n51 ,n50);
    nor g479(n676 ,n629 ,n660);
    xor g480(n1455 ,n10[8] ,n1008);
    nand g481(n1248 ,n1127 ,n1137);
    nor g482(n406 ,n294 ,n326);
    xnor g483(n625 ,n436 ,n541);
    nor g484(n144 ,n79 ,n53);
    dff g485(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[9]), .Q(n10[9]));
    dff g486(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[8]), .Q(n10[8]));
    nor g487(n336 ,n206 ,n284);
    nand g488(n1569 ,n1554 ,n1568);
    nand g489(n1258 ,n1162 ,n1121);
    nand g490(n779 ,n759 ,n778);
    dff g491(.RN(n1), .SN(1'b1), .CK(n0), .D(n1312), .Q(n12[3]));
    nor g492(n1373 ,n1204 ,n1346);
    dff g493(.RN(n1), .SN(1'b1), .CK(n0), .D(n1381), .Q(n8[7]));
    not g494(n546 ,n545);
    nor g495(n632 ,n506 ,n588);
    nor g496(n1205 ,n1061 ,n1107);
    nand g497(n970 ,n942 ,n969);
    xnor g498(n821 ,n9[10] ,n10[10]);
    not g499(n1194 ,n1088);
    nand g500(n793 ,n690 ,n792);
    nand g501(n527 ,n399 ,n495);
    xnor g502(n1554 ,n9[4] ,n10[4]);
    or g503(n389 ,n304 ,n318);
    nand g504(n1138 ,n1509 ,n1103);
    xnor g505(n455 ,n309 ,n305);
    nor g506(n994 ,n9[10] ,n993);
    nand g507(n845 ,n810 ,n844);
    not g508(n1000 ,n10[7]);
    nand g509(n1046 ,n977 ,n1012);
    nand g510(n1283 ,n1440 ,n1153);
    nor g511(n803 ,n9[5] ,n10[5]);
    nor g512(n326 ,n154 ,n247);
    nand g513(n1130 ,n1512 ,n1103);
    dff g514(.RN(n1), .SN(1'b1), .CK(n0), .D(n1328), .Q(n12[10]));
    nand g515(n1323 ,n1138 ,n1232);
    nor g516(n609 ,n520 ,n546);
    nor g517(n640 ,n525 ,n596);
    xnor g518(n593 ,n504 ,n526);
    or g519(n1387 ,n1326 ,n1380);
    xnor g520(n114 ,n10[9] ,n9[6]);
    xnor g521(n681 ,n625 ,n595);
    xor g522(n1492 ,n1528 ,n10[0]);
    xnor g523(n564 ,n300 ,n453);
    not g524(n658 ,n657);
    nand g525(n1579 ,n1557 ,n1578);
    nand g526(n1277 ,n1185 ,n1199);
    xnor g527(n451 ,n358 ,n327);
    nand g528(n949 ,n1464 ,n919);
    nand g529(n98 ,n27 ,n40);
    dff g530(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[0]), .Q(n11[0]));
    nor g531(n935 ,n929 ,n1460);
    xnor g532(n816 ,n9[4] ,n10[4]);
    nor g533(n1366 ,n1090 ,n1352);
    dff g534(.RN(n1), .SN(1'b1), .CK(n0), .D(n1315), .Q(n12[0]));
    dff g535(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[6]), .Q(n10[6]));
    dff g536(.RN(n1), .SN(1'b1), .CK(n0), .D(n1378), .Q(n8[10]));
    nand g537(n1080 ,n12[10] ,n1012);
    nand g538(n751 ,n747 ,n743);
    or g539(n664 ,n609 ,n634);
    nand g540(n1358 ,n1342 ,n1301);
    nand g541(n1379 ,n1251 ,n1365);
    not g542(n1201 ,n1194);
    nand g543(n380 ,n168 ,n307);
    xnor g544(n452 ,n346 ,n348);
    or g545(n399 ,n348 ,n346);
    nand g546(n1174 ,n1522 ,n1093);
    nand g547(n1165 ,n1512 ,n1100);
    nand g548(n292 ,n10[7] ,n210);
    not g549(n1585 ,n1584);
    or g550(n715 ,n671 ,n679);
    nand g551(n991 ,n983 ,n990);
    xnor g552(n547 ,n466 ,n373);
    nand g553(n662 ,n606 ,n630);
    not g554(n875 ,n874);
    nand g555(n667 ,n613 ,n633);
    nor g556(n308 ,n217 ,n283);
    or g557(n36 ,n23 ,n10[2]);
    nand g558(n1320 ,n1130 ,n1229);
    xnor g559(n686 ,n21 ,n550);
    not g560(n367 ,n366);
    nand g561(n164 ,n47 ,n53);
    xnor g562(n91 ,n23 ,n10[5]);
    nor g563(n1301 ,n1281 ,n1280);
    nor g564(n1208 ,n1050 ,n1120);
    not g565(n551 ,n550);
    xnor g566(n44 ,n25 ,n10[10]);
    xnor g567(n1494 ,n1564 ,n1562);
    nor g568(n216 ,n32 ,n128);
    nand g569(n1170 ,n1503 ,n1100);
    xnor g570(n1508 ,n824 ,n841);
    nand g571(n971 ,n947 ,n970);
    nor g572(n862 ,n1519 ,n12[5]);
    nand g573(n773 ,n706 ,n772);
    nor g574(n235 ,n90 ,n164);
    nand g575(n1254 ,n1161 ,n1160);
    nor g576(n412 ,n357 ,n349);
    nor g577(n643 ,n524 ,n599);
    nor g578(n318 ,n176 ,n289);
    xnor g579(n552 ,n463 ,n322);
    dff g580(.RN(n1), .SN(1'b1), .CK(n0), .D(n1379), .Q(n8[1]));
    nand g581(n1402 ,n10[3] ,n1393);
    nor g582(n885 ,n877 ,n884);
    nor g583(n1212 ,n1042 ,n1122);
    nand g584(n1004 ,n998 ,n1003);
    nor g585(n278 ,n86 ,n214);
    nand g586(n902 ,n14[11] ,n900);
    nand g587(n892 ,n864 ,n891);
    or g588(n706 ,n669 ,n678);
    nand g589(n777 ,n753 ,n776);
    nor g590(n255 ,n76 ,n165);
    xnor g591(n127 ,n10[9] ,n9[2]);
    nor g592(n208 ,n32 ,n133);
    xnor g593(n1516 ,n702 ,n767);
    nor g594(n1103 ,n1015 ,n1037);
    nor g595(n157 ,n70 ,n53);
    nor g596(n378 ,n137 ,n250);
    not g597(n918 ,n1441);
    nor g598(n1342 ,n1282 ,n1324);
    nor g599(n424 ,n316 ,n360);
    nor g600(n176 ,n107 ,n100);
    nor g601(n1339 ,n1270 ,n1321);
    nor g602(n202 ,n32 ,n118);
    not g603(n529 ,n518);
    not g604(n819 ,n818);
    nor g605(n359 ,n190 ,n277);
    nor g606(n1202 ,n1051 ,n1108);
    xnor g607(n743 ,n700 ,n662);
    nand g608(n1349 ,n1333 ,n1292);
    xor g609(n1479 ,n9[10] ,n993);
    not g610(n1026 ,n9[5]);
    nand g611(n1276 ,n1187 ,n1136);
    not g612(n1539 ,n9[2]);
    or g613(n1041 ,n1013 ,n9[11]);
    not g614(n921 ,n1445);
    nor g615(n251 ,n87 ,n163);
    buf g616(n1115 ,n1098);
    nand g617(n1467 ,n1415 ,n1412);
    nor g618(n361 ,n160 ,n274);
    or g619(n907 ,n903 ,n904);
    nor g620(n271 ,n121 ,n215);
    nor g621(n1214 ,n14[15] ,n1115);
    nor g622(n305 ,n156 ,n239);
    nand g623(n1267 ,n10[0] ,n1153);
    nor g624(n728 ,n661 ,n703);
    not g625(n569 ,n568);
    nor g626(n281 ,n64 ,n162);
    nor g627(n1371 ,n1209 ,n1357);
    nand g628(n867 ,n1514 ,n12[0]);
    dff g629(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[11]), .Q(n1388));
    not g630(n802 ,n801);
    nand g631(n1577 ,n1555 ,n1576);
    xnor g632(n573 ,n298 ,n524);
    nand g633(n1594 ,n1525 ,n19[2]);
    nor g634(n180 ,n69 ,n102);
    or g635(n34 ,n23 ,n10[6]);
    nor g636(n173 ,n31 ,n54);
    nor g637(n512 ,n387 ,n482);
    nor g638(n1032 ,n14[14] ,n14[13]);
    nand g639(n1125 ,n9[10] ,n1096);
    xnor g640(n89 ,n10[1] ,n9[8]);
    nor g641(n805 ,n9[10] ,n10[10]);
    nor g642(n946 ,n922 ,n1441);
    nand g643(n1382 ,n1275 ,n1370);
    nor g644(n154 ,n73 ,n54);
    nor g645(n1045 ,n1017 ,n10[9]);
    nand g646(n425 ,n313 ,n314);
    or g647(n419 ,n305 ,n309);
    xnor g648(n1561 ,n9[7] ,n10[7]);
    dff g649(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[3]), .Q(n10[3]));
    nand g650(n1572 ,n1547 ,n1571);
    xnor g651(n1601 ,n1598 ,n1589);
    xnor g652(n87 ,n10[1] ,n9[7]);
    nand g653(n1431 ,n1476 ,n9[11]);
    nor g654(n358 ,n171 ,n234);
    xnor g655(n75 ,n10[9] ,n9[7]);
    nand g656(n1171 ,n1500 ,n1095);
    not g657(n22 ,n9[0]);
    nand g658(n1229 ,n1466 ,n1200);
    xnor g659(n750 ,n708 ,n730);
    nand g660(n669 ,n578 ,n648);
    xnor g661(n1602 ,n1597 ,n1587);
    nor g662(n350 ,n205 ,n255);
    nand g663(n1427 ,n1454 ,n1391);
    xnor g664(n595 ,n471 ,n516);
    nand g665(n687 ,n632 ,n659);
    nand g666(n1275 ,n1442 ,n1153);
    or g667(n385 ,n361 ,n312);
    nor g668(n1300 ,n1277 ,n1276);
    xnor g669(n13[11] ,n905 ,n12[11]);
    not g670(n1525 ,n1);
    nor g671(n674 ,n583 ,n643);
    nor g672(n973 ,n948 ,n972);
    nor g673(n328 ,n152 ,n240);
    nor g674(n1001 ,n10[1] ,n996);
    xnor g675(n463 ,n169 ,n303);
    xnor g676(n1452 ,n10[5] ,n1005);
    nand g677(n1185 ,n1508 ,n1100);
    nand g678(n528 ,n415 ,n498);
    nand g679(n1429 ,n1458 ,n1391);
    dff g680(.RN(n1), .SN(1'b1), .CK(n0), .D(n1387), .Q(n7));
    nor g681(n342 ,n191 ,n252);
    nand g682(n1439 ,n1428 ,n1402);
    xnor g683(n1486 ,n870 ,n888);
    nor g684(n226 ,n103 ,n164);
    not g685(n1017 ,n9[9]);
    nand g686(n795 ,n641 ,n794);
    nand g687(n1176 ,n1499 ,n1095);
    xnor g688(n128 ,n10[1] ,n9[11]);
    nor g689(n330 ,n216 ,n267);
    xnor g690(n541 ,n459 ,n329);
    nor g691(n313 ,n140 ,n235);
    xnor g692(n831 ,n9[2] ,n10[2]);
    nor g693(n217 ,n117 ,n54);
    nand g694(n850 ,n823 ,n849);
    nand g695(n791 ,n720 ,n790);
    nand g696(n1274 ,n1183 ,n1184);
    nor g697(n1040 ,n1014 ,n11[0]);
    or g698(n744 ,n730 ,n708);
    nand g699(n1440 ,n1432 ,n1406);
    nor g700(n583 ,n297 ,n536);
    nand g701(n1356 ,n1298 ,n1335);
    nor g702(n485 ,n378 ,n397);
    not g703(n1105 ,n1104);
    nand g704(n1345 ,n1302 ,n1304);
    nand g705(n1157 ,n1502 ,n1095);
    xnor g706(n464 ,n312 ,n361);
    nor g707(n1207 ,n1065 ,n1110);
    nand g708(n705 ,n662 ,n677);
    nand g709(n947 ,n1466 ,n917);
    xnor g710(n874 ,n1524 ,n12[10]);
    nand g711(n1355 ,n1340 ,n1299);
    xnor g712(n685 ,n624 ,n566);
    dff g713(.RN(n1), .SN(1'b1), .CK(n0), .D(n1605), .Q(n6));
    nand g714(n1161 ,n1491 ,n1091);
    nor g715(n410 ,n170 ,n369);
    not g716(n1529 ,n10[11]);
    nand g717(n732 ,n696 ,n709);
    xnor g718(n45 ,n23 ,n24);
    nor g719(n227 ,n83 ,n215);
    nor g720(n937 ,n926 ,n1443);
    or g721(n1363 ,n1114 ,n1348);
    dff g722(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1600), .Q(n1604));
    xnor g723(n68 ,n10[7] ,n9[8]);
    nor g724(n1306 ,n1076 ,n1213);
    nor g725(n857 ,n1517 ,n12[3]);
    not g726(n1014 ,n11[1]);
    nand g727(n1155 ,n14[11] ,n1093);
    nand g728(n1239 ,n1489 ,n1152);
    nand g729(n1228 ,n1467 ,n1200);
    buf g730(n1480 ,n994);
    nor g731(n274 ,n91 ,n165);
    not g732(n1024 ,n9[3]);
    nand g733(n1197 ,n1484 ,n1091);
    xnor g734(n1519 ,n739 ,n774);
    xnor g735(n105 ,n10[7] ,n9[2]);
    xnor g736(n1500 ,n1576 ,n1555);
    nand g737(n910 ,n908 ,n906);
    nand g738(n1408 ,n10[8] ,n1393);
    nor g739(n992 ,n9[8] ,n991);
    not g740(n408 ,n380);
    not g741(n926 ,n1465);
    or g742(n338 ,n147 ,n275);
    xnor g743(n72 ,n10[1] ,n9[4]);
    nand g744(n516 ,n419 ,n493);
    nand g745(n1227 ,n1468 ,n1200);
    nor g746(n259 ,n111 ,n215);
    nor g747(n627 ,n547 ,n618);
    not g748(n317 ,n316);
    nor g749(n178 ,n124 ,n100);
    nor g750(n964 ,n946 ,n963);
    nand g751(n692 ,n604 ,n665);
    nand g752(n210 ,n34 ,n97);
    nor g753(n171 ,n85 ,n51);
    dff g754(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[2]), .Q(n9[2]));
    nor g755(n897 ,n876 ,n896);
    xnor g756(n678 ,n621 ,n634);
    nand g757(n788 ,n744 ,n787);
    nor g758(n586 ,n437 ,n541);
    nor g759(n150 ,n67 ,n100);
    or g760(n481 ,n327 ,n386);
    nand g761(n41 ,n23 ,n10[4]);
    nor g762(n287 ,n127 ,n162);
    nor g763(n506 ,n344 ,n503);
    nand g764(n290 ,n10[5] ,n209);
    xnor g765(n653 ,n591 ,n533);
    nor g766(n1369 ,n1206 ,n1354);
    nand g767(n556 ,n404 ,n516);
    nand g768(n1144 ,n9[2] ,n1096);
    nand g769(n1383 ,n1279 ,n1371);
    nand g770(n811 ,n9[7] ,n10[7]);
    nor g771(n984 ,n9[1] ,n979);
    or g772(n638 ,n533 ,n591);
    xnor g773(n54 ,n10[2] ,n10[1]);
    not g774(n799 ,n9[0]);
    nand g775(n1250 ,n1155 ,n1156);
    not g776(n299 ,n300);
    xnor g777(n65 ,n10[3] ,n9[10]);
    nand g778(n579 ,n522 ,n549);
    or g779(n494 ,n329 ,n445);
    nor g780(n296 ,n198 ,n246);
    nor g781(n275 ,n62 ,n214);
    nand g782(n1412 ,n9[9] ,n1392);
    nand g783(n498 ,n300 ,n431);
    nand g784(n735 ,n637 ,n723);
    nand g785(n1578 ,n1546 ,n1577);
    xnor g786(n460 ,n304 ,n318);
    nand g787(n293 ,n10[9] ,n212);
    nand g788(n1589 ,n1597 ,n1588);
    not g789(n916 ,n915);
    nand g790(n809 ,n9[11] ,n802);
    nand g791(n1260 ,n1445 ,n1153);
    nor g792(n1294 ,n1253 ,n1252);
    xnor g793(n1491 ,n898 ,n874);
    nand g794(n420 ,n315 ,n298);
    xnor g795(n633 ,n554 ,n552);
    nor g796(n239 ,n84 ,n162);
    nand g797(n1109 ,n1058 ,n1102);
    xnor g798(n1513 ,n821 ,n851);
    xnor g799(n95 ,n23 ,n10[9]);
    nand g800(n1106 ,n1054 ,n1102);
    nor g801(n1364 ,n1208 ,n1347);
    nor g802(n232 ,n67 ,n165);
    nand g803(n1461 ,n1422 ,n1399);
    nor g804(n319 ,n176 ,n229);
    xnor g805(n659 ,n574 ,n532);
    nor g806(n1009 ,n10[8] ,n1008);
    not g807(n567 ,n566);
    nor g808(n311 ,n175 ,n245);
    nor g809(n371 ,n139 ,n270);
    nand g810(n1582 ,n1545 ,n1581);
    nand g811(n792 ,n715 ,n791);
    not g812(n53 ,n52);
    nand g813(n1541 ,n10[7] ,n1531);
    nand g814(n92 ,n28 ,n43);
    xnor g815(n655 ,n573 ,n536);
    xnor g816(n93 ,n29 ,n10[4]);
    nor g817(n839 ,n804 ,n838);
    nand g818(n1251 ,n1437 ,n1153);
    or g819(n500 ,n418 ,n437);
    nand g820(n1071 ,n12[0] ,n1012);
    nand g821(n1246 ,n1149 ,n1167);
    nand g822(n1195 ,n1506 ,n1100);
    not g823(n1590 ,n1589);
    nand g824(n1316 ,n1124 ,n1225);
    nand g825(n770 ,n688 ,n769);
    not g826(n997 ,n10[5]);
    nand g827(n783 ,n782 ,n766);
    nor g828(n1335 ,n1307 ,n1258);
    nor g829(n895 ,n868 ,n894);
    xnor g830(n740 ,n697 ,n672);
    dff g831(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[0]), .Q(n10[0]));
    nand g832(n1550 ,n10[2] ,n1539);
    nand g833(n1082 ,n12[5] ,n1012);
    nand g834(n1326 ,n1285 ,n1284);
    nand g835(n1068 ,n12[3] ,n1012);
    nand g836(n1348 ,n1293 ,n1334);
    nand g837(n848 ,n819 ,n847);
    nand g838(n646 ,n528 ,n598);
    xnor g839(n1474 ,n9[5] ,n988);
    not g840(n618 ,n617);
    xnor g841(n534 ,n457 ,n476);
    nor g842(n1370 ,n1207 ,n1355);
    nand g843(n834 ,n806 ,n833);
    or g844(n854 ,n820 ,n853);
    not g845(n439 ,n411);
    nor g846(n220 ,n130 ,n215);
    not g847(n1599 ,n1595);
    xnor g848(n566 ,n473 ,n407);
    not g849(n1527 ,n9[0]);
    nand g850(n1444 ,n1434 ,n1408);
    not g851(n880 ,n879);
    or g852(n555 ,n339 ,n508);
    xnor g853(n71 ,n10[3] ,n9[4]);
    nor g854(n525 ,n391 ,n489);
    nand g855(n515 ,n398 ,n494);
    nor g856(n940 ,n928 ,n1462);
    xnor g857(n739 ,n696 ,n709);
    nand g858(n1092 ,n1015 ,n1040);
    nor g859(n225 ,n72 ,n163);
    nor g860(n289 ,n126 ,n165);
    nand g861(n1188 ,n1519 ,n1093);
    nand g862(n1273 ,n1182 ,n1199);
    or g863(n35 ,n23 ,n10[8]);
    or g864(n405 ,n293 ,n375);
    nand g865(n677 ,n521 ,n656);
    nor g866(n521 ,n402 ,n499);
    nor g867(n1298 ,n1266 ,n1263);
    nand g868(n434 ,n368 ,n302);
    nand g869(n430 ,n348 ,n346);
    nor g870(n1033 ,n14[17] ,n14[16]);
    not g871(n1019 ,n9[2]);
    nand g872(n1122 ,n1069 ,n1102);
    dff g873(.RN(n1), .SN(1'b1), .CK(n0), .D(n1329), .Q(n12[9]));
    nand g874(n712 ,n668 ,n685);
    nand g875(n582 ,n509 ,n565);
    nand g876(n1249 ,n1181 ,n1199);
    nor g877(n1334 ,n1248 ,n1317);
    nor g878(n147 ,n58 ,n102);
    nor g879(n912 ,n911 ,n909);
    nand g880(n847 ,n811 ,n846);
    not g881(n985 ,n984);
    nand g882(n1052 ,n10[10] ,n1025);
    nand g883(n1565 ,n1562 ,n1564);
    dff g884(.RN(n1), .SN(1'b1), .CK(n0), .D(n1383), .Q(n8[5]));
    nand g885(n1575 ,n1561 ,n1574);
    xor g886(n1453 ,n10[6] ,n1006);
    xnor g887(n741 ,n698 ,n684);
    nor g888(n853 ,n805 ,n852);
    xor g889(n1477 ,n9[8] ,n991);
    xnor g890(n60 ,n24 ,n9[1]);
    not g891(n1102 ,n1101);
    not g892(n1530 ,n10[0]);
    nor g893(n302 ,n189 ,n261);
    dff g894(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[2]), .Q(n10[2]));
    nand g895(n214 ,n44 ,n102);
    xnor g896(n1520 ,n764 ,n776);
    nor g897(n376 ,n143 ,n236);
    nor g898(n1088 ,n1073 ,n1078);
    nand g899(n962 ,n938 ,n961);
    xnor g900(n1495 ,n1566 ,n1553);
    xnor g901(n815 ,n9[3] ,n10[3]);
    nor g902(n386 ,n358 ,n338);
    nand g903(n1141 ,n1506 ,n1103);
    buf g904(n909 ,n904);
    nand g905(n955 ,n936 ,n943);
    not g906(n443 ,n426);
    nor g907(n387 ,n169 ,n303);
    xnor g908(n110 ,n10[7] ,n9[11]);
    nand g909(n1151 ,n1605 ,n1091);
    nor g910(n628 ,n584 ,n595);
    or g911(n393 ,n308 ,n340);
    not g912(n1013 ,n11[0]);
    not g913(n437 ,n436);
    nor g914(n195 ,n112 ,n51);
    not g915(n442 ,n425);
    nand g916(n96 ,n30 ,n41);
    nor g917(n484 ,n408 ,n377);
    nand g918(n1325 ,n1143 ,n1235);
    xnor g919(n14[16] ,n577 ,n796);
    xnor g920(n869 ,n1521 ,n12[7]);
    nand g921(n1347 ,n1332 ,n1311);
    nand g922(n723 ,n605 ,n692);
    nand g923(n1131 ,n1504 ,n1103);
    nor g924(n196 ,n82 ,n102);
    or g925(n1361 ,n1151 ,n1352);
    nor g926(n717 ,n614 ,n681);
    xnor g927(n589 ,n470 ,n523);
    not g928(n979 ,n978);
    nor g929(n571 ,n412 ,n519);
    nand g930(n1544 ,n9[11] ,n1529);
    not g931(n26 ,n10[9]);
    nor g932(n348 ,n141 ,n257);
    nand g933(n1322 ,n1135 ,n1231);
    not g934(n817 ,n816);
    nor g935(n1007 ,n10[6] ,n1006);
    xnor g936(n871 ,n1520 ,n12[6]);
    xnor g937(n1510 ,n829 ,n845);
    nor g938(n365 ,n185 ,n266);
    not g939(n297 ,n298);
    nor g940(n1586 ,n1596 ,n1585);
    not g941(n924 ,n1447);
    nand g942(n1460 ,n1421 ,n1398);
    nor g943(n183 ,n88 ,n54);
    nand g944(n1354 ,n1339 ,n1297);
    xnor g945(n536 ,n460 ,n325);
    nand g946(n1086 ,n10[3] ,n1024);
    nand g947(n1107 ,n1060 ,n1102);
    nand g948(n526 ,n384 ,n496);
    nor g949(n746 ,n718 ,n733);
    or g950(n398 ,n343 ,n342);
    nor g951(n357 ,n161 ,n280);
    xnor g952(n14[14] ,n699 ,n792);
    nor g953(n1367 ,n1211 ,n1353);
    nand g954(n1233 ,n1462 ,n1200);
    xnor g955(n868 ,n1522 ,n12[8]);
    xor g956(n1457 ,n10[10] ,n1010);
    nand g957(n814 ,n800 ,n10[0]);
    nor g958(n886 ,n857 ,n885);
    nand g959(n1069 ,n10[0] ,n1016);
    not g960(n1537 ,n9[8]);
    nor g961(n306 ,n204 ,n268);
    or g962(n37 ,n23 ,n10[4]);
    nand g963(n97 ,n29 ,n42);
    nand g964(n1060 ,n10[8] ,n1020);
    xnor g965(n102 ,n10[10] ,n10[9]);
    xnor g966(n1562 ,n9[2] ,n10[2]);
    xnor g967(n88 ,n10[3] ,n9[5]);
    not g968(n872 ,n871);
    xnor g969(n122 ,n10[7] ,n9[4]);
    nand g970(n1564 ,n1548 ,n1563);
    nor g971(n588 ,n507 ,n552);
    xnor g972(n553 ,n469 ,n321);
    nand g973(n1278 ,n1189 ,n1188);
    not g974(n340 ,n341);
    nand g975(n1378 ,n1255 ,n1360);
    nor g976(n748 ,n716 ,n734);
    nand g977(n1179 ,n1488 ,n1091);
    nor g978(n258 ,n61 ,n214);
    not g979(n446 ,n430);
    nand g980(n561 ,n420 ,n514);
    nor g981(n718 ,n594 ,n684);
    nand g982(n936 ,n1460 ,n929);
    nand g983(n785 ,n751 ,n784);
    dff g984(.RN(n1), .SN(1'b1), .CK(n0), .D(n1376), .Q(n8[2]));
    nand g985(n704 ,n590 ,n686);
    xnor g986(n591 ,n464 ,n511);
    or g987(n752 ,n747 ,n743);
    xnor g988(n14[11] ,n750 ,n786);
    nand g989(n966 ,n951 ,n965);
    nor g990(n965 ,n954 ,n964);
    nor g991(n397 ,n319 ,n356);
    not g992(n982 ,n9[9]);
    xnor g993(n1522 ,n762 ,n780);
    not g994(n980 ,n9[5]);
    xor g995(n1482 ,n873 ,n867);
    nor g996(n238 ,n79 ,n164);
    nand g997(n1432 ,n1451 ,n1391);
    xnor g998(n763 ,n743 ,n747);
    xnor g999(n113 ,n10[5] ,n9[5]);
    nand g1000(n1241 ,n1159 ,n1199);
    nor g1001(n250 ,n55 ,n214);
    xnor g1002(n115 ,n10[9] ,n9[1]);
    nand g1003(n1346 ,n1337 ,n1295);
    xnor g1004(n100 ,n10[4] ,n10[3]);
    nand g1005(n1464 ,n1430 ,n1404);
    not g1006(n444 ,n428);
    nor g1007(n961 ,n940 ,n960);
    nand g1008(n938 ,n1439 ,n927);
    xor g1009(n1503 ,n800 ,n10[0]);
    nor g1010(n323 ,n203 ,n225);
    dff g1011(.RN(n1), .SN(1'b1), .CK(n0), .D(n1330), .Q(n12[8]));
    xnor g1012(n132 ,n10[5] ,n9[7]);
    not g1013(n1093 ,n1092);
    xor g1014(n1475 ,n9[6] ,n989);
    nor g1015(n181 ,n123 ,n100);
    nor g1016(n1552 ,n1530 ,n1528);
    nand g1017(n787 ,n745 ,n786);
    nor g1018(n186 ,n66 ,n54);
    nand g1019(n974 ,n941 ,n973);
    nor g1020(n203 ,n32 ,n109);
    nand g1021(n1077 ,n14[17] ,n14[16]);
    not g1022(n535 ,n534);
    nand g1023(n510 ,n390 ,n492);
    nor g1024(n377 ,n135 ,n249);
    nand g1025(n431 ,n370 ,n353);
    nor g1026(n1341 ,n1278 ,n1323);
    xnor g1027(n1559 ,n9[6] ,n10[6]);
    or g1028(n33 ,n23 ,n10[10]);
    nand g1029(n1580 ,n1551 ,n1579);
    nor g1030(n438 ,n295 ,n335);
    nor g1031(n1011 ,n10[10] ,n1010);
    nand g1032(n404 ,n340 ,n308);
    nor g1033(n482 ,n409 ,n322);
    nand g1034(n1410 ,n9[8] ,n1392);
    xnor g1035(n129 ,n10[5] ,n9[1]);
    nand g1036(n428 ,n361 ,n312);
    nand g1037(n836 ,n807 ,n835);
    nor g1038(n1344 ,n1288 ,n1325);
    nand g1039(n617 ,n505 ,n560);
    xnor g1040(n61 ,n24 ,n9[10]);
    nand g1041(n849 ,n808 ,n848);
    not g1042(n1531 ,n9[7]);
    nand g1043(n707 ,n669 ,n678);
    nand g1044(n1173 ,n1489 ,n1091);
    nand g1045(n1415 ,n1478 ,n9[11]);
    nor g1046(n1333 ,n1246 ,n1316);
    not g1047(n565 ,n564);
    nand g1048(n607 ,n405 ,n540);
    nor g1049(n228 ,n109 ,n163);
    or g1050(n644 ,n616 ,n531);
    nand g1051(n1154 ,n1436 ,n1104);
    nand g1052(n1126 ,n16[11] ,n1103);
    nand g1053(n1350 ,n1336 ,n1294);
    nand g1054(n1183 ,n1487 ,n1091);
    xnor g1055(n626 ,n500 ,n538);
    xnor g1056(n13[15] ,n914 ,n14[15]);
    dff g1057(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[1]), .Q(n10[1]));
    not g1058(n449 ,n434);
    nand g1059(n1159 ,n1505 ,n1100);
    nor g1060(n316 ,n217 ,n272);
    nand g1061(n1386 ,n1265 ,n1368);
    nor g1062(n958 ,n955 ,n957);
    xnor g1063(n652 ,n547 ,n617);
    nand g1064(n1108 ,n1063 ,n1102);
    nand g1065(n778 ,n754 ,n777);
    nand g1066(n1353 ,n1344 ,n1303);
    nor g1067(n1293 ,n1250 ,n1249);
    nand g1068(n1433 ,n1477 ,n9[11]);
    nor g1069(n230 ,n114 ,n162);
    nor g1070(n1603 ,n1588 ,n1586);
    not g1071(n364 ,n363);
    nor g1072(n266 ,n115 ,n162);
    nor g1073(n229 ,n107 ,n165);
    nor g1074(n647 ,n512 ,n620);
    nand g1075(n1253 ,n1158 ,n1199);
    nor g1076(n310 ,n153 ,n242);
    nor g1077(n558 ,n439 ,n523);
    nor g1078(n351 ,n172 ,n253);
    nor g1079(n1027 ,n17[12] ,n16[11]);
    nor g1080(n329 ,n151 ,n248);
    not g1081(n998 ,n10[3]);
    nand g1082(n772 ,n713 ,n771);
    nand g1083(n952 ,n1437 ,n920);
    nor g1084(n418 ,n379 ,n333);
    nand g1085(n736 ,n680 ,n722);
    nand g1086(n1438 ,n1423 ,n1405);
    nand g1087(n882 ,n866 ,n881);
    nand g1088(n1187 ,n1497 ,n1095);
    nand g1089(n1400 ,n10[7] ,n1393);
    nand g1090(n1404 ,n9[6] ,n1392);
    xnor g1091(n1456 ,n10[9] ,n1009);
    nor g1092(n374 ,n187 ,n260);
    nand g1093(n1290 ,n1447 ,n1153);
    nor g1094(n969 ,n933 ,n968);
    nand g1095(n1289 ,n1439 ,n1153);
    nand g1096(n1075 ,n13[14] ,n13[13]);
    nor g1097(n135 ,n105 ,n53);
    not g1098(n30 ,n10[3]);
    nor g1099(n307 ,n207 ,n251);
    nand g1100(n1127 ,n13[11] ,n1091);
    xnor g1101(n1521 ,n761 ,n778);
    or g1102(n603 ,n334 ,n572);
    xnor g1103(n563 ,n477 ,n378);
    nand g1104(n891 ,n872 ,n890);
    nor g1105(n172 ,n110 ,n53);
    not g1106(n999 ,n10[9]);
    nor g1107(n976 ,n934 ,n975);
    nand g1108(n1182 ,n1509 ,n1100);
    not g1109(n983 ,n9[7]);
    nand g1110(n1218 ,n1486 ,n1152);
    nor g1111(n373 ,n181 ,n265);
    nor g1112(n285 ,n99 ,n215);
    not g1113(n1023 ,n9[6]);
    nand g1114(n1177 ,n1510 ,n1100);
    not g1115(n441 ,n423);
    nor g1116(n1034 ,n18[12] ,n15[11]);
    nand g1117(n789 ,n736 ,n788);
    nand g1118(n1567 ,n1553 ,n1566);
    nand g1119(n1420 ,n1448 ,n1391);
    dff g1120(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[9]), .Q(n9[9]));
    xnor g1121(n47 ,n27 ,n10[6]);
    nor g1122(n236 ,n60 ,n214);
    not g1123(n542 ,n541);
    nand g1124(n1548 ,n10[1] ,n1535);
    not g1125(n1002 ,n1001);
    xnor g1126(n1523 ,n768 ,n782);
    not g1127(n1447 ,n1429);
    nand g1128(n1119 ,n1052 ,n1102);
    nor g1129(n602 ,n501 ,n538);
    nor g1130(n721 ,n627 ,n676);
    nand g1131(n1057 ,n12[6] ,n1012);
    nand g1132(n578 ,n544 ,n566);
    nor g1133(n182 ,n64 ,n51);
    nor g1134(n262 ,n74 ,n165);
    nor g1135(n199 ,n32 ,n80);
    xnor g1136(n877 ,n1517 ,n12[3]);
    nor g1137(n948 ,n921 ,n1467);
    nor g1138(n572 ,n383 ,n517);
    nor g1139(n1351 ,n1092 ,n1345);
    xnor g1140(n829 ,n9[7] ,n10[7]);
    xnor g1141(n1488 ,n869 ,n892);
    xor g1142(n575 ,n527 ,n405);
    nand g1143(n1242 ,n1146 ,n1145);
    nor g1144(n1296 ,n1262 ,n1261);
    nand g1145(n1063 ,n10[1] ,n1018);
    xnor g1146(n77 ,n10[1] ,n9[10]);
    nand g1147(n613 ,n385 ,n557);
    xnor g1148(n1478 ,n9[9] ,n992);
    not g1149(n548 ,n547);
    dff g1150(.RN(n1), .SN(1'b1), .CK(n0), .D(n1375), .Q(n977));
    nor g1151(n483 ,n328 ,n396);
    xnor g1152(n123 ,n10[5] ,n9[6]);
    xnor g1153(n1487 ,n871 ,n890);
    not g1154(n1598 ,n1594);
    nand g1155(n1112 ,n1056 ,n1102);
    nand g1156(n1073 ,n14[14] ,n14[13]);
    nand g1157(n1049 ,n12[1] ,n1012);
    nand g1158(n1435 ,n1457 ,n1391);
    nand g1159(n1571 ,n1558 ,n1570);
    nand g1160(n295 ,n10[3] ,n213);
    nor g1161(n231 ,n132 ,n165);
    nor g1162(n140 ,n108 ,n53);
    nor g1163(n142 ,n116 ,n54);
    xnor g1164(n1499 ,n1574 ,n1561);
    nor g1165(n189 ,n103 ,n53);
    not g1166(n1469 ,n1417);
    xnor g1167(n683 ,n626 ,n571);
    nor g1168(n416 ,n366 ,n352);
    nor g1169(n253 ,n110 ,n164);
    nand g1170(n1199 ,n1604 ,n1100);
    nor g1171(n986 ,n9[2] ,n985);
    not g1172(n537 ,n536);
    xor g1173(n1451 ,n10[4] ,n1004);
    nand g1174(n1328 ,n1080 ,n1237);
    nor g1175(n244 ,n56 ,n165);
    nor g1176(n1337 ,n1259 ,n1319);
    xnor g1177(n48 ,n26 ,n10[8]);
    buf g1178(n382 ,n336);
    nor g1179(n896 ,n859 ,n895);
    nor g1180(n1050 ,n1019 ,n10[2]);
    xnor g1181(n70 ,n10[7] ,n9[3]);
    not g1182(n930 ,n1467);
    xnor g1183(n818 ,n9[8] ,n10[8]);
    xnor g1184(n55 ,n24 ,n9[5]);
    nand g1185(n637 ,n533 ,n591);
    not g1186(n23 ,n22);
    nand g1187(n1307 ,n1199 ,n1216);
    xnor g1188(n727 ,n685 ,n668);
    not g1189(n1015 ,n11[2]);
    nand g1190(n1219 ,n1460 ,n1200);
    nor g1191(n327 ,n149 ,n222);
    nand g1192(n835 ,n832 ,n834);
    not g1193(n320 ,n319);
    not g1194(n615 ,n614);
    not g1195(n46 ,n10[1]);
    nand g1196(n840 ,n817 ,n839);
    nor g1197(n286 ,n104 ,n163);
    nand g1198(n989 ,n980 ,n988);
    nor g1199(n734 ,n663 ,n717);
    or g1200(n597 ,n405 ,n540);
    nand g1201(n162 ,n48 ,n51);
    nand g1202(n605 ,n438 ,n553);
    xnor g1203(n545 ,n452 ,n331);
    not g1204(n1597 ,n1592);
    xnor g1205(n822 ,n9[9] ,n10[9]);
    nor g1206(n273 ,n105 ,n164);
    nor g1207(n1211 ,n1085 ,n1113);
    nor g1208(n391 ,n306 ,n365);
    nand g1209(n1111 ,n1066 ,n1102);
    not g1210(n24 ,n25);
    nand g1211(n1217 ,n1487 ,n1152);
    nand g1212(n411 ,n338 ,n354);
    nand g1213(n1169 ,n1490 ,n1091);
    nand g1214(n1236 ,n13[11] ,n1152);
    xnor g1215(n14[13] ,n726 ,n790);
    nand g1216(n1563 ,n1552 ,n1560);
    nand g1217(n756 ,n746 ,n742);
    nand g1218(n794 ,n695 ,n793);
    nor g1219(n321 ,n200 ,n219);
    nor g1220(n600 ,n500 ,n539);
    xnor g1221(n654 ,n563 ,n592);
    xnor g1222(n568 ,n461 ,n372);
    nand g1223(n212 ,n35 ,n98);
    nor g1224(n314 ,n183 ,n233);
    nand g1225(n1043 ,n11[0] ,n11[2]);
    nand g1226(n559 ,n339 ,n508);
    nor g1227(n167 ,n31 ,n100);
    nor g1228(n585 ,n474 ,n532);
    nand g1229(n1446 ,n1435 ,n1411);
    xor g1230(n1481 ,n1514 ,n12[0]);
    or g1231(n415 ,n370 ,n353);
    nand g1232(n1181 ,n15[11] ,n1095);
    nor g1233(n322 ,n138 ,n227);
    xnor g1234(n870 ,n1519 ,n12[5]);
    xnor g1235(n466 ,n365 ,n306);
    xnor g1236(n14[15] ,n651 ,n794);
    xnor g1237(n109 ,n10[1] ,n9[5]);
    nand g1238(n841 ,n812 ,n840);
    not g1239(n501 ,n500);
    xnor g1240(n824 ,n9[5] ,n10[5]);
    nor g1241(n353 ,n172 ,n279);
    or g1242(n942 ,n917 ,n1466);
    nand g1243(n1587 ,n1596 ,n1585);
    nand g1244(n1331 ,n1059 ,n1240);
    nor g1245(n580 ,n522 ,n549);
    nor g1246(n1061 ,n1020 ,n10[8]);
    nor g1247(n1292 ,n1244 ,n1245);
    nand g1248(n865 ,n1524 ,n12[10]);
    nor g1249(n298 ,n144 ,n256);
    dff g1250(.RN(n1), .SN(1'b1), .CK(n0), .D(n1384), .Q(n8[4]));
    nand g1251(n1083 ,n12[9] ,n1012);
    nor g1252(n335 ,n208 ,n286);
    nand g1253(n945 ,n1462 ,n928);
    nand g1254(n1397 ,n10[1] ,n1393);
    nand g1255(n1280 ,n1190 ,n1139);
    xnor g1256(n14[12] ,n738 ,n788);
    xnor g1257(n454 ,n314 ,n313);
    nor g1258(n159 ,n56 ,n100);
    nand g1259(n1377 ,n1267 ,n1362);
    nand g1260(n1545 ,n10[10] ,n1532);
    nand g1261(n1321 ,n1133 ,n1230);
    nand g1262(n648 ,n510 ,n587);
    not g1263(n544 ,n543);
    xnor g1264(n78 ,n10[9] ,n9[4]);
    nand g1265(n1414 ,n9[10] ,n1392);
    nor g1266(n722 ,n650 ,n691);
    nand g1267(n1120 ,n1047 ,n1102);
    nand g1268(n1411 ,n10[10] ,n1393);
    not g1269(n28 ,n10[1]);
    nand g1270(n581 ,n299 ,n570);
    buf g1271(n120 ,n9[1]);
    nor g1272(n324 ,n159 ,n232);
    not g1273(n291 ,n290);
    xnor g1274(n67 ,n10[5] ,n9[2]);
    nor g1275(n939 ,n927 ,n1439);
    nand g1276(n1224 ,n1481 ,n1152);
    nor g1277(n337 ,n167 ,n291);
    or g1278(n807 ,n9[2] ,n10[2]);
    xnor g1279(n540 ,n462 ,n371);
    nand g1280(n1166 ,n1495 ,n1095);
    or g1281(n1037 ,n1014 ,n11[0]);
    nor g1282(n414 ,n359 ,n317);
    nand g1283(n1286 ,n1166 ,n1142);
    nand g1284(n1094 ,n1015 ,n1039);
    nor g1285(n145 ,n75 ,n51);
    nand g1286(n1133 ,n1511 ,n1103);
    not g1287(n832 ,n831);
    nand g1288(n900 ,n865 ,n899);
    xor g1289(n1089 ,n9[11] ,n1388);
    not g1290(n450 ,n435);
    nand g1291(n422 ,n306 ,n365);
    or g1292(n688 ,n632 ,n659);
    not g1293(n906 ,n904);
    xnor g1294(n13[16] ,n913 ,n14[16]);
    or g1295(n1028 ,n13[17] ,n13[16]);
    xnor g1296(n724 ,n669 ,n678);
    nor g1297(n1117 ,n1034 ,n1094);
    nor g1298(n1039 ,n1013 ,n11[1]);
    nand g1299(n1162 ,n1492 ,n1095);
    nand g1300(n1271 ,n1443 ,n1153);
    nor g1301(n193 ,n130 ,n54);
    xnor g1302(n550 ,n341 ,n456);
    nand g1303(n689 ,n535 ,n658);
    not g1304(n1022 ,n9[4]);
    nand g1305(n1059 ,n12[7] ,n1012);
    dff g1306(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[0]), .Q(n1389));
    xnor g1307(n504 ,n406 ,n301);
    nor g1308(n1368 ,n1205 ,n1359);
    nor g1309(n223 ,n73 ,n215);
    or g1310(n505 ,n350 ,n475);
    nor g1311(n890 ,n862 ,n889);
    xnor g1312(n697 ,n534 ,n658);
    nand g1313(n1310 ,n1048 ,n1220);
    nand g1314(n1038 ,n11[2] ,n1014);
    nand g1315(n776 ,n732 ,n775);
    xnor g1316(n462 ,n170 ,n369);
    xnor g1317(n111 ,n10[3] ,n9[6]);
    xnor g1318(n554 ,n502 ,n344);
    nor g1319(n716 ,n615 ,n682);
    nand g1320(n1314 ,n1049 ,n1223);
    nor g1321(n883 ,n878 ,n882);
    nor g1322(n403 ,n355 ,n320);
    nor g1323(n194 ,n121 ,n54);
    nand g1324(n1285 ,n1074 ,n1117);
    nand g1325(n1396 ,n9[1] ,n1392);
    xnor g1326(n467 ,n290 ,n323);
    nand g1327(n1192 ,n1485 ,n1091);
    xnor g1328(n104 ,n10[1] ,n9[2]);
    nand g1329(n1463 ,n1426 ,n1409);
    xnor g1330(n543 ,n465 ,n377);
    xnor g1331(n761 ,n737 ,n741);
    or g1332(n713 ,n668 ,n685);
    xnor g1333(n1518 ,n724 ,n772);
    nor g1334(n842 ,n824 ,n841);
    nor g1335(n156 ,n78 ,n51);
    nor g1336(n631 ,n571 ,n600);
    nand g1337(n1374 ,n1260 ,n1373);
    nand g1338(n1282 ,n1192 ,n1193);
    xnor g1339(n1515 ,n675 ,n749);
    not g1340(n855 ,n12[11]);
    not g1341(n1588 ,n1587);
    not g1342(n198 ,n120);
    nor g1343(n272 ,n117 ,n215);
    xnor g1344(n477 ,n355 ,n319);
    nor g1345(n191 ,n119 ,n51);
    dff g1346(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[5]), .Q(n9[5]));
    nand g1347(n1284 ,n1079 ,n1116);
    nor g1348(n499 ,n374 ,n450);
    nor g1349(n629 ,n548 ,n617);
    not g1350(n445 ,n429);
    nor g1351(n990 ,n9[6] ,n989);
    nand g1352(n1148 ,n1504 ,n1100);
    nor g1353(n1096 ,n1041 ,n1038);
    nor g1354(n1153 ,n1436 ,n1105);
    nor g1355(n248 ,n106 ,n164);
    nor g1356(n661 ,n586 ,n628);
    not g1357(n925 ,n1443);
    xnor g1358(n530 ,n475 ,n350);
    nand g1359(n1124 ,n1505 ,n1103);
    dff g1360(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1601), .Q(n19[2]));
    nor g1361(n1210 ,n1055 ,n1112);
    nand g1362(n1592 ,n1525 ,n19[1]);
    not g1363(n978 ,n9[0]);
    nand g1364(n209 ,n37 ,n96);
    xnor g1365(n86 ,n24 ,n9[6]);
    nor g1366(n517 ,n497 ,n382);
    nand g1367(n1423 ,n1449 ,n1391);
    xnor g1368(n56 ,n10[5] ,n9[3]);
    nor g1369(n861 ,n1523 ,n12[9]);
    xnor g1370(n112 ,n10[9] ,n9[9]);
    xor g1371(n1504 ,n827 ,n814);
    nand g1372(n1143 ,n1507 ,n1103);
    xnor g1373(n121 ,n10[3] ,n9[7]);
    nand g1374(n1385 ,n1289 ,n1367);
    not g1375(n1532 ,n9[10]);
    nor g1376(n177 ,n83 ,n54);
    nand g1377(n864 ,n1520 ,n12[6]);
    nor g1378(n333 ,n148 ,n223);
    nand g1379(n1058 ,n10[7] ,n1021);
    or g1380(n1380 ,n1351 ,n1366);
    or g1381(n765 ,n748 ,n755);
    nor g1382(n143 ,n57 ,n102);
    nand g1383(n1549 ,n10[4] ,n1540);
    nand g1384(n1424 ,n1473 ,n9[11]);
    nor g1385(n151 ,n81 ,n53);
    xnor g1386(n1449 ,n10[2] ,n1001);
    nor g1387(n267 ,n77 ,n163);
    nor g1388(n1303 ,n1287 ,n1286);
    not g1389(n447 ,n432);
    xnor g1390(n1493 ,n1560 ,n1552);
    nand g1391(n1066 ,n10[5] ,n1026);
    or g1392(n1302 ,n1077 ,n1234);
    xnor g1393(n873 ,n1515 ,n12[1]);
    xnor g1394(n1471 ,n9[2] ,n984);
    not g1395(n828 ,n827);
    not g1396(n1584 ,n9[0]);
    xnor g1397(n549 ,n458 ,n330);
    nand g1398(n1222 ,n1483 ,n1152);
    not g1399(n503 ,n502);
    nand g1400(n1223 ,n1482 ,n1152);
    xnor g1401(n698 ,n673 ,n593);
    nor g1402(n903 ,n12[11] ,n902);
    nor g1403(n233 ,n71 ,n215);
    xnor g1404(n133 ,n10[1] ,n9[3]);
    xnor g1405(n726 ,n679 ,n671);
    or g1406(n881 ,n867 ,n873);
    nor g1407(n349 ,n188 ,n276);
    nand g1408(n786 ,n752 ,n785);
    nor g1409(n237 ,n89 ,n163);
    nand g1410(n899 ,n875 ,n898);
    nand g1411(n1384 ,n1283 ,n1372);
    xnor g1412(n701 ,n663 ,n615);
    dff g1413(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1602), .Q(n19[1]));
    xnor g1414(n660 ,n575 ,n540);
    nand g1415(n1237 ,n1491 ,n1152);
    nand g1416(n641 ,n616 ,n531);
    or g1417(n598 ,n299 ,n570);
    nor g1418(n402 ,n362 ,n341);
    xnor g1419(n118 ,n10[1] ,n9[9]);
    xnor g1420(n1472 ,n9[3] ,n986);
    nand g1421(n810 ,n9[6] ,n10[6]);
    nor g1422(n911 ,n856 ,n908);
    nor g1423(n139 ,n122 ,n53);
    nand g1424(n1230 ,n1465 ,n1200);
    nand g1425(n590 ,n393 ,n556);
    nand g1426(n1421 ,n1471 ,n9[11]);
    nand g1427(n1266 ,n1198 ,n1131);
    xor g1428(n472 ,n339 ,n311);
    nand g1429(n1076 ,n13[12] ,n13[11]);
    xnor g1430(n106 ,n10[7] ,n9[6]);
    nand g1431(n1128 ,n1513 ,n1103);
    nor g1432(n304 ,n197 ,n218);
    nor g1433(n804 ,n9[3] ,n10[3]);
    nand g1434(n1079 ,n17[12] ,n16[11]);
    nand g1435(n1255 ,n1446 ,n1153);
    nor g1436(n234 ,n85 ,n162);
    nor g1437(n381 ,n168 ,n307);
    not g1438(n682 ,n681);
    xnor g1439(n1511 ,n818 ,n847);
    nor g1440(n968 ,n937 ,n967);
    nand g1441(n436 ,n379 ,n333);
    nand g1442(n639 ,n619 ,n582);
    nand g1443(n636 ,n527 ,n607);
    nand g1444(n1546 ,n10[8] ,n1537);
    nand g1445(n1398 ,n9[2] ,n1392);
    buf g1446(n9[0] ,n1389);
    not g1447(n1016 ,n1389);
    nand g1448(n1140 ,n1508 ,n1103);
    xnor g1449(n476 ,n294 ,n326);
    nand g1450(n1164 ,n1501 ,n1095);
    nand g1451(n587 ,n543 ,n567);
    xnor g1452(n1514 ,n653 ,n723);
    nand g1453(n1225 ,n1459 ,n1200);
    or g1454(n495 ,n331 ,n446);
    nand g1455(n670 ,n581 ,n646);
    nand g1456(n1291 ,n1141 ,n1219);
    xnor g1457(n50 ,n27 ,n10[8]);
    nand g1458(n497 ,n38 ,n400);
    xor g1459(n1526 ,n9[11] ,n1529);
    nor g1460(n519 ,n448 ,n476);
    nor g1461(n860 ,n1516 ,n12[2]);
    nor g1462(n260 ,n81 ,n164);
    nor g1463(n1042 ,n1016 ,n10[0]);
    xnor g1464(n1556 ,n9[10] ,n10[10]);
    dff g1465(.RN(n1), .SN(1'b1), .CK(n0), .D(n1308), .Q(n12[6]));
    buf g1466(n38 ,n22);
    nand g1467(n1137 ,n17[12] ,n1103);
    nand g1468(n1191 ,n1507 ,n1100);
    nor g1469(n747 ,n710 ,n728);
    nand g1470(n1226 ,n1469 ,n1200);
    xnor g1471(n755 ,n725 ,n661);
    nand g1472(n1416 ,n1479 ,n9[11]);
    nor g1473(n1055 ,n1022 ,n10[4]);
    nand g1474(n1272 ,n1180 ,n1134);
    nor g1475(n325 ,n145 ,n230);
    xnor g1476(n475 ,n293 ,n375);
    nand g1477(n1232 ,n1463 ,n1200);
    xnor g1478(n126 ,n10[5] ,n9[10]);
    not g1479(n1533 ,n9[6]);
    nor g1480(n222 ,n58 ,n214);
    nand g1481(n1259 ,n1169 ,n1168);
    nand g1482(n215 ,n49 ,n54);
    nor g1483(n1091 ,n11[2] ,n1044);
    nand g1484(n635 ,n20 ,n610);
    xnor g1485(n103 ,n10[7] ,n9[5]);
    nor g1486(n161 ,n60 ,n102);
    or g1487(n731 ,n696 ,n709);
    nand g1488(n17[12] ,n809 ,n854);
    dff g1489(.RN(n1), .SN(1'b1), .CK(n0), .D(n1331), .Q(n12[7]));
    nand g1490(n1238 ,n1490 ,n1152);
    not g1491(n409 ,n394);
    nor g1492(n190 ,n126 ,n100);
    xnor g1493(n62 ,n24 ,n9[8]);
    dff g1494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1603), .Q(n19[0]));
    nor g1495(n511 ,n388 ,n479);
    nor g1496(n601 ,n509 ,n565);
    nand g1497(n630 ,n515 ,n612);
    nand g1498(n1074 ,n18[12] ,n15[11]);
    nor g1499(n249 ,n108 ,n164);
    xnor g1500(n14[17] ,n472 ,n798);
    not g1501(n801 ,n10[11]);
    not g1502(n101 ,n102);
    buf g1503(n914 ,n912);
    nand g1504(n714 ,n672 ,n693);
    nand g1505(n1006 ,n997 ,n1005);
    xnor g1506(n532 ,n454 ,n324);
    nand g1507(n1466 ,n1433 ,n1410);
    nand g1508(n1407 ,n9[7] ,n1392);
    xnor g1509(n456 ,n374 ,n362);
    nand g1510(n790 ,n729 ,n789);
    nor g1511(n959 ,n935 ,n958);
    xnor g1512(n1524 ,n763 ,n784);
    nand g1513(n1315 ,n1071 ,n1224);
    nor g1514(n372 ,n184 ,n269);
    xnor g1515(n16[11] ,n820 ,n853);
    xnor g1516(n1496 ,n1568 ,n1554);
    nand g1517(n1180 ,n1498 ,n1095);
    xnor g1518(n99 ,n23 ,n10[3]);
    nand g1519(n1244 ,n1148 ,n1199);
    nand g1520(n1142 ,n9[3] ,n1096);
    nand g1521(n1425 ,n1456 ,n1391);
    nand g1522(n1193 ,n1518 ,n1093);
    nand g1523(n1147 ,n1493 ,n1095);
    nand g1524(n1097 ,n1036 ,n1031);
    not g1525(n710 ,n704);
    not g1526(n174 ,n173);
    nor g1527(n486 ,n372 ,n424);
    dff g1528(.RN(n1), .SN(1'b1), .CK(n0), .D(n1327), .Q(n12[11]));
    nand g1529(n798 ,n559 ,n797);
    nand g1530(n1595 ,n1525 ,n1604);
    nand g1531(n1287 ,n1195 ,n1199);
    nor g1532(n300 ,n195 ,n288);
    xnor g1533(n130 ,n10[3] ,n9[1]);
    nand g1534(n1121 ,n1389 ,n1096);
    dff g1535(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[2]), .Q(n11[2]));
    nand g1536(n1573 ,n1559 ,n1572);
    nor g1537(n185 ,n127 ,n51);
    not g1538(n929 ,n1438);
    xnor g1539(n13[17] ,n14[17] ,n916);
    not g1540(n1538 ,n9[5]);
    nor g1541(n894 ,n858 ,n893);
    nand g1542(n168 ,n23 ,n50);
    xnor g1543(n125 ,n10[9] ,n9[8]);
    nor g1544(n261 ,n122 ,n164);
    nand g1545(n813 ,n9[9] ,n10[9]);
    xnor g1546(n85 ,n10[9] ,n9[11]);
    nor g1547(n1065 ,n1023 ,n10[6]);
    xnor g1548(n1497 ,n1570 ,n1558);
    nor g1549(n207 ,n32 ,n89);
    nand g1550(n967 ,n949 ,n966);
    nor g1551(n339 ,n175 ,n258);
    or g1552(n163 ,n10[0] ,n46);
    nand g1553(n1008 ,n1000 ,n1007);
    nor g1554(n268 ,n118 ,n163);
    xnor g1555(n76 ,n10[5] ,n9[4]);
    not g1556(n1099 ,n1100);
    nor g1557(n219 ,n133 ,n163);
    nand g1558(n1139 ,n9[4] ,n1096);
    nand g1559(n394 ,n169 ,n303);
    not g1560(n345 ,n344);
    not g1561(n360 ,n359);
    or g1562(n557 ,n444 ,n511);
    nand g1563(n1234 ,n14[15] ,n1201);
    nand g1564(n767 ,n667 ,n760);
    not g1565(n246 ,n163);
    nand g1566(n1070 ,n12[2] ,n1012);
    nand g1567(n1146 ,n1483 ,n1091);
    xnor g1568(n82 ,n24 ,n9[3]);
    xnor g1569(n634 ,n530 ,n513);
    nand g1570(n1264 ,n1173 ,n1174);
    nor g1571(n668 ,n585 ,n647);
    nor g1572(n148 ,n65 ,n54);
    nand g1573(n1056 ,n10[4] ,n1022);
    xnor g1574(n738 ,n680 ,n722);
    not g1575(n1200 ,n1154);
    nor g1576(n134 ,n74 ,n100);
    nor g1577(n1343 ,n1306 ,n1305);
    nand g1578(n1304 ,n1033 ,n1214);
    nor g1579(n332 ,n201 ,n241);
    nand g1580(n696 ,n611 ,n664);
    nand g1581(n812 ,n9[4] ,n10[4]);
    nand g1582(n1172 ,n1511 ,n1100);
    xnor g1583(n1507 ,n839 ,n816);
    nand g1584(n1419 ,n1453 ,n1391);
    nor g1585(n1035 ,n14[12] ,n14[11]);
    nand g1586(n963 ,n945 ,n962);
    nor g1587(n663 ,n602 ,n631);
    dff g1588(.RN(n1), .SN(1'b1), .CK(n0), .D(n1314), .Q(n12[1]));
    dff g1589(.RN(n1), .SN(1'b1), .CK(n0), .D(n1309), .Q(n12[5]));
    not g1590(n908 ,n903);
    not g1591(n25 ,n10[11]);
    nor g1592(n288 ,n125 ,n162);
    xnor g1593(n1485 ,n886 ,n879);
    nand g1594(n1136 ,n9[5] ,n1096);
    or g1595(n757 ,n746 ,n742);
    nand g1596(n1113 ,n1086 ,n1102);
    xnor g1597(n461 ,n359 ,n316);
    nand g1598(n1158 ,n1513 ,n1100);
    not g1599(n1596 ,n1593);
    not g1600(n922 ,n1463);
    nand g1601(n518 ,n350 ,n475);
    nand g1602(n94 ,n26 ,n39);
    not g1603(n919 ,n1442);
    nand g1604(n1263 ,n1163 ,n1170);
    nor g1605(n241 ,n80 ,n163);
    nor g1606(n341 ,n178 ,n262);
    nor g1607(n146 ,n76 ,n100);
    nand g1608(n769 ,n687 ,n767);
    nand g1609(n433 ,n357 ,n349);
    or g1610(n560 ,n513 ,n529);
    nand g1611(n784 ,n765 ,n783);
    nand g1612(n1313 ,n1070 ,n1222);
    not g1613(n29 ,n10[5]);
    nand g1614(n488 ,n301 ,n406);
    xnor g1615(n1490 ,n896 ,n876);
    nor g1616(n136 ,n106 ,n53);
    xnor g1617(n709 ,n652 ,n660);
    nand g1618(n614 ,n488 ,n562);
    nand g1619(n1269 ,n1177 ,n1199);
    not g1620(n356 ,n355);
    nand g1621(n1413 ,n10[5] ,n1393);
    xnor g1622(n1517 ,n727 ,n770);
    nand g1623(n797 ,n555 ,n796);
    nand g1624(n611 ,n520 ,n546);
    not g1625(n502 ,n421);
    nand g1626(n758 ,n737 ,n741);
    nand g1627(n1190 ,n1496 ,n1095);
    nor g1628(n283 ,n65 ,n215);
    dff g1629(.RN(n1), .SN(1'b1), .CK(n0), .D(n1374), .Q(n8[9]));
    nor g1630(n240 ,n63 ,n214);
    nor g1631(n1203 ,n1053 ,n1119);
    or g1632(n604 ,n438 ,n553);
    not g1633(n1540 ,n9[4]);
    dff g1634(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[4]), .Q(n10[4]));
    nand g1635(n612 ,n550 ,n569);
    nor g1636(n1311 ,n1241 ,n1247);
    nand g1637(n753 ,n721 ,n740);
    nor g1638(n137 ,n86 ,n102);
    nor g1639(n155 ,n125 ,n51);
    nand g1640(n1198 ,n1481 ,n1091);
    dff g1641(.RN(n1), .SN(1'b1), .CK(n0), .D(n1385), .Q(n8[3]));
    nor g1642(n303 ,n199 ,n228);
    nand g1643(n487 ,n407 ,n427);
    nor g1644(n277 ,n124 ,n165);
    nor g1645(n206 ,n32 ,n104);
    nand g1646(n1591 ,n1598 ,n1590);
    nor g1647(n197 ,n55 ,n102);
    nand g1648(n1252 ,n1157 ,n1125);
    nand g1649(n672 ,n597 ,n636);
    nand g1650(n851 ,n813 ,n850);
    nor g1651(n205 ,n113 ,n100);
    dff g1652(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[8]), .Q(n9[8]));
    nand g1653(n1581 ,n1556 ,n1580);
    nand g1654(n1437 ,n1420 ,n1397);
    nor g1655(n257 ,n95 ,n162);
    xnor g1656(n1458 ,n10[11] ,n1011);
    nor g1657(n1029 ,n11[0] ,n11[1]);
    nor g1658(n1362 ,n1212 ,n1356);
    nand g1659(n1098 ,n1032 ,n1035);
endmodule
