module top (n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11);
    input [127:0] n0;
    input [255:0] n1;
    input [63:0] n2;
    input [3:0] n3;
    input [31:0] n4;
    input [4:0] n5;
    input n6, n7, n8;
    output [127:0] n9;
    output [31:0] n10;
    output n11;
    wire [127:0] n0;
    wire [255:0] n1;
    wire [63:0] n2;
    wire [3:0] n3;
    wire [31:0] n4;
    wire [4:0] n5;
    wire n6, n7, n8;
    wire [127:0] n9;
    wire [31:0] n10;
    wire n11;
    wire n12, n13, n14, n15, n16, n17, n18, n19;
    wire n20, n21, n22, n23, n24, n25, n26, n27;
    wire n28, n29, n30, n31, n32, n33, n34, n35;
    wire n36, n37, n38, n39, n40, n41, n42, n43;
    wire n44, n45, n46, n47, n48, n49, n50, n51;
    wire n52, n53, n54, n55, n56, n57, n58, n59;
    wire n60, n61, n62, n63, n64, n65, n66, n67;
    wire n68, n69, n70, n71, n72, n73, n74, n75;
    wire n76, n77, n78, n79, n80, n81, n82, n83;
    wire n84, n85, n86, n87, n88, n89, n90, n91;
    wire n92, n93, n94, n95, n96, n97, n98, n99;
    wire n100, n101, n102, n103, n104, n105, n106, n107;
    wire n108, n109, n110, n111, n112, n113, n114, n115;
    wire n116, n117, n118, n119, n120, n121, n122, n123;
    wire n124, n125, n126, n127, n128, n129, n130, n131;
    wire n132, n133, n134, n135, n136, n137, n138, n139;
    wire n140, n141, n142, n143, n144, n145, n146, n147;
    wire n148, n149, n150, n151, n152, n153, n154, n155;
    wire n156, n157, n158, n159, n160, n161, n162, n163;
    wire n164, n165, n166, n167, n168, n169, n170, n171;
    wire n172, n173, n174, n175, n176, n177, n178, n179;
    wire n180, n181, n182, n183, n184, n185, n186, n187;
    wire n188, n189, n190, n191, n192, n193, n194, n195;
    wire n196, n197, n198, n199, n200, n201, n202, n203;
    wire n204, n205, n206, n207, n208, n209, n210, n211;
    wire n212, n213, n214, n215, n216, n217, n218, n219;
    wire n220, n221, n222, n223, n224, n225, n226, n227;
    wire n228, n229, n230, n231, n232, n233, n234, n235;
    wire n236, n237, n238, n239, n240, n241, n242, n243;
    wire n244, n245, n246, n247, n248, n249, n250, n251;
    wire n252, n253, n254, n255, n256, n257, n258, n259;
    wire n260, n261, n262, n263, n264, n265, n266, n267;
    wire n268, n269, n270, n271, n272, n273, n274, n275;
    wire n276, n277, n278, n279, n280, n281, n282, n283;
    wire n284, n285, n286, n287, n288, n289, n290, n291;
    wire n292, n293, n294, n295, n296, n297, n298, n299;
    wire n300, n301, n302, n303, n304, n305, n306, n307;
    wire n308, n309, n310, n311, n312, n313, n314, n315;
    wire n316, n317, n318, n319, n320, n321, n322, n323;
    wire n324, n325, n326, n327, n328, n329, n330, n331;
    wire n332, n333, n334, n335, n336, n337, n338, n339;
    wire n340, n341, n342, n343, n344, n345, n346, n347;
    wire n348, n349, n350, n351, n352, n353, n354, n355;
    wire n356, n357, n358, n359, n360, n361, n362, n363;
    wire n364, n365, n366, n367, n368, n369, n370, n371;
    wire n372, n373, n374, n375, n376, n377, n378, n379;
    wire n380, n381, n382, n383, n384, n385, n386, n387;
    wire n388, n389, n390, n391, n392, n393, n394, n395;
    wire n396, n397, n398, n399, n400, n401, n402, n403;
    wire n404, n405, n406, n407, n408, n409, n410, n411;
    wire n412, n413, n414, n415, n416, n417, n418, n419;
    wire n420, n421, n422, n423, n424, n425, n426, n427;
    wire n428, n429, n430, n431, n432, n433, n434, n435;
    wire n436, n437, n438, n439, n440, n441, n442, n443;
    wire n444, n445, n446, n447, n448, n449, n450, n451;
    wire n452, n453, n454, n455, n456, n457, n458, n459;
    wire n460, n461, n462, n463, n464, n465, n466, n467;
    wire n468, n469, n470, n471, n472, n473, n474, n475;
    wire n476, n477, n478, n479, n480, n481, n482, n483;
    wire n484, n485, n486, n487, n488, n489, n490, n491;
    wire n492, n493, n494, n495, n496, n497, n498, n499;
    wire n500, n501, n502, n503, n504, n505, n506, n507;
    wire n508, n509, n510, n511, n512, n513, n514, n515;
    wire n516, n517, n518, n519, n520, n521, n522, n523;
    wire n524, n525, n526, n527, n528, n529, n530, n531;
    wire n532, n533, n534, n535, n536, n537, n538, n539;
    wire n540, n541, n542, n543, n544, n545, n546, n547;
    wire n548, n549, n550, n551, n552, n553, n554, n555;
    wire n556, n557, n558, n559, n560, n561, n562, n563;
    wire n564, n565, n566, n567, n568, n569, n570, n571;
    wire n572, n573, n574, n575, n576, n577, n578, n579;
    wire n580, n581, n582, n583, n584, n585, n586, n587;
    wire n588, n589, n590, n591, n592, n593, n594, n595;
    wire n596, n597, n598, n599, n600, n601, n602, n603;
    wire n604, n605, n606, n607, n608, n609, n610, n611;
    wire n612, n613, n614, n615, n616, n617, n618, n619;
    wire n620, n621, n622, n623, n624, n625, n626, n627;
    wire n628, n629, n630, n631, n632, n633, n634, n635;
    wire n636, n637, n638, n639, n640, n641, n642, n643;
    wire n644, n645, n646, n647, n648, n649, n650, n651;
    wire n652, n653, n654, n655, n656, n657, n658, n659;
    wire n660, n661, n662, n663, n664, n665, n666, n667;
    wire n668, n669, n670, n671, n672, n673, n674, n675;
    wire n676, n677, n678, n679, n680, n681, n682, n683;
    wire n684, n685, n686, n687, n688, n689, n690, n691;
    wire n692, n693, n694, n695, n696, n697, n698, n699;
    wire n700, n701, n702, n703, n704, n705, n706, n707;
    wire n708, n709, n710, n711, n712, n713, n714, n715;
    wire n716, n717, n718, n719, n720, n721, n722, n723;
    wire n724, n725, n726, n727, n728, n729, n730, n731;
    wire n732, n733, n734, n735, n736, n737, n738, n739;
    wire n740, n741, n742, n743, n744, n745, n746, n747;
    wire n748, n749, n750, n751, n752, n753, n754, n755;
    wire n756, n757, n758, n759, n760, n761, n762, n763;
    wire n764, n765, n766, n767, n768, n769, n770, n771;
    wire n772, n773, n774, n775, n776, n777, n778, n779;
    wire n780, n781, n782, n783, n784, n785, n786, n787;
    wire n788, n789, n790, n791, n792, n793, n794, n795;
    wire n796, n797, n798, n799, n800, n801, n802, n803;
    wire n804, n805, n806, n807, n808, n809, n810, n811;
    wire n812, n813, n814, n815, n816, n817, n818, n819;
    wire n820, n821, n822, n823, n824, n825, n826, n827;
    wire n828, n829, n830, n831, n832, n833, n834, n835;
    wire n836, n837, n838, n839, n840, n841, n842, n843;
    wire n844, n845, n846, n847, n848, n849, n850, n851;
    wire n852, n853, n854, n855, n856, n857, n858, n859;
    wire n860, n861, n862, n863, n864, n865, n866, n867;
    wire n868, n869, n870, n871, n872, n873, n874, n875;
    wire n876, n877, n878, n879, n880, n881, n882, n883;
    wire n884, n885, n886, n887, n888, n889, n890, n891;
    wire n892, n893, n894, n895, n896, n897, n898, n899;
    wire n900, n901, n902, n903, n904, n905, n906, n907;
    wire n908, n909, n910, n911, n912, n913, n914, n915;
    wire n916, n917, n918, n919, n920, n921, n922, n923;
    wire n924, n925, n926, n927, n928, n929, n930, n931;
    wire n932, n933, n934, n935, n936, n937, n938, n939;
    wire n940, n941, n942, n943, n944, n945, n946, n947;
    wire n948, n949, n950, n951, n952, n953, n954, n955;
    wire n956, n957, n958, n959, n960, n961, n962, n963;
    wire n964, n965, n966, n967, n968, n969, n970, n971;
    wire n972, n973, n974, n975, n976, n977, n978, n979;
    wire n980, n981, n982, n983, n984, n985, n986, n987;
    wire n988, n989, n990, n991, n992, n993, n994, n995;
    wire n996, n997, n998, n999, n1000, n1001, n1002, n1003;
    wire n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011;
    wire n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
    wire n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
    wire n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
    wire n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
    wire n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051;
    wire n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059;
    wire n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067;
    wire n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075;
    wire n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083;
    wire n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091;
    wire n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099;
    wire n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107;
    wire n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115;
    wire n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123;
    wire n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131;
    wire n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139;
    wire n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147;
    wire n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155;
    wire n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163;
    wire n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171;
    wire n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179;
    wire n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187;
    wire n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195;
    wire n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203;
    wire n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
    wire n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219;
    wire n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227;
    wire n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235;
    wire n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243;
    wire n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251;
    wire n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259;
    wire n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267;
    wire n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275;
    wire n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;
    wire n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291;
    wire n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;
    wire n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307;
    wire n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315;
    wire n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323;
    wire n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331;
    wire n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;
    wire n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;
    wire n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;
    wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
    wire n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;
    wire n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;
    wire n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387;
    wire n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395;
    wire n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403;
    wire n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411;
    wire n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419;
    wire n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427;
    wire n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435;
    wire n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443;
    wire n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451;
    wire n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459;
    wire n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467;
    wire n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475;
    wire n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483;
    wire n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491;
    wire n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499;
    wire n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507;
    wire n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515;
    wire n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523;
    wire n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531;
    wire n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539;
    wire n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547;
    wire n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555;
    wire n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563;
    wire n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571;
    wire n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579;
    wire n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587;
    wire n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595;
    wire n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603;
    wire n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611;
    wire n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619;
    wire n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627;
    wire n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635;
    wire n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643;
    wire n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651;
    wire n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659;
    wire n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667;
    wire n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675;
    wire n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683;
    wire n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691;
    wire n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699;
    wire n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707;
    wire n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715;
    wire n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723;
    wire n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731;
    wire n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739;
    wire n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747;
    wire n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755;
    wire n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763;
    wire n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771;
    wire n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779;
    wire n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787;
    wire n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795;
    wire n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803;
    wire n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811;
    wire n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819;
    wire n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827;
    wire n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835;
    wire n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843;
    wire n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851;
    wire n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859;
    wire n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867;
    wire n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875;
    wire n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883;
    wire n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891;
    wire n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899;
    wire n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907;
    wire n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915;
    wire n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923;
    wire n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931;
    wire n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939;
    wire n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947;
    wire n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955;
    wire n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963;
    wire n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971;
    wire n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979;
    wire n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987;
    wire n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995;
    wire n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003;
    wire n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011;
    wire n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019;
    wire n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027;
    wire n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035;
    wire n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043;
    wire n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051;
    wire n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059;
    wire n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067;
    wire n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075;
    wire n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083;
    wire n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091;
    wire n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099;
    wire n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107;
    wire n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115;
    wire n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123;
    wire n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131;
    wire n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139;
    wire n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147;
    wire n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155;
    wire n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163;
    wire n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171;
    wire n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179;
    wire n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187;
    wire n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195;
    wire n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203;
    wire n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211;
    wire n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219;
    wire n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227;
    wire n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235;
    wire n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243;
    wire n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251;
    wire n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259;
    wire n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267;
    wire n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275;
    wire n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283;
    wire n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291;
    wire n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299;
    wire n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307;
    wire n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315;
    wire n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323;
    wire n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331;
    wire n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339;
    wire n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347;
    wire n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355;
    wire n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363;
    wire n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371;
    wire n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379;
    wire n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387;
    wire n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395;
    wire n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403;
    wire n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411;
    wire n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419;
    wire n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427;
    wire n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435;
    wire n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443;
    wire n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451;
    wire n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459;
    wire n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467;
    wire n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475;
    wire n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483;
    wire n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491;
    wire n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499;
    wire n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507;
    wire n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515;
    wire n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523;
    wire n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531;
    wire n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539;
    wire n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547;
    wire n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555;
    wire n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563;
    wire n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571;
    wire n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579;
    wire n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587;
    wire n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595;
    wire n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603;
    wire n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611;
    wire n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619;
    wire n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627;
    wire n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635;
    wire n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643;
    wire n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651;
    wire n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659;
    wire n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667;
    wire n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675;
    wire n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683;
    wire n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691;
    wire n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699;
    wire n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707;
    wire n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715;
    wire n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723;
    wire n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731;
    wire n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739;
    wire n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747;
    wire n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755;
    wire n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763;
    wire n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771;
    wire n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779;
    wire n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787;
    wire n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795;
    wire n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803;
    wire n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811;
    wire n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819;
    wire n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827;
    wire n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835;
    wire n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843;
    wire n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851;
    wire n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859;
    wire n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867;
    wire n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875;
    wire n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883;
    wire n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891;
    wire n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899;
    wire n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907;
    wire n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915;
    wire n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923;
    wire n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931;
    wire n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939;
    wire n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947;
    wire n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955;
    wire n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963;
    wire n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971;
    wire n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979;
    wire n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987;
    wire n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995;
    wire n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003;
    wire n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011;
    wire n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019;
    wire n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027;
    wire n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035;
    wire n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043;
    wire n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051;
    wire n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059;
    wire n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067;
    wire n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075;
    wire n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083;
    wire n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091;
    wire n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099;
    wire n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107;
    wire n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115;
    wire n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123;
    wire n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131;
    wire n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139;
    wire n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147;
    wire n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155;
    wire n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163;
    wire n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171;
    wire n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179;
    wire n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187;
    wire n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195;
    wire n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203;
    wire n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211;
    wire n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219;
    wire n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227;
    wire n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235;
    wire n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243;
    wire n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251;
    wire n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259;
    wire n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267;
    wire n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275;
    wire n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283;
    wire n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291;
    wire n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299;
    wire n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307;
    wire n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315;
    wire n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323;
    wire n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331;
    wire n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339;
    wire n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347;
    wire n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355;
    wire n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363;
    wire n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371;
    wire n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379;
    wire n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387;
    wire n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395;
    wire n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403;
    wire n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411;
    wire n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419;
    wire n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427;
    wire n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435;
    wire n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443;
    wire n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451;
    wire n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459;
    wire n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467;
    wire n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475;
    wire n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483;
    wire n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491;
    wire n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499;
    wire n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507;
    wire n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515;
    wire n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523;
    wire n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531;
    wire n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539;
    wire n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547;
    wire n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555;
    wire n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563;
    wire n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571;
    wire n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579;
    wire n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587;
    wire n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595;
    wire n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603;
    wire n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611;
    wire n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619;
    wire n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627;
    wire n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635;
    wire n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643;
    wire n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651;
    wire n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659;
    wire n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667;
    wire n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675;
    wire n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683;
    wire n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691;
    wire n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699;
    wire n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707;
    wire n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715;
    wire n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723;
    wire n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731;
    wire n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739;
    wire n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747;
    wire n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755;
    wire n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763;
    wire n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771;
    wire n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779;
    wire n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787;
    wire n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795;
    wire n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803;
    wire n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811;
    wire n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819;
    wire n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827;
    wire n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835;
    wire n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843;
    wire n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851;
    wire n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859;
    wire n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867;
    wire n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875;
    wire n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883;
    wire n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891;
    wire n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899;
    wire n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907;
    wire n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915;
    wire n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923;
    wire n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931;
    wire n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939;
    wire n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947;
    wire n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955;
    wire n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963;
    wire n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971;
    wire n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979;
    wire n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987;
    wire n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995;
    wire n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003;
    wire n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011;
    wire n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019;
    wire n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027;
    wire n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035;
    wire n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043;
    wire n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051;
    wire n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059;
    wire n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067;
    wire n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075;
    wire n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083;
    wire n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091;
    wire n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099;
    wire n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107;
    wire n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115;
    wire n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123;
    wire n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131;
    wire n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139;
    wire n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147;
    wire n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155;
    wire n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163;
    wire n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171;
    wire n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179;
    wire n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187;
    wire n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195;
    wire n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203;
    wire n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211;
    wire n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219;
    wire n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227;
    wire n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235;
    wire n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243;
    wire n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251;
    wire n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259;
    wire n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267;
    wire n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275;
    wire n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283;
    wire n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291;
    wire n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299;
    wire n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307;
    wire n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315;
    wire n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323;
    wire n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331;
    wire n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339;
    wire n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347;
    wire n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355;
    wire n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363;
    wire n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371;
    wire n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379;
    wire n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387;
    wire n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395;
    wire n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403;
    wire n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411;
    wire n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419;
    wire n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427;
    wire n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435;
    wire n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443;
    wire n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451;
    wire n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459;
    wire n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467;
    wire n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475;
    wire n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483;
    wire n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491;
    wire n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499;
    wire n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507;
    wire n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515;
    wire n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523;
    wire n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531;
    wire n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539;
    wire n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547;
    wire n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555;
    wire n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563;
    wire n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571;
    wire n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579;
    wire n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587;
    wire n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595;
    wire n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603;
    wire n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611;
    wire n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619;
    wire n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627;
    wire n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635;
    wire n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643;
    wire n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651;
    wire n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659;
    wire n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667;
    wire n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675;
    wire n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683;
    wire n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691;
    wire n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699;
    wire n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707;
    wire n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715;
    wire n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723;
    wire n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731;
    wire n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739;
    wire n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747;
    wire n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755;
    wire n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763;
    wire n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771;
    wire n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779;
    wire n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787;
    wire n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795;
    wire n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803;
    wire n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811;
    wire n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819;
    wire n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827;
    wire n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835;
    wire n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843;
    wire n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851;
    wire n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859;
    wire n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867;
    wire n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875;
    wire n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883;
    wire n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891;
    wire n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899;
    wire n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907;
    wire n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915;
    wire n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923;
    wire n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931;
    wire n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939;
    wire n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947;
    wire n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955;
    wire n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963;
    wire n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971;
    wire n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979;
    wire n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987;
    wire n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995;
    wire n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003;
    wire n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011;
    wire n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019;
    wire n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027;
    wire n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035;
    wire n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043;
    wire n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051;
    wire n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059;
    wire n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067;
    wire n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075;
    wire n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083;
    wire n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091;
    wire n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099;
    wire n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107;
    wire n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115;
    wire n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123;
    wire n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131;
    wire n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139;
    wire n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147;
    wire n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155;
    wire n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163;
    wire n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171;
    wire n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179;
    wire n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187;
    wire n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195;
    wire n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203;
    wire n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211;
    wire n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219;
    wire n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227;
    wire n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235;
    wire n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243;
    wire n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251;
    wire n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259;
    wire n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267;
    wire n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275;
    wire n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283;
    wire n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291;
    wire n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299;
    wire n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307;
    wire n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315;
    wire n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323;
    wire n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331;
    wire n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339;
    wire n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347;
    wire n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355;
    wire n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363;
    wire n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371;
    wire n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379;
    wire n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387;
    wire n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395;
    wire n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403;
    wire n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411;
    wire n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419;
    wire n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427;
    wire n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435;
    wire n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443;
    wire n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451;
    wire n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459;
    wire n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467;
    wire n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475;
    wire n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483;
    wire n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491;
    wire n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499;
    wire n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507;
    wire n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515;
    wire n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523;
    wire n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531;
    wire n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539;
    wire n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547;
    wire n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555;
    wire n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563;
    wire n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571;
    wire n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579;
    wire n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587;
    wire n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595;
    wire n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603;
    wire n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611;
    wire n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619;
    wire n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627;
    wire n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635;
    wire n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643;
    wire n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651;
    wire n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659;
    wire n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667;
    wire n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675;
    wire n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683;
    wire n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691;
    wire n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699;
    wire n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707;
    wire n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715;
    wire n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723;
    wire n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731;
    wire n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739;
    wire n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747;
    wire n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755;
    wire n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763;
    wire n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771;
    wire n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779;
    wire n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787;
    wire n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795;
    wire n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803;
    wire n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811;
    wire n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819;
    wire n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827;
    wire n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835;
    wire n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843;
    wire n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851;
    wire n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859;
    wire n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867;
    wire n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875;
    wire n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883;
    wire n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891;
    wire n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899;
    wire n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907;
    wire n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915;
    wire n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923;
    wire n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931;
    wire n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939;
    wire n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947;
    wire n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955;
    wire n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963;
    wire n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971;
    wire n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979;
    wire n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987;
    wire n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995;
    wire n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003;
    wire n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011;
    wire n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019;
    wire n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027;
    wire n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035;
    wire n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043;
    wire n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051;
    wire n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059;
    wire n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067;
    wire n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075;
    wire n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083;
    wire n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091;
    wire n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099;
    wire n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107;
    wire n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115;
    wire n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123;
    wire n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131;
    wire n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139;
    wire n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147;
    wire n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155;
    wire n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163;
    wire n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171;
    wire n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179;
    wire n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187;
    wire n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195;
    wire n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203;
    wire n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211;
    wire n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219;
    wire n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227;
    wire n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235;
    wire n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243;
    wire n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251;
    wire n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259;
    wire n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267;
    wire n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275;
    wire n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283;
    wire n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291;
    wire n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299;
    wire n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307;
    wire n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315;
    wire n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323;
    wire n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331;
    wire n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339;
    wire n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347;
    wire n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355;
    wire n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363;
    wire n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371;
    wire n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379;
    wire n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387;
    wire n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395;
    wire n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403;
    wire n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411;
    wire n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419;
    wire n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427;
    wire n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435;
    wire n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443;
    wire n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451;
    wire n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459;
    wire n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467;
    wire n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475;
    wire n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483;
    wire n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491;
    wire n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499;
    wire n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507;
    wire n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515;
    wire n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523;
    wire n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531;
    wire n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539;
    wire n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547;
    wire n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555;
    wire n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563;
    wire n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571;
    wire n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579;
    wire n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587;
    wire n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595;
    wire n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603;
    wire n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611;
    wire n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619;
    wire n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627;
    wire n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635;
    wire n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643;
    wire n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651;
    wire n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659;
    wire n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667;
    wire n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675;
    wire n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683;
    wire n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691;
    wire n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699;
    wire n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707;
    wire n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715;
    wire n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723;
    wire n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731;
    wire n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739;
    wire n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747;
    wire n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755;
    wire n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763;
    wire n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771;
    wire n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779;
    wire n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787;
    wire n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795;
    wire n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803;
    wire n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811;
    wire n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819;
    wire n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827;
    wire n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835;
    wire n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843;
    wire n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851;
    wire n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859;
    wire n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867;
    wire n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875;
    wire n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883;
    wire n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891;
    wire n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899;
    wire n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907;
    wire n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915;
    wire n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923;
    wire n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931;
    wire n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939;
    wire n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947;
    wire n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955;
    wire n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963;
    wire n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971;
    wire n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979;
    wire n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987;
    wire n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995;
    wire n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003;
    wire n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011;
    wire n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019;
    wire n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027;
    wire n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035;
    wire n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043;
    wire n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051;
    wire n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059;
    wire n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067;
    wire n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075;
    wire n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083;
    wire n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091;
    wire n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099;
    wire n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107;
    wire n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115;
    wire n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123;
    wire n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131;
    wire n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139;
    wire n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147;
    wire n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155;
    wire n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163;
    wire n7164, n7165, n7166, n7167, n7168;
    nand g0(n670 ,n1[16] ,n621);
    nand g1(n436 ,n326 ,n435);
    nand g2(n6663 ,n0[119] ,n0[87]);
    nor g3(n4931 ,n6 ,n4808);
    xnor g4(n1428 ,n1[13] ,n2[13]);
    xnor g5(n4872 ,n4571 ,n4454);
    xnor g6(n1486 ,n0[27] ,n1[27]);
    nor g7(n5901 ,n713 ,n5833);
    or g8(n4407 ,n722 ,n4223);
    nand g9(n9[20] ,n5761 ,n5965);
    not g10(n6071 ,n6070);
    nor g11(n6323 ,n706 ,n6310);
    nor g12(n3507 ,n1222 ,n2825);
    xnor g13(n5580 ,n4569 ,n5271);
    not g14(n750 ,n0[9]);
    nor g15(n2277 ,n709 ,n1602);
    nand g16(n1971 ,n963 ,n1100);
    nand g17(n450 ,n330 ,n449);
    nand g18(n6454 ,n3446 ,n6351);
    nor g19(n4728 ,n722 ,n4584);
    nor g20(n6006 ,n3350 ,n5904);
    nand g21(n4372 ,n791 ,n4236);
    xnor g22(n102 ,n0[18] ,n7074);
    nor g23(n5422 ,n4997 ,n5278);
    nor g24(n2118 ,n1959 ,n1473);
    xnor g25(n4449 ,n3942 ,n2838);
    nand g26(n4833 ,n1966 ,n4436);
    nor g27(n4207 ,n3552 ,n4082);
    xnor g28(n94 ,n0[10] ,n7066);
    nand g29(n457 ,n371 ,n456);
    nor g30(n3140 ,n1852 ,n2592);
    nand g31(n6992 ,n6627 ,n6816);
    nand g32(n4579 ,n1104 ,n4230);
    xnor g33(n1681 ,n0[115] ,n4[3]);
    not g34(n833 ,n0[119]);
    nor g35(n5876 ,n712 ,n5835);
    nor g36(n2728 ,n1055 ,n2610);
    nand g37(n3778 ,n1179 ,n2768);
    nand g38(n42 ,n7077 ,n0[21]);
    nor g39(n2042 ,n1004 ,n1761);
    nand g40(n4366 ,n2017 ,n3850);
    nand g41(n648 ,n0[65] ,n622);
    not g42(n812 ,n0[65]);
    xnor g43(n1710 ,n0[33] ,n1[49]);
    nor g44(n4250 ,n2325 ,n3962);
    not g45(n743 ,n0[42]);
    nand g46(n6640 ,n1[78] ,n6579);
    nor g47(n2219 ,n1961 ,n1933);
    nand g48(n5821 ,n1953 ,n5589);
    nor g49(n3064 ,n1821 ,n2295);
    xnor g50(n5728 ,n5457 ,n2698);
    nor g51(n3039 ,n1221 ,n2347);
    nand g52(n4093 ,n7141 ,n3468);
    nand g53(n4604 ,n717 ,n4573);
    nor g54(n3063 ,n1808 ,n2288);
    nor g55(n4421 ,n4335 ,n4203);
    xnor g56(n543 ,n6956 ,n0[99]);
    or g57(n174 ,n0[47] ,n1[47]);
    nand g58(n5560 ,n4831 ,n5238);
    xnor g59(n1269 ,n0[92] ,n7120);
    nand g60(n1040 ,n714 ,n805);
    xnor g61(n1675 ,n0[16] ,n4[24]);
    nand g62(n6753 ,n0[32] ,n6737);
    nand g63(n561 ,n507 ,n560);
    nand g64(n1909 ,n0[99] ,n1043);
    nand g65(n437 ,n357 ,n436);
    nand g66(n1142 ,n6911 ,n795);
    nor g67(n2425 ,n1956 ,n1542);
    nand g68(n356 ,n7041 ,n7009);
    nor g69(n3641 ,n840 ,n3038);
    nand g70(n3197 ,n1053 ,n2578);
    or g71(n171 ,n0[56] ,n1[56]);
    nand g72(n3966 ,n0[6] ,n3491);
    nand g73(n6497 ,n6453 ,n6348);
    nand g74(n5843 ,n4390 ,n5642);
    xnor g75(n5205 ,n1644 ,n4839);
    xnor g76(n1607 ,n0[111] ,n1[111]);
    nand g77(n6675 ,n0[123] ,n0[91]);
    or g78(n2998 ,n968 ,n2418);
    nor g79(n5863 ,n706 ,n5842);
    nand g80(n3653 ,n3135 ,n2776);
    or g81(n485 ,n0[125] ,n6982);
    nor g82(n2993 ,n1789 ,n2327);
    nor g83(n4283 ,n827 ,n3879);
    nand g84(n3590 ,n3112 ,n3037);
    nand g85(n3736 ,n6819 ,n3137);
    xnor g86(n2852 ,n0[114] ,n1374);
    xnor g87(n534 ,n6978 ,n0[121]);
    nand g88(n461 ,n353 ,n460);
    xnor g89(n2815 ,n1382 ,n1695);
    nand g90(n9[16] ,n6409 ,n6474);
    nand g91(n6304 ,n6164 ,n6225);
    nor g92(n3174 ,n1977 ,n2325);
    xnor g93(n1679 ,n0[10] ,n4[26]);
    nand g94(n2535 ,n1234 ,n1949);
    not g95(n1488 ,n1487);
    or g96(n3357 ,n1[50] ,n3158);
    nand g97(n7039 ,n6660 ,n7134);
    xnor g98(n1405 ,n1[60] ,n2[60]);
    or g99(n3335 ,n2339 ,n2796);
    not g100(n840 ,n0[86]);
    xor g101(n6832 ,n541 ,n528);
    nand g102(n371 ,n7043 ,n7011);
    nand g103(n1114 ,n6847 ,n795);
    nor g104(n1020 ,n804 ,n0[3]);
    nand g105(n5478 ,n4640 ,n5289);
    xnor g106(n393 ,n6991 ,n7023);
    nor g107(n2753 ,n2073 ,n2117);
    nor g108(n2971 ,n2605 ,n2372);
    xnor g109(n1654 ,n0[46] ,n1[62]);
    or g110(n3414 ,n1954 ,n2855);
    nand g111(n6749 ,n0[47] ,n6737);
    nand g112(n1869 ,n0[84] ,n964);
    not g113(n5454 ,n5453);
    or g114(n2257 ,n721 ,n1527);
    xnor g115(n5064 ,n4664 ,n4671);
    not g116(n5937 ,n5938);
    nand g117(n6986 ,n6693 ,n6822);
    nor g118(n2116 ,n6 ,n1993);
    nor g119(n1806 ,n739 ,n1037);
    not g120(n2941 ,n2940);
    nand g121(n6028 ,n3378 ,n5877);
    nor g122(n3293 ,n1954 ,n2868);
    nor g123(n2189 ,n1956 ,n1597);
    nand g124(n7064 ,n673 ,n626);
    nand g125(n4427 ,n2262 ,n4224);
    nand g126(n1794 ,n733 ,n1014);
    or g127(n6024 ,n5553 ,n5856);
    or g128(n4649 ,n3808 ,n4538);
    xnor g129(n1309 ,n6918 ,n6917);
    nor g130(n3912 ,n2224 ,n3757);
    nor g131(n5159 ,n6824 ,n4923);
    nand g132(n5107 ,n717 ,n4990);
    nand g133(n3556 ,n2440 ,n2723);
    not g134(n5378 ,n5377);
    nand g135(n1085 ,n0[55] ,n793);
    nand g136(n134 ,n20 ,n133);
    xnor g137(n6211 ,n6068 ,n5973);
    nand g138(n4069 ,n787 ,n3525);
    nor g139(n5659 ,n3370 ,n5407);
    nor g140(n4392 ,n3202 ,n4285);
    nor g141(n915 ,n807 ,n0[106]);
    xnor g142(n1304 ,n0[8] ,n4[24]);
    xnor g143(n6870 ,n246 ,n273);
    nand g144(n6786 ,n1[118] ,n7088);
    not g145(n970 ,n969);
    nand g146(n7022 ,n6641 ,n7151);
    nor g147(n1820 ,n740 ,n11);
    nand g148(n3110 ,n0[99] ,n2140);
    nand g149(n1822 ,n0[48] ,n1221);
    nand g150(n1082 ,n0[92] ,n715);
    xnor g151(n1432 ,n1[79] ,n2[15]);
    nand g152(n4344 ,n3646 ,n3867);
    nand g153(n1833 ,n0[35] ,n1221);
    nand g154(n5389 ,n3496 ,n5121);
    nand g155(n1227 ,n0[106] ,n0[104]);
    nand g156(n9[118] ,n5655 ,n5616);
    nand g157(n5790 ,n3281 ,n5638);
    nor g158(n3304 ,n1954 ,n2875);
    nor g159(n1827 ,n741 ,n11);
    nor g160(n4260 ,n710 ,n4114);
    not g161(n5284 ,n5283);
    xor g162(n4901 ,n4458 ,n2853);
    nand g163(n6654 ,n0[74] ,n6579);
    nand g164(n4123 ,n790 ,n3963);
    nor g165(n3176 ,n2567 ,n2495);
    nor g166(n2303 ,n721 ,n1639);
    nor g167(n2297 ,n1956 ,n1589);
    nand g168(n6956 ,n6748 ,n6789);
    nand g169(n4082 ,n720 ,n3701);
    nand g170(n4334 ,n2581 ,n3900);
    xnor g171(n2950 ,n1698 ,n1517);
    nor g172(n6190 ,n5028 ,n6142);
    nand g173(n4305 ,n2782 ,n3866);
    xnor g174(n1535 ,n1[53] ,n1[21]);
    nand g175(n4690 ,n1966 ,n4450);
    nand g176(n3181 ,n1981 ,n2326);
    xnor g177(n6208 ,n6066 ,n6032);
    nand g178(n581 ,n527 ,n580);
    not g179(n2906 ,n2905);
    not g180(n5773 ,n5772);
    nand g181(n6769 ,n0[58] ,n6737);
    nor g182(n4516 ,n3762 ,n4299);
    nand g183(n1908 ,n0[58] ,n996);
    nand g184(n301 ,n204 ,n300);
    nor g185(n5785 ,n1954 ,n5594);
    nor g186(n5154 ,n2228 ,n4883);
    nand g187(n209 ,n0[34] ,n1[34]);
    or g188(n5052 ,n4930 ,n4886);
    nand g189(n6797 ,n1[117] ,n7088);
    nor g190(n2789 ,n1963 ,n2430);
    nand g191(n9[106] ,n6076 ,n6153);
    xnor g192(n6213 ,n6110 ,n5974);
    nand g193(n5248 ,n4862 ,n5070);
    nand g194(n5354 ,n3417 ,n5077);
    nor g195(n5152 ,n3617 ,n4944);
    nor g196(n3887 ,n3353 ,n3352);
    or g197(n2106 ,n719 ,n1507);
    or g198(n3549 ,n2411 ,n3256);
    nor g199(n6729 ,n6826 ,n6589);
    or g200(n494 ,n0[119] ,n6976);
    nand g201(n3935 ,n2159 ,n3634);
    nand g202(n5698 ,n5106 ,n5465);
    nand g203(n4091 ,n7143 ,n3458);
    nor g204(n6104 ,n5998 ,n5986);
    nor g205(n2347 ,n1[87] ,n1957);
    nand g206(n4381 ,n787 ,n4236);
    xnor g207(n245 ,n1[41] ,n0[41]);
    nor g208(n4700 ,n6824 ,n4479);
    nand g209(n3093 ,n1220 ,n2355);
    nand g210(n2537 ,n1183 ,n1860);
    nand g211(n5137 ,n6827 ,n4899);
    xnor g212(n1482 ,n0[30] ,n1[30]);
    nor g213(n5636 ,n5098 ,n5458);
    nor g214(n5140 ,n727 ,n4907);
    nand g215(n1891 ,n0[36] ,n966);
    nor g216(n4258 ,n710 ,n4112);
    xnor g217(n2926 ,n1601 ,n1536);
    nor g218(n4669 ,n882 ,n4469);
    xnor g219(n5017 ,n4360 ,n4680);
    not g220(n1956 ,n718);
    nand g221(n4551 ,n1151 ,n4281);
    xnor g222(n551 ,n6964 ,n0[107]);
    nor g223(n4733 ,n2325 ,n4448);
    nand g224(n2964 ,n2253 ,n2524);
    xnor g225(n5853 ,n5568 ,n4591);
    nand g226(n1112 ,n6944 ,n796);
    nand g227(n6464 ,n5776 ,n6425);
    nand g228(n3212 ,n1185 ,n2100);
    nor g229(n939 ,n0[83] ,n0[80]);
    nor g230(n1798 ,n803 ,n1220);
    xnor g231(n1575 ,n0[53] ,n4[13]);
    nor g232(n5023 ,n4937 ,n4928);
    nor g233(n866 ,n710 ,n0[103]);
    nor g234(n5336 ,n4806 ,n5108);
    nor g235(n3882 ,n3218 ,n3495);
    nand g236(n4297 ,n2577 ,n4090);
    nand g237(n6233 ,n3437 ,n6127);
    nand g238(n5637 ,n5249 ,n5475);
    or g239(n2167 ,n719 ,n1548);
    nand g240(n5290 ,n4701 ,n5086);
    nand g241(n4682 ,n4123 ,n4378);
    or g242(n9[126] ,n5417 ,n5805);
    nand g243(n293 ,n216 ,n292);
    nand g244(n6689 ,n1[94] ,n6580);
    xnor g245(n1298 ,n1[38] ,n4[30]);
    nand g246(n6669 ,n0[121] ,n0[89]);
    nand g247(n3149 ,n1[119] ,n2415);
    nor g248(n3411 ,n1954 ,n2938);
    or g249(n22 ,n7071 ,n0[15]);
    nand g250(n6561 ,n4531 ,n6521);
    xnor g251(n1940 ,n1[85] ,n2[21]);
    nand g252(n5043 ,n4697 ,n4880);
    nand g253(n5922 ,n3610 ,n5756);
    nand g254(n2000 ,n961 ,n1103);
    xnor g255(n529 ,n6973 ,n0[116]);
    nor g256(n4118 ,n793 ,n3931);
    nor g257(n5547 ,n4821 ,n5364);
    xnor g258(n1257 ,n1[46] ,n4[6]);
    nor g259(n3412 ,n1222 ,n2846);
    not g260(n5062 ,n5063);
    nand g261(n1226 ,n0[96] ,n714);
    nor g262(n6705 ,n6826 ,n6609);
    nand g263(n6684 ,n0[78] ,n6580);
    nor g264(n5235 ,n3669 ,n5174);
    xnor g265(n1931 ,n1[110] ,n2[46]);
    nor g266(n6083 ,n3344 ,n5959);
    nor g267(n5366 ,n3515 ,n5148);
    not g268(n757 ,n0[67]);
    xnor g269(n5281 ,n4989 ,n4660);
    nand g270(n3587 ,n0[85] ,n2794);
    nand g271(n2562 ,n0[23] ,n707);
    xnor g272(n1260 ,n1[33] ,n1[1]);
    nand g273(n6804 ,n6581 ,n7110);
    xnor g274(n253 ,n1[49] ,n0[49]);
    not g275(n2949 ,n2948);
    xnor g276(n6891 ,n99 ,n131);
    nand g277(n6692 ,n1[95] ,n6580);
    nor g278(n5774 ,n793 ,n5640);
    nand g279(n1090 ,n0[46] ,n715);
    nor g280(n2014 ,n0[11] ,n1053);
    or g281(n1053 ,n0[10] ,n0[8]);
    xnor g282(n2903 ,n1673 ,n1573);
    or g283(n2199 ,n908 ,n2019);
    nand g284(n6988 ,n6639 ,n6820);
    or g285(n5653 ,n5508 ,n4903);
    nor g286(n4034 ,n3736 ,n2784);
    nand g287(n2591 ,n0[2] ,n1964);
    nor g288(n6122 ,n6097 ,n6078);
    xnor g289(n1285 ,n6842 ,n6840);
    nand g290(n4423 ,n792 ,n4217);
    xnor g291(n1609 ,n0[66] ,n1[66]);
    xnor g292(n4593 ,n4105 ,n4358);
    nand g293(n3589 ,n6827 ,n2822);
    not g294(n5832 ,n5833);
    xnor g295(n6202 ,n5974 ,n6112);
    nand g296(n3397 ,n1952 ,n2932);
    nand g297(n3390 ,n1953 ,n2919);
    nor g298(n4935 ,n3472 ,n4603);
    xnor g299(n5080 ,n4666 ,n4431);
    or g300(n4287 ,n4003 ,n3680);
    or g301(n476 ,n0[112] ,n6969);
    nand g302(n4586 ,n2519 ,n4232);
    nand g303(n2595 ,n714 ,n1795);
    not g304(n2951 ,n2950);
    nor g305(n3528 ,n6825 ,n2840);
    nor g306(n6602 ,n0[125] ,n0[93]);
    nor g307(n2350 ,n1[33] ,n1963);
    nand g308(n683 ,n1[5] ,n621);
    nor g309(n3328 ,n1954 ,n2890);
    nand g310(n3584 ,n0[126] ,n2794);
    nand g311(n7148 ,n6617 ,n6704);
    nor g312(n6534 ,n6477 ,n6501);
    nand g313(n3656 ,n0[3] ,n3077);
    nor g314(n4308 ,n2548 ,n3889);
    nor g315(n3130 ,n839 ,n2639);
    nand g316(n6301 ,n6158 ,n6191);
    nor g317(n4704 ,n1965 ,n4464);
    nand g318(n56 ,n7072 ,n0[16]);
    nand g319(n4498 ,n3689 ,n4173);
    nor g320(n4199 ,n6 ,n4099);
    nand g321(n2529 ,n971 ,n1902);
    nand g322(n6152 ,n3355 ,n6051);
    nand g323(n3103 ,n2596 ,n2436);
    not g324(n803 ,n0[105]);
    nand g325(n1881 ,n0[110] ,n966);
    nor g326(n2232 ,n6 ,n1755);
    nor g327(n4942 ,n6 ,n4811);
    nor g328(n3007 ,n2225 ,n2223);
    nor g329(n3073 ,n1841 ,n2499);
    xor g330(n7121 ,n0[61] ,n0[29]);
    nand g331(n4499 ,n2326 ,n4359);
    xnor g332(n5948 ,n5834 ,n1314);
    nand g333(n7012 ,n6651 ,n7161);
    nand g334(n4282 ,n2115 ,n3990);
    nand g335(n5034 ,n4859 ,n4892);
    nor g336(n6434 ,n3448 ,n6350);
    nand g337(n6140 ,n3282 ,n6048);
    nand g338(n6789 ,n1[99] ,n7088);
    nand g339(n2779 ,n1529 ,n2615);
    or g340(n4721 ,n711 ,n4583);
    nor g341(n4300 ,n2747 ,n3913);
    nand g342(n4014 ,n0[71] ,n3490);
    not g343(n4834 ,n4833);
    nand g344(n3678 ,n791 ,n3261);
    nor g345(n1760 ,n725 ,n915);
    nor g346(n6605 ,n0[101] ,n0[69]);
    xnor g347(n4894 ,n2821 ,n4450);
    nand g348(n1075 ,n0[50] ,n725);
    or g349(n330 ,n7040 ,n7008);
    nor g350(n2385 ,n0[30] ,n721);
    nand g351(n1782 ,n1245 ,n1007);
    nand g352(n3573 ,n1814 ,n3252);
    not g353(n3496 ,n3495);
    nand g354(n4004 ,n0[95] ,n3490);
    nand g355(n202 ,n0[46] ,n1[46]);
    nor g356(n5033 ,n4965 ,n4892);
    nand g357(n4328 ,n2594 ,n3880);
    nor g358(n959 ,n0[118] ,n6);
    nand g359(n9[3] ,n4953 ,n6559);
    nor g360(n942 ,n0[102] ,n715);
    nand g361(n4533 ,n2326 ,n4222);
    nor g362(n3288 ,n1954 ,n2864);
    or g363(n12 ,n7067 ,n0[11]);
    nand g364(n667 ,n1[14] ,n621);
    nand g365(n1019 ,n0[41] ,n751);
    nand g366(n4860 ,n3373 ,n4605);
    nand g367(n6399 ,n5903 ,n6339);
    xnor g368(n4887 ,n4213 ,n4574);
    nand g369(n6100 ,n6019 ,n5783);
    xnor g370(n1316 ,n0[80] ,n7108);
    nor g371(n5878 ,n706 ,n5840);
    or g372(n3857 ,n0[19] ,n3440);
    not g373(n4679 ,n4678);
    xnor g374(n5849 ,n5570 ,n1559);
    xnor g375(n1475 ,n1[68] ,n2[4]);
    not g376(n4460 ,n4459);
    nor g377(n3279 ,n2398 ,n2796);
    xnor g378(n5447 ,n5059 ,n2682);
    xnor g379(n1327 ,n0[112] ,n4[0]);
    nor g380(n5619 ,n5103 ,n5467);
    nand g381(n4803 ,n715 ,n4588);
    nor g382(n4647 ,n4124 ,n4375);
    nor g383(n2416 ,n0[33] ,n1754);
    xnor g384(n1449 ,n1[107] ,n2[43]);
    not g385(n735 ,n0[3]);
    or g386(n5441 ,n4025 ,n5288);
    nand g387(n6744 ,n0[61] ,n6737);
    xnor g388(n5866 ,n5571 ,n1717);
    xnor g389(n5848 ,n5574 ,n5529);
    nand g390(n1241 ,n0[58] ,n765);
    nor g391(n1724 ,n1050 ,n1027);
    xnor g392(n1274 ,n0[113] ,n7109);
    xnor g393(n6145 ,n5970 ,n5639);
    or g394(n4705 ,n1965 ,n4465);
    xnor g395(n6345 ,n6243 ,n6174);
    nand g396(n651 ,n0[69] ,n622);
    nor g397(n5324 ,n4630 ,n5089);
    xnor g398(n6913 ,n378 ,n447);
    xor g399(n6834 ,n237 ,n224);
    xnor g400(n2667 ,n1[98] ,n1550);
    xor g401(n7103 ,n0[43] ,n0[11]);
    nand g402(n7124 ,n6691 ,n6728);
    nand g403(n3734 ,n6820 ,n3140);
    nor g404(n2376 ,n0[118] ,n1956);
    nand g405(n1102 ,n0[77] ,n792);
    nor g406(n4461 ,n3895 ,n4183);
    xnor g407(n6283 ,n5938 ,n6171);
    xnor g408(n1657 ,n6879 ,n6877);
    not g409(n5775 ,n5774);
    nor g410(n6598 ,n0[121] ,n0[89]);
    nor g411(n3125 ,n1[32] ,n2598);
    or g412(n4848 ,n6 ,n4677);
    nor g413(n4854 ,n6 ,n4682);
    nand g414(n6574 ,n2997 ,n6564);
    nand g415(n5144 ,n6827 ,n4913);
    nand g416(n5098 ,n1955 ,n4991);
    nand g417(n4948 ,n3314 ,n4735);
    xnor g418(n1614 ,n0[89] ,n1[89]);
    xnor g419(n1638 ,n0[6] ,n1[6]);
    nand g420(n2617 ,n742 ,n707);
    nor g421(n5909 ,n5753 ,n5816);
    nand g422(n58 ,n7060 ,n0[4]);
    nor g423(n2997 ,n2204 ,n2203);
    nand g424(n7011 ,n6624 ,n7162);
    nand g425(n264 ,n179 ,n263);
    xnor g426(n6839 ,n86 ,n105);
    xnor g427(n1503 ,n1[50] ,n1[18]);
    nand g428(n2611 ,n890 ,n1825);
    or g429(n9[92] ,n4514 ,n5884);
    xnor g430(n2690 ,n1[105] ,n1574);
    nand g431(n7071 ,n669 ,n639);
    nor g432(n4040 ,n3751 ,n3012);
    nand g433(n1855 ,n0[26] ,n1025);
    xnor g434(n1421 ,n1[48] ,n2[48]);
    nor g435(n4666 ,n2155 ,n4470);
    nor g436(n4043 ,n3758 ,n3032);
    nor g437(n4182 ,n2550 ,n3862);
    xnor g438(n5988 ,n5836 ,n5527);
    nand g439(n5411 ,n717 ,n5270);
    nor g440(n858 ,n791 ,n0[14]);
    nor g441(n5223 ,n713 ,n5060);
    nor g442(n3925 ,n2560 ,n3497);
    nand g443(n2612 ,n750 ,n707);
    nor g444(n6026 ,n5543 ,n5921);
    nand g445(n6356 ,n6274 ,n6273);
    not g446(n6426 ,n6408);
    xnor g447(n1325 ,n0[52] ,n0[36]);
    nor g448(n2608 ,n725 ,n1920);
    nor g449(n6562 ,n5823 ,n6539);
    xnor g450(n1466 ,n1[106] ,n2[42]);
    nand g451(n3696 ,n2238 ,n3161);
    nand g452(n5183 ,n798 ,n4906);
    nor g453(n1049 ,n709 ,n0[7]);
    nand g454(n284 ,n174 ,n283);
    nand g455(n131 ,n50 ,n130);
    nor g456(n3081 ,n1221 ,n2356);
    nor g457(n3466 ,n6823 ,n2818);
    nor g458(n6603 ,n0[126] ,n0[94]);
    xnor g459(n6419 ,n6309 ,n6141);
    xnor g460(n6200 ,n5972 ,n6105);
    nor g461(n4648 ,n715 ,n4475);
    xnor g462(n1596 ,n0[33] ,n1[33]);
    xnor g463(n1667 ,n6834 ,n6835);
    nand g464(n5541 ,n4829 ,n5360);
    not g465(n3493 ,n3492);
    nand g466(n3735 ,n2644 ,n3233);
    nor g467(n5914 ,n5555 ,n5806);
    nor g468(n6708 ,n6826 ,n6585);
    xnor g469(n2848 ,n1315 ,n1657);
    xnor g470(n1293 ,n1[39] ,n4[31]);
    xnor g471(n1502 ,n0[118] ,n0[102]);
    nand g472(n3154 ,n1[87] ,n2346);
    nand g473(n282 ,n191 ,n281);
    nor g474(n3473 ,n1222 ,n2815);
    nor g475(n5349 ,n4718 ,n5194);
    nand g476(n6118 ,n1955 ,n6066);
    xnor g477(n226 ,n1[53] ,n0[53]);
    nand g478(n1111 ,n6876 ,n795);
    not g479(n1562 ,n1561);
    nor g480(n4567 ,n722 ,n4217);
    nand g481(n636 ,n0[94] ,n622);
    xnor g482(n1337 ,n6847 ,n6845);
    nor g483(n2041 ,n1017 ,n1732);
    nand g484(n5031 ,n717 ,n4999);
    nor g485(n2101 ,n954 ,n1962);
    nand g486(n9[116] ,n5868 ,n6103);
    xnor g487(n4905 ,n2841 ,n4465);
    nand g488(n3094 ,n1220 ,n2357);
    xnor g489(n2873 ,n1675 ,n1597);
    nand g490(n1804 ,n0[15] ,n1221);
    or g491(n4037 ,n2553 ,n3391);
    xnor g492(n6850 ,n241 ,n263);
    nand g493(n6054 ,n5895 ,n5977);
    nor g494(n3008 ,n2231 ,n2229);
    xnor g495(n4877 ,n4572 ,n4586);
    xnor g496(n2832 ,n0[119] ,n1263);
    xnor g497(n1495 ,n1[45] ,n1[13]);
    nand g498(n1981 ,n1081 ,n1066);
    nor g499(n2783 ,n1020 ,n2085);
    nand g500(n3673 ,n1953 ,n2945);
    nor g501(n6727 ,n6826 ,n6603);
    nand g502(n5762 ,n4698 ,n5656);
    nor g503(n2181 ,n1962 ,n1396);
    nand g504(n3784 ,n6817 ,n3237);
    nor g505(n853 ,n0[75] ,n0[74]);
    nor g506(n4488 ,n3772 ,n4152);
    xnor g507(n6861 ,n396 ,n421);
    nor g508(n3906 ,n3753 ,n3502);
    nand g509(n1990 ,n1237 ,n1072);
    or g510(n40 ,n7062 ,n0[6]);
    nor g511(n4374 ,n4293 ,n4283);
    nand g512(n6178 ,n1953 ,n6121);
    nand g513(n3773 ,n1117 ,n2753);
    nand g514(n5192 ,n4244 ,n4855);
    nand g515(n3976 ,n748 ,n3571);
    not g516(n4681 ,n4680);
    or g517(n891 ,n743 ,n0[41]);
    nand g518(n4608 ,n717 ,n4430);
    nor g519(n3692 ,n773 ,n3091);
    xnor g520(n6910 ,n225 ,n293);
    nor g521(n2295 ,n1958 ,n1623);
    nand g522(n6690 ,n0[108] ,n0[76]);
    xnor g523(n1922 ,n0[81] ,n1[81]);
    nor g524(n4036 ,n3725 ,n3387);
    xnor g525(n239 ,n1[35] ,n0[35]);
    or g526(n6052 ,n5894 ,n5975);
    nand g527(n6955 ,n6756 ,n6787);
    nand g528(n1903 ,n0[122] ,n999);
    nand g529(n4352 ,n3981 ,n3628);
    nor g530(n2126 ,n1958 ,n1598);
    xnor g531(n1411 ,n1[37] ,n2[37]);
    xnor g532(n2859 ,n1663 ,n1605);
    xor g533(n3826 ,n2662 ,n1[75]);
    xnor g534(n1385 ,n1[56] ,n2[56]);
    nor g535(n2226 ,n1963 ,n1492);
    nand g536(n1092 ,n0[86] ,n789);
    nor g537(n2287 ,n719 ,n1619);
    xnor g538(n81 ,n0[28] ,n7084);
    xnor g539(n1627 ,n0[127] ,n1[127]);
    nor g540(n3856 ,n2556 ,n3715);
    nand g541(n3223 ,n1200 ,n2298);
    nor g542(n5451 ,n4654 ,n5386);
    xnor g543(n3828 ,n1[83] ,n2692);
    nand g544(n3117 ,n763 ,n2586);
    xnor g545(n5203 ,n4431 ,n4837);
    nand g546(n6412 ,n5542 ,n6331);
    xnor g547(n5941 ,n1356 ,n5771);
    nor g548(n6146 ,n5889 ,n6074);
    nor g549(n3364 ,n1954 ,n2906);
    xnor g550(n1265 ,n6830 ,n6829);
    nor g551(n2043 ,n1026 ,n1762);
    nand g552(n4103 ,n3436 ,n3561);
    nor g553(n2352 ,n721 ,n1551);
    nand g554(n2521 ,n794 ,n1979);
    not g555(n2588 ,n2587);
    nand g556(n1774 ,n714 ,n889);
    nor g557(n5949 ,n1954 ,n5854);
    nor g558(n2210 ,n896 ,n1734);
    nand g559(n10[25] ,n4622 ,n5322);
    nand g560(n665 ,n1[27] ,n621);
    nand g561(n7030 ,n6634 ,n7143);
    or g562(n6558 ,n5168 ,n6526);
    xnor g563(n1436 ,n1[88] ,n2[24]);
    xnor g564(n4458 ,n2833 ,n3949);
    nor g565(n3909 ,n6 ,n3494);
    not g566(n751 ,n0[40]);
    nand g567(n6748 ,n0[35] ,n6737);
    nand g568(n4431 ,n2078 ,n4229);
    or g569(n2192 ,n1960 ,n1432);
    nor g570(n3356 ,n1954 ,n2904);
    nor g571(n3066 ,n1827 ,n2318);
    not g572(n5280 ,n5279);
    nor g573(n3311 ,n1[35] ,n3145);
    nor g574(n5614 ,n5481 ,n5395);
    nand g575(n5100 ,n717 ,n4988);
    nor g576(n929 ,n819 ,n0[8]);
    nand g577(n1094 ,n0[61] ,n791);
    nor g578(n6734 ,n7090 ,n7091);
    nor g579(n6236 ,n3553 ,n6129);
    nand g580(n6076 ,n5601 ,n5980);
    nor g581(n5862 ,n713 ,n5845);
    nor g582(n6599 ,n0[122] ,n0[90]);
    nand g583(n4368 ,n3998 ,n4074);
    xnor g584(n1560 ,n0[56] ,n4[16]);
    nor g585(n2418 ,n803 ,n1753);
    not g586(n4365 ,n4364);
    nand g587(n5515 ,n2896 ,n5282);
    nand g588(n3682 ,n1[34] ,n2715);
    nand g589(n1815 ,n809 ,n989);
    not g590(n788 ,n709);
    or g591(n5303 ,n4324 ,n5030);
    nor g592(n3016 ,n2420 ,n2258);
    nor g593(n3141 ,n1817 ,n2575);
    nand g594(n6798 ,n1[103] ,n7088);
    nand g595(n1172 ,n6849 ,n795);
    nand g596(n364 ,n7024 ,n6992);
    nor g597(n1844 ,n0[99] ,n1044);
    nor g598(n4934 ,n3508 ,n4612);
    nand g599(n1809 ,n740 ,n986);
    xnor g600(n6932 ,n535 ,n609);
    or g601(n326 ,n7033 ,n7001);
    xnor g602(n2671 ,n1647 ,n1617);
    not g603(n717 ,n706);
    nand g604(n409 ,n355 ,n408);
    nand g605(n4830 ,n1966 ,n4432);
    not g606(n5065 ,n5064);
    not g607(n5780 ,n5779);
    xnor g608(n4437 ,n2842 ,n3956);
    nand g609(n3722 ,n1114 ,n3047);
    xnor g610(n1470 ,n1[118] ,n2[54]);
    xnor g611(n2900 ,n1710 ,n1543);
    nand g612(n3596 ,n1[63] ,n3006);
    nor g613(n4031 ,n3767 ,n3042);
    xnor g614(n1305 ,n6985 ,n6952);
    not g615(n5273 ,n5272);
    xnor g616(n5771 ,n4874 ,n5457);
    nand g617(n198 ,n0[54] ,n1[54]);
    xnor g618(n2802 ,n0[91] ,n1321);
    xnor g619(n530 ,n6974 ,n0[117]);
    nand g620(n6816 ,n6581 ,n7098);
    nand g621(n1122 ,n6943 ,n795);
    nand g622(n7161 ,n6581 ,n7118);
    nor g623(n2466 ,n1961 ,n1417);
    nand g624(n1870 ,n0[85] ,n964);
    nand g625(n5691 ,n5500 ,n5499);
    nor g626(n4050 ,n3754 ,n3572);
    nor g627(n3321 ,n1954 ,n2885);
    xnor g628(n2821 ,n1256 ,n1696);
    nand g629(n2457 ,n0[0] ,n1765);
    nor g630(n2414 ,n0[41] ,n1758);
    xnor g631(n1322 ,n6846 ,n6844);
    nand g632(n3155 ,n2574 ,n2431);
    nor g633(n5321 ,n4628 ,n5087);
    not g634(n4826 ,n4825);
    nand g635(n4274 ,n2163 ,n3975);
    xnor g636(n5953 ,n697 ,n1581);
    nand g637(n4126 ,n2560 ,n3947);
    nand g638(n267 ,n212 ,n266);
    xnor g639(n1334 ,n7095 ,n7053);
    nand g640(n5288 ,n4687 ,n5088);
    nor g641(n878 ,n756 ,n710);
    nand g642(n6644 ,n0[84] ,n6579);
    nor g643(n951 ,n757 ,n0[65]);
    xor g644(n4923 ,n4445 ,n2801);
    xnor g645(n2803 ,n0[110] ,n1320);
    nand g646(n2589 ,n0[25] ,n1964);
    or g647(n5694 ,n722 ,n5528);
    nor g648(n5703 ,n3533 ,n5511);
    nor g649(n5635 ,n5193 ,n5401);
    xnor g650(n3955 ,n2814 ,n2800);
    not g651(n5538 ,n5537);
    nor g652(n1888 ,n835 ,n11);
    nor g653(n4597 ,n6 ,n4456);
    nand g654(n4800 ,n4072 ,n4533);
    xnor g655(n1701 ,n6855 ,n6853);
    nand g656(n4240 ,n1966 ,n3942);
    xnor g657(n2812 ,n1268 ,n1714);
    nor g658(n2137 ,n1961 ,n1442);
    nand g659(n4565 ,n1173 ,n4126);
    nand g660(n519 ,n0[104] ,n6961);
    nand g661(n4233 ,n3111 ,n3976);
    xor g662(n6835 ,n85 ,n72);
    nand g663(n4379 ,n788 ,n4235);
    nand g664(n4560 ,n1145 ,n4261);
    nor g665(n5376 ,n3877 ,n5044);
    nor g666(n4697 ,n712 ,n4425);
    nand g667(n7144 ,n6630 ,n6708);
    nand g668(n6451 ,n6098 ,n6338);
    not g669(n778 ,n0[54]);
    nand g670(n1219 ,n6828 ,n796);
    not g671(n5484 ,n5483);
    nand g672(n435 ,n354 ,n434);
    nor g673(n2076 ,n1960 ,n1914);
    nor g674(n3895 ,n708 ,n3517);
    nand g675(n1077 ,n0[124] ,n787);
    nand g676(n5401 ,n5213 ,n5221);
    nand g677(n205 ,n0[47] ,n1[47]);
    nand g678(n1982 ,n1236 ,n1105);
    nor g679(n2279 ,n1961 ,n1393);
    nand g680(n6656 ,n1[84] ,n6579);
    not g681(n5165 ,n5164);
    xnor g682(n1916 ,n0[80] ,n1[80]);
    not g683(n5092 ,n5091);
    nor g684(n953 ,n0[53] ,n6);
    not g685(n4824 ,n4823);
    nor g686(n5370 ,n3707 ,n5033);
    nor g687(n5175 ,n6824 ,n4900);
    nor g688(n5109 ,n4971 ,n4814);
    nand g689(n576 ,n487 ,n575);
    nor g690(n3352 ,n2369 ,n3129);
    nand g691(n121 ,n66 ,n120);
    xnor g692(n5768 ,n5392 ,n1357);
    nand g693(n1132 ,n6879 ,n797);
    nand g694(n2989 ,n11 ,n2363);
    nor g695(n4223 ,n4070 ,n3868);
    nand g696(n49 ,n7083 ,n0[27]);
    or g697(n32 ,n7059 ,n0[3]);
    nor g698(n4732 ,n3516 ,n4530);
    nand g699(n217 ,n0[52] ,n1[52]);
    nor g700(n3431 ,n1954 ,n2931);
    nor g701(n4968 ,n981 ,n4797);
    nor g702(n4041 ,n3752 ,n3019);
    nand g703(n1236 ,n0[71] ,n789);
    or g704(n35 ,n7063 ,n0[7]);
    xnor g705(n2670 ,n1324 ,n1546);
    nor g706(n6396 ,n5473 ,n6376);
    or g707(n6238 ,n5704 ,n6166);
    nand g708(n4735 ,n717 ,n4580);
    nand g709(n314 ,n177 ,n313);
    xnor g710(n2834 ,n0[68] ,n1300);
    nor g711(n6291 ,n6047 ,n6238);
    xnor g712(n3829 ,n1[80] ,n2689);
    nand g713(n7139 ,n6679 ,n6729);
    nand g714(n7021 ,n6671 ,n7152);
    xnor g715(n6316 ,n6175 ,n1304);
    nor g716(n945 ,n0[101] ,n715);
    nand g717(n600 ,n486 ,n599);
    xnor g718(n2839 ,n1282 ,n1329);
    nand g719(n4326 ,n2326 ,n4105);
    nor g720(n2260 ,n6 ,n1731);
    nand g721(n2580 ,n0[9] ,n707);
    xnor g722(n2934 ,n1592 ,n1546);
    not g723(n4907 ,n4906);
    nand g724(n369 ,n7038 ,n7006);
    xnor g725(n6210 ,n6068 ,n5838);
    or g726(n2255 ,n1962 ,n1408);
    nand g727(n6984 ,n6757 ,n6788);
    nand g728(n6166 ,n4535 ,n6046);
    nand g729(n7141 ,n6638 ,n6711);
    or g730(n4725 ,n713 ,n4574);
    xnor g731(n401 ,n6999 ,n7031);
    or g732(n3309 ,n1954 ,n2880);
    nand g733(n6032 ,n4656 ,n5888);
    nand g734(n368 ,n7037 ,n7005);
    nor g735(n2719 ,n1735 ,n2442);
    xnor g736(n5072 ,n4659 ,n4666);
    nand g737(n4889 ,n1955 ,n4659);
    nand g738(n413 ,n373 ,n412);
    nand g739(n7143 ,n6690 ,n6709);
    xnor g740(n5945 ,n5839 ,n1548);
    nand g741(n1895 ,n0[60] ,n1221);
    nand g742(n4430 ,n2114 ,n4215);
    xnor g743(n553 ,n6966 ,n0[109]);
    xnor g744(n2892 ,n1292 ,n1685);
    xnor g745(n4920 ,n2807 ,n4443);
    nand g746(n6025 ,n3292 ,n5892);
    nand g747(n5919 ,n4420 ,n5809);
    xnor g748(n6349 ,n5934 ,n6244);
    or g749(n3283 ,n2404 ,n2796);
    nand g750(n7151 ,n6610 ,n6713);
    nor g751(n3252 ,n979 ,n2590);
    nand g752(n6459 ,n6372 ,n6281);
    nor g753(n3273 ,n1954 ,n2923);
    nand g754(n1988 ,n1073 ,n1065);
    or g755(n2063 ,n719 ,n1605);
    nand g756(n1216 ,n1[7] ,n2[7]);
    nand g757(n3771 ,n1110 ,n2777);
    nor g758(n2197 ,n1959 ,n1425);
    nor g759(n4983 ,n6 ,n4810);
    nand g760(n5674 ,n4188 ,n5546);
    nor g761(n3369 ,n1954 ,n2909);
    nand g762(n5708 ,n5515 ,n5523);
    nor g763(n3808 ,n6825 ,n2801);
    nor g764(n2110 ,n1962 ,n1409);
    nor g765(n2276 ,n1001 ,n1997);
    or g766(n190 ,n0[55] ,n1[55]);
    nand g767(n5816 ,n4977 ,n5624);
    nand g768(n6650 ,n1[82] ,n6580);
    xnor g769(n1346 ,n0[126] ,n4[14]);
    nand g770(n6470 ,n6400 ,n6399);
    nor g771(n4188 ,n4079 ,n3788);
    not g772(n766 ,n0[123]);
    nor g773(n5177 ,n6824 ,n4904);
    nor g774(n5188 ,n706 ,n4992);
    nand g775(n983 ,n714 ,n734);
    xor g776(n3834 ,n2690 ,n1[73]);
    nand g777(n4330 ,n2586 ,n3912);
    xnor g778(n1438 ,n1[72] ,n2[8]);
    nand g779(n7125 ,n6687 ,n6727);
    nand g780(n7135 ,n6655 ,n6717);
    xnor g781(n1689 ,n0[107] ,n4[3]);
    xnor g782(n6869 ,n398 ,n425);
    nand g783(n1084 ,n0[54] ,n794);
    xnor g784(n2918 ,n1344 ,n1628);
    nor g785(n6089 ,n3476 ,n5961);
    xnor g786(n6923 ,n76 ,n147);
    nor g787(n5025 ,n4689 ,n4877);
    xnor g788(n6045 ,n5847 ,n4584);
    nor g789(n2924 ,n1866 ,n2610);
    nor g790(n1787 ,n0[80] ,n1023);
    nand g791(n4547 ,n1188 ,n4133);
    nor g792(n5646 ,n5254 ,n5475);
    not g793(n5096 ,n5095);
    nor g794(n947 ,n758 ,n0[34]);
    nor g795(n5365 ,n3500 ,n5147);
    xnor g796(n548 ,n6961 ,n0[104]);
    xnor g797(n1376 ,n0[72] ,n7100);
    xnor g798(n5983 ,n5837 ,n5269);
    nand g799(n4059 ,n2763 ,n3656);
    nand g800(n315 ,n214 ,n314);
    xnor g801(n1254 ,n6857 ,n6856);
    xnor g802(n90 ,n0[6] ,n7062);
    nand g803(n6795 ,n1[102] ,n7088);
    or g804(n324 ,n7034 ,n7002);
    nor g805(n5148 ,n727 ,n4921);
    or g806(n6472 ,n6406 ,n6346);
    xnor g807(n6882 ,n249 ,n279);
    nand g808(n662 ,n1[11] ,n621);
    xnor g809(n1711 ,n0[113] ,n4[1]);
    nand g810(n4607 ,n717 ,n4570);
    nand g811(n852 ,n0[17] ,n742);
    not g812(n800 ,n0[122]);
    nand g813(n6075 ,n5685 ,n5975);
    nand g814(n1974 ,n1070 ,n930);
    xnor g815(n3811 ,n2647 ,n1969);
    nor g816(n5300 ,n3317 ,n5038);
    nand g817(n1765 ,n723 ,n1028);
    not g818(n2027 ,n2026);
    nor g819(n2227 ,n719 ,n1583);
    or g820(n5955 ,n712 ,n5938);
    not g821(n1995 ,n1994);
    nand g822(n3797 ,n2481 ,n2785);
    xnor g823(n2869 ,n1290 ,n1687);
    nand g824(n3201 ,n765 ,n2534);
    xnor g825(n1564 ,n0[117] ,n0[101]);
    xnor g826(n3842 ,n1[94] ,n2655);
    nor g827(n2766 ,n1498 ,n2614);
    nand g828(n4114 ,n3110 ,n3315);
    nand g829(n6402 ,n3399 ,n702);
    nand g830(n1076 ,n0[29] ,n715);
    nand g831(n410 ,n332 ,n409);
    nor g832(n3532 ,n6825 ,n2844);
    nand g833(n291 ,n211 ,n290);
    nand g834(n4383 ,n4196 ,n4020);
    nand g835(n1009 ,n0[122] ,n714);
    nand g836(n3396 ,n2220 ,n2750);
    or g837(n342 ,n7041 ,n7009);
    or g838(n2995 ,n1[57] ,n2589);
    nor g839(n5318 ,n4739 ,n5180);
    xnor g840(n1538 ,n0[17] ,n1[17]);
    nand g841(n3358 ,n1953 ,n2878);
    or g842(n2764 ,n1566 ,n2617);
    xnor g843(n6860 ,n548 ,n573);
    nand g844(n3180 ,n1986 ,n2326);
    xnor g845(n554 ,n6967 ,n0[110]);
    not g846(n710 ,n715);
    nand g847(n3392 ,n2087 ,n2764);
    xnor g848(n6939 ,n80 ,n155);
    nand g849(n6445 ,n6090 ,n6336);
    nand g850(n1992 ,n820 ,n990);
    nor g851(n3865 ,n969 ,n3291);
    nor g852(n4086 ,n791 ,n3791);
    xnor g853(n5195 ,n4990 ,n1350);
    nor g854(n3420 ,n1222 ,n2841);
    xnor g855(n1363 ,n0[11] ,n4[27]);
    xnor g856(n4370 ,n4102 ,n3950);
    xnor g857(n7055 ,n84 ,n163);
    xnor g858(n254 ,n1[50] ,n0[50]);
    or g859(n6158 ,n3475 ,n6041);
    xnor g860(n6905 ,n407 ,n443);
    nand g861(n2450 ,n990 ,n1784);
    nor g862(n5141 ,n727 ,n4909);
    xnor g863(n539 ,n6983 ,n0[126]);
    nor g864(n6473 ,n6368 ,n6461);
    or g865(n5748 ,n711 ,n5639);
    nand g866(n3218 ,n1121 ,n2046);
    xnor g867(n1317 ,n0[35] ,n1[51]);
    nand g868(n7126 ,n6685 ,n6726);
    not g869(n737 ,n0[24]);
    nor g870(n5428 ,n5099 ,n5265);
    nand g871(n678 ,n1[3] ,n621);
    nand g872(n1182 ,n6895 ,n797);
    or g873(n3898 ,n2332 ,n3490);
    nand g874(n2601 ,n0[18] ,n707);
    nand g875(n5002 ,n2509 ,n4674);
    nor g876(n1753 ,n724 ,n881);
    or g877(n2469 ,n830 ,n1485);
    xnor g878(n2952 ,n1700 ,n1610);
    nand g879(n5715 ,n4804 ,n5488);
    or g880(n5523 ,n2896 ,n5283);
    nand g881(n2483 ,n1244 ,n1992);
    xnor g882(n4915 ,n2818 ,n4439);
    xnor g883(n5453 ,n4570 ,n5158);
    nand g884(n10[21] ,n4762 ,n5341);
    or g885(n479 ,n0[109] ,n6966);
    xnor g886(n6920 ,n532 ,n603);
    nor g887(n5147 ,n727 ,n4919);
    nor g888(n3900 ,n2227 ,n3745);
    xnor g889(n83 ,n0[30] ,n7086);
    nand g890(n4967 ,n3338 ,n4637);
    nand g891(n4333 ,n2582 ,n3893);
    nand g892(n3078 ,n11 ,n2389);
    nor g893(n956 ,n815 ,n791);
    nor g894(n6501 ,n6380 ,n6420);
    nand g895(n3746 ,n7155 ,n3100);
    nand g896(n2491 ,n0[51] ,n1786);
    xnor g897(n5219 ,n4877 ,n2668);
    nand g898(n4125 ,n2560 ,n3948);
    xnor g899(n6874 ,n247 ,n275);
    xnor g900(n97 ,n0[13] ,n7069);
    xnor g901(n74 ,n0[21] ,n7077);
    not g902(n1031 ,n1030);
    nand g903(n656 ,n1[29] ,n621);
    xor g904(n5276 ,n4660 ,n5003);
    nor g905(n3659 ,n805 ,n3090);
    nor g906(n3257 ,n2012 ,n2611);
    nand g907(n3557 ,n789 ,n2916);
    nor g908(n3524 ,n6825 ,n2835);
    nand g909(n4361 ,n2018 ,n3844);
    nor g910(n5312 ,n3420 ,n5180);
    nor g911(n5951 ,n712 ,n5939);
    nand g912(n4574 ,n2521 ,n4229);
    nor g913(n5393 ,n2325 ,n5380);
    nand g914(n6277 ,n6148 ,n6219);
    nor g915(n720 ,n7091 ,n1240);
    nand g916(n4002 ,n0[94] ,n3490);
    not g917(n4100 ,n4099);
    not g918(n2630 ,n2629);
    not g919(n4921 ,n4920);
    nand g920(n4019 ,n789 ,n3799);
    xnor g921(n5260 ,n4999 ,n5003);
    nand g922(n4087 ,n6808 ,n3648);
    not g923(n4107 ,n4106);
    or g924(n343 ,n7032 ,n7000);
    nand g925(n7070 ,n667 ,n637);
    not g926(n723 ,n724);
    or g927(n334 ,n7039 ,n7007);
    nor g928(n6261 ,n713 ,n6244);
    nand g929(n7003 ,n6700 ,n6805);
    xnor g930(n3821 ,n1[66] ,n2667);
    nand g931(n219 ,n0[57] ,n1[57]);
    nand g932(n4791 ,n2326 ,n4587);
    nor g933(n3004 ,n1[62] ,n2571);
    xnor g934(n6916 ,n531 ,n601);
    nand g935(n3631 ,n0[63] ,n2794);
    nor g936(n2622 ,n0[26] ,n1963);
    xnor g937(n5944 ,n4[2] ,n5837);
    xnor g938(n1659 ,n6930 ,n6931);
    nor g939(n2406 ,n0[80] ,n1772);
    nor g940(n2038 ,n1957 ,n1485);
    nand g941(n580 ,n468 ,n579);
    nand g942(n7165 ,n6581 ,n7114);
    xnor g943(n1921 ,n1[116] ,n2[52]);
    nor g944(n3914 ,n2400 ,n3490);
    nor g945(n5688 ,n4788 ,n5556);
    nand g946(n3167 ,n2569 ,n2473);
    xnor g947(n6893 ,n404 ,n437);
    nor g948(n4178 ,n3223 ,n4076);
    xnor g949(n5209 ,n4996 ,n4569);
    nand g950(n449 ,n346 ,n448);
    nor g951(n6060 ,n5659 ,n5977);
    nand g952(n2769 ,n1497 ,n2627);
    nor g953(n2274 ,n1961 ,n1467);
    xnor g954(n1633 ,n0[69] ,n1[69]);
    nor g955(n1033 ,n811 ,n0[1]);
    nand g956(n4587 ,n4253 ,n4256);
    xnor g957(n541 ,n6954 ,n0[97]);
    nand g958(n5406 ,n5097 ,n5260);
    nor g959(n5864 ,n712 ,n5844);
    nand g960(n2604 ,n824 ,n707);
    nor g961(n5516 ,n5170 ,n5262);
    nor g962(n3571 ,n725 ,n3132);
    nor g963(n6719 ,n6826 ,n6595);
    nand g964(n7154 ,n6581 ,n7051);
    or g965(n474 ,n0[124] ,n6981);
    xnor g966(n1663 ,n0[76] ,n4[4]);
    nor g967(n5360 ,n3524 ,n5141);
    nand g968(n459 ,n372 ,n458);
    or g969(n4311 ,n3897 ,n3704);
    nand g970(n3730 ,n3231 ,n3211);
    nand g971(n5001 ,n2251 ,n4673);
    nor g972(n1746 ,n0[99] ,n1002);
    or g973(n6481 ,n6430 ,n6424);
    nor g974(n5818 ,n1954 ,n5590);
    nor g975(n2312 ,n1959 ,n1394);
    nand g976(n69 ,n7059 ,n0[3]);
    xnor g977(n3938 ,n1367 ,n2830);
    or g978(n3873 ,n2403 ,n3490);
    xnor g979(n1375 ,n6901 ,n6900);
    nor g980(n4869 ,n3438 ,n4696);
    nand g981(n1137 ,n6851 ,n795);
    nor g982(n5718 ,n794 ,n5452);
    or g983(n4170 ,n788 ,n4116);
    nor g984(n3383 ,n1[59] ,n3169);
    or g985(n2100 ,n719 ,n1558);
    nor g986(n5496 ,n4972 ,n5288);
    nand g987(n9[8] ,n6365 ,n6473);
    nand g988(n6156 ,n3991 ,n6037);
    or g989(n6442 ,n5163 ,n6367);
    nor g990(n2251 ,n1778 ,n1780);
    xnor g991(n2895 ,n1352 ,n1603);
    or g992(n6480 ,n6373 ,n703);
    nor g993(n2771 ,n2098 ,n2055);
    nand g994(n7032 ,n6640 ,n7141);
    nor g995(n3580 ,n806 ,n2773);
    or g996(n5129 ,n4668 ,n4882);
    nor g997(n2221 ,n1961 ,n1440);
    nand g998(n3756 ,n7126 ,n3116);
    nand g999(n3729 ,n6822 ,n3108);
    nor g1000(n5189 ,n6824 ,n4914);
    xnor g1001(n1390 ,n1[47] ,n2[47]);
    or g1002(n5241 ,n4694 ,n5066);
    nor g1003(n2732 ,n891 ,n2165);
    nor g1004(n2012 ,n803 ,n1229);
    nand g1005(n2566 ,n0[22] ,n1964);
    or g1006(n482 ,n0[118] ,n6975);
    nand g1007(n5093 ,n4242 ,n4959);
    xnor g1008(n6925 ,n381 ,n453);
    nand g1009(n11 ,n3[3] ,n3[2]);
    nand g1010(n5868 ,n717 ,n5729);
    xnor g1011(n1913 ,n0[82] ,n1[82]);
    nand g1012(n3974 ,n968 ,n3803);
    or g1013(n192 ,n0[38] ,n1[38]);
    or g1014(n9[51] ,n4510 ,n6566);
    nor g1015(n2495 ,n778 ,n1958);
    nor g1016(n865 ,n791 ,n0[102]);
    nand g1017(n4485 ,n4278 ,n3874);
    not g1018(n1545 ,n1544);
    xnor g1019(n397 ,n6995 ,n7027);
    nand g1020(n639 ,n0[79] ,n622);
    nand g1021(n3220 ,n1132 ,n2160);
    or g1022(n9[85] ,n5750 ,n5925);
    nand g1023(n5713 ,n5438 ,n4903);
    xnor g1024(n4841 ,n4580 ,n1572);
    nand g1025(n3687 ,n3152 ,n2464);
    nand g1026(n2018 ,n723 ,n1014);
    nand g1027(n4973 ,n4021 ,n4727);
    nand g1028(n10[6] ,n4610 ,n5318);
    xor g1029(n7114 ,n0[54] ,n0[22]);
    xnor g1030(n6336 ,n5935 ,n6245);
    xnor g1031(n4457 ,n2802 ,n3951);
    xnor g1032(n2828 ,n1310 ,n1655);
    nand g1033(n5105 ,n717 ,n5000);
    nand g1034(n4513 ,n3710 ,n4177);
    nand g1035(n448 ,n334 ,n447);
    or g1036(n2762 ,n1493 ,n2620);
    nand g1037(n3189 ,n2010 ,n2157);
    xnor g1038(n5067 ,n4661 ,n4585);
    or g1039(n4720 ,n713 ,n4580);
    nand g1040(n6334 ,n1955 ,n6306);
    nor g1041(n4046 ,n3763 ,n3035);
    nand g1042(n5894 ,n717 ,n5846);
    nor g1043(n6079 ,n5671 ,n5980);
    nand g1044(n5243 ,n4939 ,n5068);
    nor g1045(n5155 ,n2120 ,n4883);
    not g1046(n836 ,n0[118]);
    nor g1047(n3128 ,n1[42] ,n2583);
    nor g1048(n3506 ,n1222 ,n2843);
    nor g1049(n2231 ,n1961 ,n1402);
    nand g1050(n5320 ,n4033 ,n5127);
    nand g1051(n7147 ,n6678 ,n6705);
    xnor g1052(n3848 ,n1[90] ,n2707);
    nor g1053(n849 ,n0[3] ,n0[2]);
    nor g1054(n955 ,n0[46] ,n787);
    nand g1055(n3436 ,n708 ,n3251);
    nor g1056(n5924 ,n5818 ,n5825);
    nand g1057(n2473 ,n0[52] ,n718);
    or g1058(n4055 ,n3652 ,n3506);
    nand g1059(n2539 ,n1115 ,n1889);
    not g1060(n6384 ,n6354);
    nand g1061(n6962 ,n6738 ,n6800);
    nor g1062(n3085 ,n1221 ,n2366);
    nor g1063(n6395 ,n5541 ,n6355);
    nor g1064(n4933 ,n3505 ,n4614);
    nand g1065(n5741 ,n1953 ,n5579);
    xnor g1066(n1930 ,n0[60] ,n1[60]);
    nand g1067(n5412 ,n5284 ,n5282);
    nor g1068(n4710 ,n6824 ,n4478);
    nand g1069(n3219 ,n1175 ,n2192);
    nor g1070(n2388 ,n0[38] ,n1957);
    nand g1071(n2490 ,n805 ,n2007);
    xor g1072(n7052 ,n0[98] ,n0[66]);
    xor g1073(n7123 ,n0[63] ,n0[31]);
    nand g1074(n4874 ,n2058 ,n4679);
    nand g1075(n2165 ,n1010 ,n1737);
    nand g1076(n4112 ,n1901 ,n3297);
    nand g1077(n9[19] ,n5513 ,n6573);
    xnor g1078(n2894 ,n1257 ,n1720);
    nor g1079(n6576 ,n5672 ,n6574);
    nor g1080(n2438 ,n1956 ,n1595);
    xnor g1081(n5452 ,n5019 ,n3248);
    nor g1082(n5437 ,n3296 ,n5287);
    nand g1083(n4338 ,n2573 ,n3916);
    xnor g1084(n2845 ,n1277 ,n1661);
    or g1085(n2086 ,n1962 ,n1452);
    nand g1086(n1799 ,n800 ,n1021);
    nand g1087(n9[123] ,n4413 ,n6571);
    or g1088(n4156 ,n4048 ,n3775);
    nor g1089(n2398 ,n1[119] ,n1958);
    nand g1090(n1100 ,n0[20] ,n709);
    nand g1091(n6392 ,n1952 ,n6316);
    xnor g1092(n5071 ,n4665 ,n4582);
    nand g1093(n3800 ,n921 ,n2731);
    nor g1094(n3522 ,n2414 ,n2729);
    or g1095(n471 ,n0[114] ,n6971);
    xnor g1096(n5777 ,n5268 ,n5462);
    not g1097(n769 ,n0[96]);
    xnor g1098(n2699 ,n1[119] ,n1579);
    nand g1099(n4752 ,n715 ,n4589);
    nor g1100(n5624 ,n5185 ,n5402);
    nand g1101(n676 ,n1[2] ,n621);
    nor g1102(n6488 ,n4398 ,n6442);
    nor g1103(n940 ,n0[18] ,n723);
    nand g1104(n289 ,n200 ,n288);
    nand g1105(n6686 ,n1[93] ,n6580);
    nor g1106(n5118 ,n4329 ,n4847);
    nand g1107(n452 ,n342 ,n451);
    nor g1108(n4959 ,n3536 ,n4775);
    nor g1109(n6474 ,n5387 ,n6444);
    not g1110(n2572 ,n2571);
    nor g1111(n6013 ,n3332 ,n5864);
    or g1112(n497 ,n0[122] ,n6979);
    nand g1113(n6817 ,n6581 ,n7097);
    xnor g1114(n5577 ,n1284 ,n5203);
    nor g1115(n2479 ,n825 ,n721);
    nor g1116(n1189 ,n847 ,n716);
    nor g1117(n5670 ,n6 ,n5529);
    nand g1118(n2344 ,n840 ,n718);
    nor g1119(n3868 ,n787 ,n3793);
    nand g1120(n4685 ,n717 ,n4429);
    nor g1121(n5604 ,n4685 ,n5453);
    nand g1122(n3749 ,n7162 ,n3060);
    or g1123(n2213 ,n1961 ,n1465);
    nand g1124(n7137 ,n6649 ,n6715);
    nor g1125(n2122 ,n719 ,n1930);
    nand g1126(n6738 ,n0[41] ,n6737);
    xnor g1127(n247 ,n1[43] ,n0[43]);
    xnor g1128(n558 ,n6971 ,n0[114]);
    nand g1129(n4153 ,n2326 ,n4109);
    nand g1130(n4242 ,n1966 ,n3948);
    xnor g1131(n1512 ,n1[42] ,n1[10]);
    nor g1132(n2401 ,n0[1] ,n1769);
    or g1133(n3042 ,n2237 ,n2424);
    or g1134(n5117 ,n4068 ,n4976);
    xnor g1135(n5640 ,n5297 ,n4363);
    nor g1136(n2449 ,n854 ,n1962);
    nor g1137(n5934 ,n4194 ,n5774);
    nor g1138(n3472 ,n1954 ,n2942);
    nand g1139(n3203 ,n1201 ,n2057);
    xor g1140(n7111 ,n0[51] ,n0[19]);
    nand g1141(n3698 ,n1[67] ,n2910);
    nor g1142(n4474 ,n2412 ,n4349);
    not g1143(n976 ,n975);
    nand g1144(n263 ,n210 ,n262);
    nand g1145(n9[108] ,n5859 ,n6087);
    or g1146(n4870 ,n3987 ,n4638);
    nor g1147(n2756 ,n2037 ,n2216);
    xnor g1148(n5969 ,n5784 ,n5009);
    nand g1149(n6502 ,n6454 ,n6341);
    nand g1150(n512 ,n0[112] ,n6969);
    xnor g1151(n6414 ,n6311 ,n6310);
    nor g1152(n2179 ,n1957 ,n1596);
    nor g1153(n2039 ,n721 ,n1487);
    nand g1154(n502 ,n0[118] ,n6975);
    nand g1155(n6168 ,n6101 ,n6086);
    nor g1156(n908 ,n808 ,n0[41]);
    or g1157(n318 ,n7022 ,n6990);
    nor g1158(n5497 ,n5320 ,n5290);
    nor g1159(n4559 ,n1168 ,n4263);
    nand g1160(n10[11] ,n4770 ,n5347);
    nor g1161(n1166 ,n848 ,n716);
    nand g1162(n5185 ,n4238 ,n4858);
    nand g1163(n3258 ,n948 ,n2031);
    nand g1164(n3191 ,n809 ,n2529);
    xnor g1165(n4913 ,n2848 ,n4436);
    xnor g1166(n6948 ,n539 ,n617);
    nor g1167(n1997 ,n0[112] ,n978);
    xnor g1168(n1356 ,n0[124] ,n4[12]);
    nor g1169(n2150 ,n1956 ,n1628);
    nand g1170(n653 ,n0[70] ,n622);
    nor g1171(n5809 ,n5721 ,n5557);
    nand g1172(n47 ,n7069 ,n0[13]);
    nand g1173(n2107 ,n978 ,n1743);
    nand g1174(n6223 ,n3326 ,n6130);
    nand g1175(n148 ,n38 ,n147);
    nor g1176(n3368 ,n1954 ,n2908);
    nor g1177(n4144 ,n709 ,n4115);
    nand g1178(n598 ,n472 ,n597);
    nand g1179(n3105 ,n1806 ,n2049);
    nor g1180(n854 ,n1[55] ,n2[55]);
    nand g1181(n3595 ,n0[57] ,n3022);
    nand g1182(n6784 ,n1[96] ,n7088);
    nand g1183(n1204 ,n6928 ,n795);
    nand g1184(n365 ,n7025 ,n6993);
    nand g1185(n6975 ,n6739 ,n6786);
    xnor g1186(n1360 ,n1[22] ,n4[22]);
    nor g1187(n5554 ,n4826 ,n5369);
    nand g1188(n297 ,n194 ,n296);
    xnor g1189(n2885 ,n1364 ,n1616);
    nand g1190(n6294 ,n6161 ,n6207);
    not g1191(n1242 ,n1241);
    nor g1192(n1752 ,n0[56] ,n992);
    nor g1193(n6280 ,n4853 ,n6192);
    nand g1194(n4359 ,n4052 ,n3883);
    xnor g1195(n6187 ,n6033 ,n6035);
    nand g1196(n7159 ,n6581 ,n7120);
    nor g1197(n990 ,n725 ,n0[67]);
    nand g1198(n9[72] ,n5489 ,n6533);
    xnor g1199(n3917 ,n1[84] ,n2694);
    xnor g1200(n2793 ,n1643 ,n1582);
    not g1201(n847 ,n6904);
    nand g1202(n5548 ,n4819 ,n5365);
    xnor g1203(n1587 ,n0[36] ,n0[20]);
    xnor g1204(n1528 ,n1[57] ,n1[25]);
    not g1205(n5088 ,n5087);
    nand g1206(n4256 ,n715 ,n3964);
    nand g1207(n7074 ,n680 ,n649);
    or g1208(n2417 ,n0[113] ,n1770);
    nor g1209(n6249 ,n4641 ,n6142);
    not g1210(n4668 ,n4667);
    nand g1211(n3629 ,n0[60] ,n2794);
    xnor g1212(n1431 ,n1[25] ,n2[25]);
    nand g1213(n361 ,n7020 ,n6988);
    nand g1214(n5531 ,n4396 ,n5327);
    nor g1215(n6309 ,n4983 ,n6194);
    nor g1216(n3492 ,n2410 ,n2733);
    or g1217(n3033 ,n2312 ,n2309);
    nand g1218(n5355 ,n3463 ,n5066);
    nor g1219(n5347 ,n4716 ,n5160);
    xnor g1220(n6921 ,n380 ,n451);
    xnor g1221(n6114 ,n5843 ,n5944);
    nand g1222(n432 ,n327 ,n431);
    xnor g1223(n3833 ,n1[77] ,n2673);
    nand g1224(n9[79] ,n4341 ,n5914);
    nand g1225(n272 ,n183 ,n271);
    nand g1226(n9[21] ,n5427 ,n5924);
    xnor g1227(n79 ,n0[26] ,n7082);
    nand g1228(n884 ,n0[122] ,n725);
    nor g1229(n4481 ,n2977 ,n4296);
    or g1230(n3036 ,n2171 ,n2485);
    nor g1231(n6001 ,n3406 ,n5873);
    nand g1232(n2564 ,n0[29] ,n707);
    or g1233(n4196 ,n722 ,n4103);
    nand g1234(n2750 ,n1540 ,n2634);
    nand g1235(n626 ,n0[72] ,n622);
    or g1236(n9[48] ,n3969 ,n6561);
    nand g1237(n163 ,n62 ,n162);
    not g1238(n756 ,n0[22]);
    nand g1239(n2502 ,n1867 ,n1831);
    xnor g1240(n1695 ,n6891 ,n6889);
    nor g1241(n898 ,n0[92] ,n790);
    nor g1242(n2270 ,n1959 ,n1395);
    nor g1243(n4963 ,n985 ,n4782);
    xor g1244(n690 ,n4872 ,n2675);
    not g1245(n715 ,n791);
    nand g1246(n6240 ,n4635 ,n6157);
    nor g1247(n5051 ,n713 ,n4873);
    nor g1248(n6260 ,n713 ,n6245);
    nand g1249(n3663 ,n3139 ,n2772);
    nand g1250(n9[13] ,n5950 ,n5908);
    or g1251(n4139 ,n1961 ,n3835);
    nor g1252(n3076 ,n1221 ,n2352);
    xnor g1253(n4837 ,n4430 ,n1296);
    nor g1254(n3738 ,n2540 ,n3264);
    xnor g1255(n5572 ,n1328 ,n5274);
    nor g1256(n3091 ,n1221 ,n2362);
    xnor g1257(n2867 ,n1613 ,n1516);
    nand g1258(n4818 ,n1966 ,n4443);
    nor g1259(n6313 ,n6289 ,n6286);
    nor g1260(n1733 ,n0[72] ,n982);
    xnor g1261(n4434 ,n2830 ,n3958);
    xnor g1262(n251 ,n1[47] ,n0[47]);
    nand g1263(n1177 ,n6885 ,n797);
    nor g1264(n5358 ,n3513 ,n5139);
    nor g1265(n3086 ,n1221 ,n2358);
    xnor g1266(n4906 ,n2843 ,n4432);
    nor g1267(n1769 ,n724 ,n1020);
    not g1268(n724 ,n7);
    nor g1269(n4667 ,n2149 ,n4472);
    nor g1270(n2246 ,n1962 ,n1431);
    nand g1271(n3640 ,n1[58] ,n2999);
    xnor g1272(n5245 ,n4835 ,n4842);
    not g1273(n781 ,n1[58]);
    xnor g1274(n2856 ,n1333 ,n1526);
    nor g1275(n6368 ,n5992 ,n6281);
    nor g1276(n5160 ,n6824 ,n4912);
    xnor g1277(n1268 ,n6893 ,n6892);
    xnor g1278(n1361 ,n0[38] ,n0[22]);
    nor g1279(n2391 ,n721 ,n1497);
    nand g1280(n4810 ,n4381 ,n4201);
    or g1281(n3000 ,n1227 ,n2611);
    nand g1282(n3985 ,n787 ,n3511);
    xnor g1283(n6862 ,n244 ,n269);
    nor g1284(n4867 ,n4146 ,n4710);
    nand g1285(n9[87] ,n4794 ,n5916);
    or g1286(n5686 ,n4935 ,n5469);
    nor g1287(n3299 ,n1954 ,n2859);
    nand g1288(n4566 ,n7132 ,n4132);
    nor g1289(n4145 ,n1960 ,n3842);
    nor g1290(n5742 ,n5600 ,n5599);
    nand g1291(n5992 ,n717 ,n5931);
    nand g1292(n1067 ,n0[33] ,n714);
    nand g1293(n3139 ,n1535 ,n2563);
    not g1294(n4995 ,n4996);
    nand g1295(n4503 ,n3695 ,n4182);
    nand g1296(n2527 ,n792 ,n1967);
    nand g1297(n1124 ,n6861 ,n795);
    nand g1298(n3776 ,n1111 ,n3182);
    nor g1299(n3278 ,n790 ,n3255);
    xnor g1300(n1464 ,n1[99] ,n2[35]);
    nand g1301(n3394 ,n1953 ,n2920);
    nor g1302(n6244 ,n3909 ,n6142);
    nand g1303(n1915 ,n714 ,n1247);
    xnor g1304(n5752 ,n2703 ,n5465);
    nor g1305(n6436 ,n6089 ,n6343);
    or g1306(n4198 ,n3771 ,n4059);
    nor g1307(n6524 ,n5474 ,n6468);
    nand g1308(n9[59] ,n5695 ,n6556);
    not g1309(n821 ,n0[98]);
    nand g1310(n4426 ,n2259 ,n4230);
    nor g1311(n2339 ,n1[116] ,n1957);
    nand g1312(n6462 ,n6093 ,n6349);
    or g1313(n4061 ,n3658 ,n3806);
    or g1314(n2159 ,n1962 ,n1481);
    nor g1315(n3432 ,n788 ,n2925);
    nand g1316(n3661 ,n3138 ,n2306);
    nor g1317(n3162 ,n2584 ,n2470);
    nand g1318(n7149 ,n6637 ,n6703);
    nand g1319(n1008 ,n0[90] ,n714);
    not g1320(n4448 ,n4447);
    or g1321(n9[14] ,n5738 ,n5927);
    or g1322(n3928 ,n2792 ,n3776);
    nor g1323(n3276 ,n1954 ,n2860);
    nor g1324(n6023 ,n3346 ,n5917);
    or g1325(n4252 ,n2325 ,n4104);
    nand g1326(n925 ,n0[114] ,n724);
    or g1327(n3011 ,n2242 ,n2241);
    nand g1328(n6773 ,n1[119] ,n7088);
    nand g1329(n3597 ,n0[100] ,n2794);
    xor g1330(n7115 ,n0[55] ,n0[23]);
    xnor g1331(n3827 ,n1[76] ,n2661);
    nor g1332(n3567 ,n1222 ,n2810);
    not g1333(n4873 ,n4874);
    nor g1334(n5605 ,n706 ,n5512);
    nand g1335(n7056 ,n682 ,n642);
    xnor g1336(n6347 ,n6245 ,n6171);
    nor g1337(n1810 ,n809 ,n11);
    or g1338(n4304 ,n2536 ,n3861);
    xnor g1339(n3949 ,n2806 ,n2852);
    nand g1340(n3686 ,n3151 ,n2169);
    nand g1341(n1985 ,n997 ,n1062);
    nand g1342(n661 ,n1[21] ,n621);
    nor g1343(n1732 ,n1019 ,n851);
    nand g1344(n5527 ,n4318 ,n5273);
    nor g1345(n2083 ,n1960 ,n1406);
    nand g1346(n4089 ,n7148 ,n3429);
    nand g1347(n3320 ,n1953 ,n2883);
    xnor g1348(n1446 ,n1[113] ,n2[49]);
    nand g1349(n3633 ,n1[39] ,n3014);
    xnor g1350(n4836 ,n4427 ,n1563);
    nor g1351(n6586 ,n0[109] ,n0[77]);
    or g1352(n4695 ,n712 ,n4431);
    nor g1353(n4936 ,n3499 ,n4613);
    nand g1354(n5709 ,n5517 ,n5446);
    xnor g1355(n6131 ,n5947 ,n4214);
    nor g1356(n5132 ,n727 ,n4893);
    xnor g1357(n2666 ,n1[100] ,n1498);
    nand g1358(n3439 ,n714 ,n3121);
    nand g1359(n195 ,n0[61] ,n1[61]);
    not g1360(n5995 ,n5994);
    nor g1361(n2293 ,n1956 ,n1637);
    nor g1362(n4943 ,n2325 ,n4810);
    nor g1363(n2371 ,n1[45] ,n1956);
    nand g1364(n2513 ,n1882 ,n1869);
    nand g1365(n4636 ,n717 ,n4428);
    not g1366(n5467 ,n5466);
    nand g1367(n5692 ,n5502 ,n5501);
    nand g1368(n5519 ,n4481 ,n5302);
    xnor g1369(n6915 ,n74 ,n143);
    xnor g1370(n1591 ,n0[91] ,n1[91]);
    nand g1371(n2594 ,n0[24] ,n1964);
    xnor g1372(n1419 ,n1[26] ,n2[26]);
    nor g1373(n3669 ,n1222 ,n2845);
    nand g1374(n617 ,n499 ,n616);
    nand g1375(n2526 ,n794 ,n1970);
    nand g1376(n6806 ,n6581 ,n7108);
    nor g1377(n1027 ,n0[108] ,n790);
    xnor g1378(n6386 ,n0[3] ,n6307);
    nor g1379(n2216 ,n1962 ,n1459);
    xnor g1380(n1547 ,n0[85] ,n4[29]);
    or g1381(n4628 ,n3528 ,n4542);
    xnor g1382(n73 ,n0[20] ,n7076);
    nand g1383(n428 ,n316 ,n427);
    nor g1384(n2178 ,n1959 ,n1900);
    not g1385(n6207 ,n6206);
    or g1386(n29 ,n7085 ,n0[29]);
    nand g1387(n7062 ,n684 ,n653);
    nand g1388(n3097 ,n1514 ,n2600);
    nand g1389(n3762 ,n7137 ,n3066);
    nor g1390(n3533 ,n1222 ,n2807);
    not g1391(n986 ,n985);
    nand g1392(n4321 ,n793 ,n4105);
    xnor g1393(n4843 ,n4568 ,n2686);
    nand g1394(n4808 ,n4372 ,n4257);
    or g1395(n3469 ,n1487 ,n2743);
    or g1396(n495 ,n0[110] ,n6967);
    not g1397(n1961 ,n720);
    nand g1398(n3185 ,n2426 ,n1942);
    nand g1399(n5305 ,n709 ,n5173);
    xor g1400(n7093 ,n0[33] ,n0[1]);
    nand g1401(n3261 ,n897 ,n2480);
    xnor g1402(n2907 ,n1713 ,n1575);
    nor g1403(n3296 ,n1954 ,n2858);
    nand g1404(n3435 ,n788 ,n2963);
    or g1405(n3017 ,n2125 ,n2261);
    nor g1406(n892 ,n733 ,n0[88]);
    nand g1407(n5925 ,n4747 ,n5810);
    xnor g1408(n6918 ,n227 ,n297);
    xnor g1409(n2872 ,n1270 ,n1524);
    not g1410(n2889 ,n2888);
    or g1411(n3923 ,n790 ,n3797);
    not g1412(n6199 ,n6198);
    nand g1413(n4684 ,n717 ,n4426);
    nor g1414(n1984 ,n862 ,n898);
    nor g1415(n1789 ,n987 ,n1036);
    xnor g1416(n4840 ,n4577 ,n1289);
    nor g1417(n3336 ,n1954 ,n2892);
    nand g1418(n3727 ,n1890 ,n3181);
    nand g1419(n6974 ,n6766 ,n6797);
    xnor g1420(n1914 ,n1[108] ,n2[44]);
    nand g1421(n4577 ,n1068 ,n4216);
    nor g1422(n1021 ,n0[121] ,n0[120]);
    xnor g1423(n1277 ,n6909 ,n6908);
    nand g1424(n9[86] ,n4793 ,n5690);
    xnor g1425(n5056 ,n4595 ,n4447);
    nor g1426(n2345 ,n1[86] ,n1957);
    nor g1427(n5544 ,n4828 ,n5361);
    xnor g1428(n1571 ,n781 ,n1[26]);
    nor g1429(n3106 ,n1488 ,n2568);
    not g1430(n5534 ,n5533);
    nand g1431(n5250 ,n3318 ,n5031);
    nand g1432(n5553 ,n4833 ,n5232);
    or g1433(n4397 ,n3784 ,n4273);
    nand g1434(n1923 ,n0[48] ,n1243);
    nor g1435(n6125 ,n713 ,n6108);
    nand g1436(n1867 ,n0[37] ,n966);
    nand g1437(n3715 ,n3156 ,n2760);
    nand g1438(n570 ,n496 ,n569);
    xnor g1439(n2714 ,n1[118] ,n1506);
    xnor g1440(n85 ,n0[1] ,n7057);
    nand g1441(n6623 ,n1[73] ,n6579);
    xnor g1442(n5015 ,n4[7] ,n4658);
    nor g1443(n2730 ,n724 ,n2042);
    or g1444(n5638 ,n706 ,n5527);
    xnor g1445(n1280 ,n6850 ,n6848);
    or g1446(n170 ,n0[60] ,n1[60]);
    or g1447(n9[37] ,n4485 ,n5898);
    nor g1448(n4884 ,n794 ,n4658);
    xnor g1449(n390 ,n6988 ,n7020);
    nand g1450(n5442 ,n793 ,n5275);
    nor g1451(n3880 ,n2168 ,n3739);
    not g1452(n6189 ,n6190);
    nor g1453(n2488 ,n876 ,n1847);
    nand g1454(n1079 ,n0[127] ,n787);
    nand g1455(n3224 ,n1164 ,n2048);
    nand g1456(n6648 ,n1[81] ,n6579);
    nor g1457(n1007 ,n814 ,n0[64]);
    nor g1458(n5706 ,n5516 ,n5439);
    or g1459(n3029 ,n2162 ,n2297);
    nand g1460(n4502 ,n3938 ,n4155);
    xnor g1461(n2673 ,n1[109] ,n1495);
    or g1462(n2220 ,n1959 ,n1450);
    nor g1463(n3612 ,n834 ,n2971);
    or g1464(n2363 ,n1[56] ,n1958);
    nand g1465(n2461 ,n0[49] ,n718);
    nand g1466(n5434 ,n5243 ,n5247);
    xnor g1467(n1463 ,n1[31] ,n2[31]);
    nand g1468(n2379 ,n707 ,n1512);
    or g1469(n193 ,n0[58] ,n1[58]);
    not g1470(n4900 ,n4899);
    nand g1471(n2459 ,n0[16] ,n1774);
    nand g1472(n115 ,n60 ,n114);
    nor g1473(n3116 ,n1888 ,n2065);
    nor g1474(n2314 ,n721 ,n1538);
    nor g1475(n932 ,n0[94] ,n787);
    nor g1476(n4160 ,n715 ,n4113);
    not g1477(n994 ,n993);
    xnor g1478(n236 ,n0[63] ,n1[63]);
    nand g1479(n2569 ,n0[20] ,n1964);
    nor g1480(n1018 ,n0[91] ,n0[88]);
    nor g1481(n2984 ,n0[65] ,n2483);
    nor g1482(n3388 ,n1954 ,n2917);
    not g1483(n5170 ,n5169);
    nand g1484(n3740 ,n6814 ,n3099);
    nor g1485(n4774 ,n727 ,n687);
    nor g1486(n3979 ,n708 ,n3793);
    xnor g1487(n1266 ,n6933 ,n6932);
    nand g1488(n3982 ,n0[84] ,n3490);
    xnor g1489(n1725 ,n0[29] ,n4[5]);
    not g1490(n6826 ,n6737);
    nor g1491(n5039 ,n727 ,n4927);
    xnor g1492(n1500 ,n0[16] ,n1[16]);
    nand g1493(n302 ,n171 ,n301);
    nor g1494(n3400 ,n1222 ,n2849);
    nor g1495(n4974 ,n4327 ,n4729);
    nand g1496(n1208 ,n1[6] ,n2[6]);
    nor g1497(n5856 ,n713 ,n5771);
    nor g1498(n2292 ,n1961 ,n1941);
    xnor g1499(n6899 ,n101 ,n135);
    nand g1500(n5394 ,n5214 ,n5211);
    xnor g1501(n6901 ,n406 ,n441);
    nand g1502(n4518 ,n2010 ,n4365);
    nand g1503(n3788 ,n6810 ,n3007);
    nand g1504(n5239 ,n5100 ,n5065);
    or g1505(n186 ,n0[42] ,n1[42]);
    nand g1506(n1899 ,n0[63] ,n1221);
    xnor g1507(n229 ,n1[56] ,n0[56]);
    or g1508(n1784 ,n0[65] ,n1004);
    xnor g1509(n2678 ,n1[110] ,n1515);
    not g1510(n785 ,n6869);
    nor g1511(n3398 ,n1954 ,n2921);
    nand g1512(n2579 ,n0[19] ,n1964);
    nand g1513(n4937 ,n4039 ,n4732);
    xnor g1514(n385 ,n7014 ,n7046);
    not g1515(n1011 ,n1010);
    xnor g1516(n1481 ,n1[75] ,n2[11]);
    nand g1517(n5371 ,n4181 ,n5152);
    nand g1518(n2016 ,n714 ,n1021);
    nor g1519(n1763 ,n866 ,n1051);
    nor g1520(n3870 ,n2557 ,n3717);
    nand g1521(n659 ,n1[4] ,n621);
    or g1522(n6484 ,n6434 ,n6341);
    xnor g1523(n1398 ,n1[35] ,n2[35]);
    xnor g1524(n2865 ,n1665 ,n1508);
    not g1525(n5644 ,n5630);
    nand g1526(n3664 ,n0[9] ,n3092);
    xnor g1527(n5568 ,n5377 ,n4811);
    nand g1528(n564 ,n488 ,n563);
    not g1529(n6732 ,n7089);
    xnor g1530(n5198 ,n4991 ,n4841);
    nor g1531(n6573 ,n4851 ,n6565);
    not g1532(n709 ,n715);
    xor g1533(n6346 ,n6246 ,n6143);
    nor g1534(n6406 ,n3447 ,n6332);
    nand g1535(n5899 ,n1953 ,n5768);
    nor g1536(n2976 ,n1046 ,n2176);
    nand g1537(n5133 ,n6827 ,n4894);
    not g1538(n3802 ,n3801);
    xnor g1539(n1282 ,n6945 ,n6944);
    nor g1540(n6709 ,n6826 ,n6584);
    xnor g1541(n2943 ,n1645 ,n1624);
    xnor g1542(n1697 ,n0[77] ,n4[5]);
    xnor g1543(n5455 ,n4430 ,n5157);
    nand g1544(n6661 ,n0[118] ,n0[86]);
    nand g1545(n4273 ,n2142 ,n3973);
    nand g1546(n6683 ,n1[92] ,n6580);
    nand g1547(n5253 ,n791 ,n5082);
    nand g1548(n1949 ,n0[33] ,n1231);
    nor g1549(n912 ,n735 ,n0[1]);
    or g1550(n1239 ,n822 ,n0[50]);
    not g1551(n2565 ,n2564);
    xnor g1552(n6342 ,n5970 ,n6190);
    nand g1553(n130 ,n39 ,n129);
    nand g1554(n7083 ,n665 ,n631);
    not g1555(n825 ,n0[14]);
    nand g1556(n1217 ,n1[65] ,n2[1]);
    nor g1557(n3072 ,n1842 ,n2451);
    nor g1558(n3381 ,n1954 ,n2915);
    or g1559(n31 ,n7065 ,n0[9]);
    nand g1560(n6815 ,n6581 ,n7099);
    nor g1561(n5258 ,n4323 ,n5094);
    nand g1562(n9[5] ,n5404 ,n5906);
    nor g1563(n6297 ,n6236 ,n6202);
    nor g1564(n2030 ,n725 ,n957);
    nor g1565(n1001 ,n738 ,n0[115]);
    nand g1566(n625 ,n0[84] ,n622);
    xnor g1567(n6851 ,n89 ,n111);
    or g1568(n2169 ,n721 ,n1572);
    xnor g1569(n2799 ,n1308 ,n1667);
    nor g1570(n6324 ,n706 ,n6280);
    nor g1571(n896 ,n804 ,n0[2]);
    nand g1572(n6754 ,n0[33] ,n6737);
    nor g1573(n6552 ,n6398 ,n6523);
    nand g1574(n5356 ,n3521 ,n5137);
    nand g1575(n660 ,n1[10] ,n621);
    nor g1576(n3310 ,n2335 ,n3126);
    nand g1577(n4532 ,n2326 ,n4221);
    nor g1578(n4977 ,n3672 ,n4796);
    not g1579(n6205 ,n6204);
    nor g1580(n6595 ,n0[118] ,n0[86]);
    xnor g1581(n1440 ,n1[27] ,n2[27]);
    nor g1582(n2489 ,n993 ,n2008);
    nand g1583(n3742 ,n6812 ,n3053);
    nand g1584(n6064 ,n5789 ,n5995);
    nand g1585(n4819 ,n1966 ,n4442);
    xnor g1586(n1932 ,n0[62] ,n1[62]);
    nor g1587(n3863 ,n2537 ,n3720);
    nor g1588(n3500 ,n6825 ,n2812);
    not g1589(n771 ,n1[46]);
    nand g1590(n222 ,n0[42] ,n1[42]);
    nor g1591(n2204 ,n1958 ,n1617);
    nor g1592(n3427 ,n1222 ,n2837);
    nor g1593(n5180 ,n6824 ,n4905);
    nor g1594(n5416 ,n1954 ,n5245);
    nor g1595(n4401 ,n2544 ,n4355);
    nor g1596(n2477 ,n1956 ,n1610);
    nor g1597(n2994 ,n2615 ,n2354);
    nor g1598(n2407 ,n724 ,n1836);
    not g1599(n5542 ,n5541);
    nand g1600(n220 ,n0[58] ,n1[58]);
    nand g1601(n9[80] ,n5493 ,n6508);
    nand g1602(n3969 ,n3467 ,n3626);
    not g1603(n5472 ,n5471);
    nand g1604(n9[44] ,n5881 ,n5870);
    not g1605(n5068 ,n5067);
    nand g1606(n9[6] ,n5651 ,n5907);
    nor g1607(n2786 ,n721 ,n2429);
    or g1608(n2239 ,n719 ,n1638);
    not g1609(n3251 ,n3250);
    nand g1610(n3157 ,n2599 ,n2471);
    xnor g1611(n5989 ,n5374 ,n5846);
    nand g1612(n6232 ,n3401 ,n6117);
    nor g1613(n3552 ,n1[64] ,n2914);
    xnor g1614(n1286 ,n1[52] ,n4[12]);
    nor g1615(n4603 ,n711 ,n4581);
    xnor g1616(n1404 ,n1[119] ,n2[55]);
    or g1617(n3023 ,n2279 ,n2278);
    nand g1618(n4609 ,n798 ,n4473);
    nand g1619(n9[70] ,n5677 ,n5691);
    nor g1620(n2978 ,n2628 ,n2367);
    nand g1621(n6617 ,n0[103] ,n0[71]);
    nor g1622(n2300 ,n1956 ,n1612);
    nor g1623(n3546 ,n1222 ,n2851);
    xnor g1624(n6204 ,n5770 ,n6110);
    nand g1625(n963 ,n0[84] ,n788);
    nand g1626(n6673 ,n1[90] ,n6580);
    nor g1627(n1803 ,n802 ,n1220);
    nand g1628(n62 ,n7086 ,n0[30]);
    xnor g1629(n5196 ,n4876 ,n1558);
    xnor g1630(n1381 ,n6882 ,n6881);
    nand g1631(n9[33] ,n4599 ,n6391);
    nand g1632(n5720 ,n4822 ,n5492);
    nand g1633(n157 ,n49 ,n156);
    xnor g1634(n1549 ,n0[84] ,n4[28]);
    xnor g1635(n2931 ,n1620 ,n1560);
    nor g1636(n3067 ,n1828 ,n2487);
    nand g1637(n60 ,n7062 ,n0[6]);
    nor g1638(n4624 ,n712 ,n4430);
    xnor g1639(n1371 ,n6905 ,n6904);
    nor g1640(n5173 ,n2991 ,n4963);
    or g1641(n6237 ,n5556 ,n6136);
    xnor g1642(n5465 ,n4663 ,n5154);
    or g1643(n2186 ,n868 ,n2014);
    nor g1644(n2223 ,n1958 ,n1600);
    nor g1645(n5333 ,n3512 ,n5134);
    nor g1646(n2963 ,n1893 ,n2606);
    nand g1647(n5012 ,n4239 ,n4734);
    xnor g1648(n2676 ,n1982 ,n1999);
    nor g1649(n6007 ,n5636 ,n5905);
    nand g1650(n4411 ,n791 ,n4365);
    xnor g1651(n2878 ,n1317 ,n1536);
    xnor g1652(n6871 ,n94 ,n121);
    xnor g1653(n1665 ,n0[9] ,n4[25]);
    xnor g1654(n5570 ,n5276 ,n1637);
    nand g1655(n3791 ,n3190 ,n3189);
    nand g1656(n7000 ,n6684 ,n6808);
    nor g1657(n5448 ,n6 ,n5376);
    nand g1658(n351 ,n7031 ,n6999);
    nand g1659(n223 ,n0[43] ,n1[43]);
    nand g1660(n985 ,n714 ,n766);
    nor g1661(n3737 ,n2558 ,n3263);
    nand g1662(n7040 ,n6662 ,n7133);
    nand g1663(n6487 ,n5997 ,n6438);
    not g1664(n5830 ,n5831);
    xnor g1665(n6198 ,n6106 ,n5838);
    nand g1666(n3470 ,n1953 ,n2942);
    nand g1667(n7073 ,n677 ,n645);
    or g1668(n9[52] ,n4508 ,n5829);
    xnor g1669(n2827 ,n0[103] ,n1251);
    nand g1670(n5510 ,n2326 ,n5379);
    nand g1671(n585 ,n503 ,n584);
    xnor g1672(n6941 ,n385 ,n461);
    nor g1673(n5304 ,n3365 ,n5024);
    or g1674(n2725 ,n725 ,n2643);
    xnor g1675(n1278 ,n0[70] ,n7098);
    xnor g1676(n5018 ,n4594 ,n4104);
    nand g1677(n5007 ,n4803 ,n4748);
    nor g1678(n3911 ,n722 ,n3494);
    nor g1679(n5343 ,n4657 ,n5177);
    xnor g1680(n6947 ,n82 ,n159);
    nand g1681(n6622 ,n0[105] ,n0[73]);
    not g1682(n974 ,n973);
    xnor g1683(n1444 ,n1[120] ,n2[56]);
    nor g1684(n3079 ,n1221 ,n2392);
    nor g1685(n2470 ,n826 ,n1957);
    nand g1686(n4501 ,n3691 ,n4169);
    nand g1687(n6776 ,n1[110] ,n7088);
    nand g1688(n4108 ,n3435 ,n3434);
    nand g1689(n2609 ,n887 ,n1815);
    nor g1690(n4947 ,n2325 ,n4812);
    or g1691(n9[110] ,n5605 ,n5715);
    nor g1692(n1862 ,n759 ,n1220);
    nor g1693(n1808 ,n734 ,n1220);
    nand g1694(n110 ,n14 ,n109);
    nand g1695(n977 ,n0[120] ,n723);
    nor g1696(n5683 ,n5491 ,n5490);
    nand g1697(n4011 ,n0[108] ,n3490);
    nor g1698(n4010 ,n3219 ,n3615);
    nor g1699(n5341 ,n4644 ,n5175);
    xnor g1700(n5977 ,n5843 ,n5461);
    nor g1701(n6608 ,n0[100] ,n0[68]);
    xnor g1702(n4910 ,n2819 ,n4434);
    nor g1703(n2782 ,n2137 ,n2217);
    nand g1704(n363 ,n7036 ,n7004);
    nor g1705(n2746 ,n1[36] ,n2475);
    nand g1706(n6761 ,n0[37] ,n6737);
    or g1707(n486 ,n0[117] ,n6974);
    or g1708(n2464 ,n721 ,n1558);
    nand g1709(n4768 ,n2560 ,n4432);
    nand g1710(n2468 ,n0[67] ,n2028);
    nor g1711(n850 ,n0[19] ,n0[18]);
    xnor g1712(n1451 ,n1[121] ,n2[57]);
    not g1713(n752 ,n0[58]);
    xnor g1714(n1415 ,n1[12] ,n2[12]);
    xor g1715(n7119 ,n0[59] ,n0[27]);
    not g1716(n6425 ,n6402);
    nand g1717(n6636 ,n1[77] ,n6579);
    nand g1718(n4545 ,n1158 ,n4122);
    nand g1719(n4208 ,n791 ,n4117);
    nand g1720(n5004 ,n2516 ,n4674);
    not g1721(n6418 ,n6417);
    nand g1722(n1814 ,n0[48] ,n1225);
    or g1723(n6048 ,n712 ,n5973);
    xor g1724(n696 ,n4664 ,n5458);
    xnor g1725(n2846 ,n1322 ,n1337);
    nand g1726(n669 ,n1[15] ,n621);
    nor g1727(n1744 ,n857 ,n1013);
    or g1728(n189 ,n0[49] ,n1[49]);
    xnor g1729(n1338 ,n6851 ,n6849);
    xnor g1730(n1708 ,n0[71] ,n1[87]);
    nand g1731(n6517 ,n6471 ,n6469);
    nor g1732(n4707 ,n6824 ,n687);
    nand g1733(n4190 ,n792 ,n3953);
    nand g1734(n5122 ,n4043 ,n4946);
    nand g1735(n1831 ,n0[69] ,n964);
    nor g1736(n4340 ,n3607 ,n4093);
    nand g1737(n5386 ,n5037 ,n4795);
    nor g1738(n6507 ,n6456 ,n6404);
    not g1739(n831 ,n0[79]);
    buf g1740(n1954 ,n1642);
    xnor g1741(n1527 ,n0[5] ,n1[5]);
    xnor g1742(n1328 ,n0[45] ,n1[45]);
    or g1743(n2033 ,n719 ,n1486);
    xnor g1744(n6894 ,n252 ,n285);
    nor g1745(n6087 ,n5674 ,n6030);
    xnor g1746(n1947 ,n0[48] ,n1[48]);
    nor g1747(n4982 ,n4185 ,n4784);
    not g1748(n4812 ,n4811);
    nand g1749(n685 ,n1[19] ,n621);
    nand g1750(n930 ,n0[5] ,n709);
    xnor g1751(n5587 ,n5001 ,n5274);
    xnor g1752(n93 ,n0[9] ,n7065);
    nor g1753(n5089 ,n6824 ,n4895);
    nand g1754(n48 ,n7073 ,n0[17]);
    nand g1755(n3599 ,n0[38] ,n2794);
    nand g1756(n4625 ,n3805 ,n4539);
    or g1757(n340 ,n7030 ,n6998);
    nand g1758(n6687 ,n0[126] ,n0[94]);
    xnor g1759(n4880 ,n4428 ,n4585);
    xnor g1760(n1595 ,n0[115] ,n1[115]);
    nor g1761(n5166 ,n6824 ,n4922);
    nor g1762(n2336 ,n1[68] ,n1958);
    nand g1763(n1973 ,n1090 ,n1078);
    nor g1764(n4853 ,n6 ,n4683);
    nand g1765(n4809 ,n3985 ,n4411);
    nor g1766(n4883 ,n792 ,n4671);
    not g1767(n834 ,n1[44]);
    nand g1768(n3999 ,n0[117] ,n3283);
    nor g1769(n1845 ,n813 ,n11);
    xnor g1770(n6852 ,n546 ,n569);
    nand g1771(n637 ,n0[78] ,n622);
    nand g1772(n3269 ,n1952 ,n2857);
    nand g1773(n45 ,n7068 ,n0[12]);
    xnor g1774(n1292 ,n1[43] ,n4[3]);
    nor g1775(n6550 ,n5160 ,n6535);
    nor g1776(n1987 ,n858 ,n955);
    nand g1777(n4779 ,n984 ,n4404);
    nand g1778(n3739 ,n7163 ,n3058);
    nor g1779(n2445 ,n1963 ,n1641);
    xnor g1780(n5449 ,n5018 ,n4221);
    nor g1781(n2484 ,n721 ,n1578);
    xnor g1782(n1344 ,n0[74] ,n4[2]);
    nor g1783(n4635 ,n4058 ,n4383);
    nand g1784(n1202 ,n6947 ,n795);
    nor g1785(n4166 ,n722 ,n4098);
    nand g1786(n150 ,n19 ,n149);
    nor g1787(n6257 ,n711 ,n6249);
    or g1788(n3047 ,n997 ,n2325);
    nor g1789(n5917 ,n711 ,n5830);
    xnor g1790(n1494 ,n0[80] ,n4[24]);
    nor g1791(n2368 ,n0[39] ,n719);
    xnor g1792(n1680 ,n6926 ,n6927);
    nand g1793(n7041 ,n6665 ,n7132);
    or g1794(n2121 ,n1959 ,n1403);
    nand g1795(n9[25] ,n5443 ,n6313);
    nor g1796(n5536 ,n4704 ,n5310);
    nand g1797(n4718 ,n3504 ,n4561);
    or g1798(n13 ,n7075 ,n0[19]);
    nand g1799(n7027 ,n6623 ,n7146);
    nand g1800(n644 ,n0[67] ,n622);
    nor g1801(n5887 ,n792 ,n5731);
    nand g1802(n6774 ,n1[108] ,n7088);
    xnor g1803(n4592 ,n4103 ,n4218);
    nor g1804(n4357 ,n3550 ,n4083);
    xnor g1805(n1368 ,n0[34] ,n0[18]);
    nand g1806(n9[76] ,n5717 ,n6031);
    nand g1807(n4785 ,n2735 ,n4382);
    nand g1808(n287 ,n208 ,n286);
    or g1809(n20 ,n7072 ,n0[16]);
    or g1810(n2442 ,n813 ,n2013);
    not g1811(n6216 ,n6215);
    nand g1812(n3132 ,n1855 ,n2490);
    nand g1813(n507 ,n0[97] ,n6954);
    nor g1814(n2141 ,n1959 ,n1411);
    xor g1815(n7099 ,n0[39] ,n0[7]);
    nand g1816(n140 ,n13 ,n139);
    nor g1817(n3497 ,n6825 ,n2798);
    nor g1818(n6263 ,n1954 ,n6187);
    nand g1819(n5858 ,n1955 ,n5770);
    xor g1820(n2707 ,n1[122] ,n1571);
    nor g1821(n5885 ,n706 ,n696);
    not g1822(n1958 ,n718);
    nand g1823(n517 ,n0[103] ,n6960);
    not g1824(n1965 ,n1966);
    nand g1825(n618 ,n481 ,n617);
    nor g1826(n2267 ,n6 ,n2026);
    nand g1827(n10[2] ,n4502 ,n4982);
    nor g1828(n3266 ,n1222 ,n2839);
    xnor g1829(n5200 ,n4[13] ,n4992);
    or g1830(n4134 ,n1962 ,n3828);
    nand g1831(n3240 ,n1216 ,n2166);
    xnor g1832(n2698 ,n1651 ,n1600);
    xnor g1833(n1324 ,n0[44] ,n1[60]);
    nand g1834(n414 ,n318 ,n413);
    nor g1835(n2327 ,n1997 ,n2030);
    xnor g1836(n5591 ,n5207 ,n1625);
    xnor g1837(n402 ,n7000 ,n7032);
    nand g1838(n416 ,n331 ,n415);
    nor g1839(n4452 ,n4164 ,n4130);
    nor g1840(n1892 ,n821 ,n1226);
    nor g1841(n4039 ,n3748 ,n3011);
    nor g1842(n2761 ,n2083 ,n2089);
    xnor g1843(n1314 ,n0[122] ,n4[10]);
    xnor g1844(n6513 ,n6170 ,n6414);
    nand g1845(n503 ,n0[109] ,n6966);
    nor g1846(n5906 ,n5745 ,n5820);
    nor g1847(n1723 ,n1052 ,n1022);
    nor g1848(n5418 ,n5095 ,n5295);
    xnor g1849(n550 ,n6963 ,n0[106]);
    nand g1850(n3077 ,n1220 ,n2353);
    nand g1851(n6814 ,n6581 ,n7100);
    nor g1852(n4471 ,n792 ,n4209);
    xnor g1853(n6463 ,n6312 ,n1716);
    nor g1854(n5492 ,n3466 ,n5389);
    or g1855(n979 ,n725 ,n0[51]);
    or g1856(n4792 ,n3697 ,n4512);
    nand g1857(n286 ,n172 ,n285);
    nand g1858(n6505 ,n5660 ,n6405);
    nor g1859(n4353 ,n3174 ,n4096);
    not g1860(n1534 ,n1533);
    xnor g1861(n1694 ,n0[65] ,n1[81]);
    nor g1862(n6722 ,n6826 ,n6598);
    nand g1863(n3123 ,n972 ,n2111);
    nand g1864(n3790 ,n3154 ,n3175);
    nand g1865(n6652 ,n0[115] ,n0[83]);
    nor g1866(n6404 ,n3286 ,n6352);
    nor g1867(n2638 ,n0[7] ,n721);
    nor g1868(n4070 ,n708 ,n3792);
    or g1869(n6081 ,n6025 ,n5781);
    nand g1870(n3339 ,n1953 ,n2917);
    nand g1871(n3207 ,n1108 ,n2077);
    nor g1872(n6124 ,n706 ,n6110);
    not g1873(n1056 ,n1055);
    or g1874(n9[49] ,n4801 ,n6394);
    nor g1875(n4960 ,n3535 ,n4776);
    or g1876(n3391 ,n3004 ,n2135);
    nand g1877(n6177 ,n1955 ,n6141);
    or g1878(n4062 ,n3659 ,n3507);
    xnor g1879(n238 ,n1[34] ,n0[34]);
    xnor g1880(n1460 ,n0[83] ,n1[83]);
    nor g1881(n2372 ,n0[44] ,n719);
    nand g1882(n883 ,n0[15] ,n710);
    nand g1883(n3151 ,n1[68] ,n2337);
    nand g1884(n2559 ,n1195 ,n1863);
    nor g1885(n902 ,n0[103] ,n790);
    nor g1886(n2202 ,n715 ,n1445);
    nand g1887(n961 ,n0[85] ,n790);
    nand g1888(n3395 ,n2316 ,n2755);
    or g1889(n9[17] ,n6537 ,n6388);
    nand g1890(n2563 ,n0[21] ,n707);
    xnor g1891(n1626 ,n0[88] ,n1[88]);
    nor g1892(n877 ,n0[24] ,n723);
    not g1893(n4676 ,n4675);
    nor g1894(n5754 ,n5646 ,n5645);
    nor g1895(n5882 ,n5766 ,n5758);
    nand g1896(n3229 ,n1204 ,n2109);
    nand g1897(n6460 ,n6374 ,n6283);
    nand g1898(n299 ,n198 ,n298);
    nand g1899(n1042 ,n723 ,n754);
    nand g1900(n50 ,n7070 ,n0[14]);
    nor g1901(n6128 ,n713 ,n6111);
    xnor g1902(n5595 ,n5197 ,n5210);
    nand g1903(n1175 ,n6891 ,n795);
    nand g1904(n3793 ,n3201 ,n3200);
    nand g1905(n3281 ,n1952 ,n2861);
    nor g1906(n5736 ,n712 ,n5582);
    nand g1907(n1055 ,n0[122] ,n740);
    nand g1908(n5625 ,n4957 ,n5471);
    xnor g1909(n3825 ,n1[74] ,n2663);
    nor g1910(n2320 ,n1958 ,n1640);
    xnor g1911(n1719 ,n7093 ,n7051);
    not g1912(n817 ,n0[13]);
    xnor g1913(n246 ,n1[42] ,n0[42]);
    nand g1914(n1188 ,n6901 ,n797);
    nor g1915(n2047 ,n1963 ,n1548);
    nor g1916(n5296 ,n794 ,n5057);
    nand g1917(n1028 ,n0[1] ,n811);
    xnor g1918(n1505 ,n0[63] ,n4[23]);
    xnor g1919(n2910 ,n1[99] ,n1557);
    nor g1920(n6333 ,n711 ,n6305);
    nand g1921(n113 ,n55 ,n112);
    nand g1922(n3479 ,n714 ,n2726);
    nand g1923(n4289 ,n0[36] ,n3873);
    nor g1924(n5631 ,n3288 ,n5405);
    xnor g1925(n4211 ,n3538 ,n1996);
    or g1926(n5103 ,n706 ,n4994);
    xnor g1927(n6900 ,n558 ,n593);
    or g1928(n5446 ,n5300 ,n5281);
    xnor g1929(n1565 ,n1[16] ,n763);
    nand g1930(n5757 ,n1955 ,n5585);
    nand g1931(n4115 ,n3000 ,n3609);
    nand g1932(n4755 ,n717 ,n4583);
    nand g1933(n6982 ,n6744 ,n6771);
    nand g1934(n3846 ,n2033 ,n3477);
    nor g1935(n1951 ,n0[0] ,n1029);
    nand g1936(n3217 ,n1150 ,n2086);
    nor g1937(n5487 ,n3413 ,n5285);
    nor g1938(n4850 ,n6 ,n4809);
    nand g1939(n3450 ,n709 ,n3257);
    nand g1940(n6495 ,n6450 ,n6345);
    nand g1941(n1143 ,n6917 ,n795);
    nand g1942(n1163 ,n6905 ,n796);
    nand g1943(n5865 ,n1953 ,n5728);
    xnor g1944(n5975 ,n5839 ,n5462);
    or g1945(n2980 ,n2023 ,n2329);
    nand g1946(n6050 ,n717 ,n5973);
    or g1947(n6427 ,n6083 ,n6336);
    nor g1948(n1880 ,n829 ,n11);
    xnor g1949(n2936 ,n1683 ,n1623);
    nand g1950(n308 ,n169 ,n307);
    nor g1951(n3009 ,n1872 ,n2235);
    or g1952(n2075 ,n719 ,n1625);
    nand g1953(n2518 ,n793 ,n1982);
    nand g1954(n421 ,n365 ,n420);
    or g1955(n5664 ,n4395 ,n5470);
    nor g1956(n3484 ,n1954 ,n2950);
    or g1957(n4395 ,n3783 ,n4282);
    nor g1958(n6726 ,n6826 ,n6602);
    nand g1959(n5399 ,n5222 ,n5220);
    xnor g1960(n1939 ,n1[84] ,n2[20]);
    xnor g1961(n5476 ,n4662 ,n5155);
    nand g1962(n2024 ,n723 ,n1024);
    xnor g1963(n4445 ,n2800 ,n3951);
    not g1964(n798 ,n6824);
    nor g1965(n1013 ,n0[109] ,n787);
    nand g1966(n630 ,n0[75] ,n622);
    or g1967(n4787 ,n6823 ,n4438);
    nand g1968(n2548 ,n1165 ,n1876);
    nand g1969(n4128 ,n2560 ,n3940);
    nand g1970(n2365 ,n1964 ,n1515);
    nand g1971(n9[0] ,n5329 ,n6377);
    nand g1972(n6179 ,n1952 ,n6120);
    nor g1973(n2034 ,n1963 ,n1486);
    xnor g1974(n1579 ,n1[55] ,n1[23]);
    xor g1975(n7094 ,n0[34] ,n0[2]);
    nand g1976(n72 ,n7056 ,n0[0]);
    xnor g1977(n6514 ,n6386 ,n6387);
    nand g1978(n3724 ,n1144 ,n3049);
    nor g1979(n5306 ,n4311 ,n5171);
    nand g1980(n6268 ,n1955 ,n6246);
    nand g1981(n2467 ,n0[3] ,n2029);
    nand g1982(n3957 ,n3451 ,n3450);
    xnor g1983(n1660 ,n1[126] ,n4[6]);
    xnor g1984(n1635 ,n0[73] ,n1[73]);
    nor g1985(n6256 ,n6012 ,n6215);
    nand g1986(n281 ,n199 ,n280);
    nand g1987(n3929 ,n2990 ,n3594);
    nand g1988(n4406 ,n793 ,n4218);
    nor g1989(n4876 ,n953 ,n4672);
    not g1990(n3804 ,n3803);
    or g1991(n2145 ,n721 ,n1453);
    nand g1992(n1173 ,n6841 ,n796);
    nand g1993(n1073 ,n0[31] ,n787);
    nand g1994(n969 ,n723 ,n822);
    xnor g1995(n1554 ,n1[56] ,n1[24]);
    xnor g1996(n2875 ,n1295 ,n1368);
    nor g1997(n4026 ,n3229 ,n3384);
    or g1998(n3301 ,n1954 ,n2874);
    nor g1999(n6184 ,n5551 ,n6159);
    nand g2000(n5875 ,n1952 ,n5734);
    xnor g2001(n4885 ,n4213 ,n4568);
    nor g2002(n2405 ,n724 ,n1791);
    nor g2003(n4008 ,n3220 ,n3612);
    or g2004(n6303 ,n6162 ,n6191);
    nand g2005(n5388 ,n4818 ,n5164);
    xnor g2006(n1693 ,n1[117] ,n4[13]);
    xnor g2007(n1496 ,n1[51] ,n1[19]);
    nor g2008(n1728 ,n0[48] ,n1243);
    xor g2009(n7100 ,n0[40] ,n0[8]);
    xnor g2010(n1255 ,n1[44] ,n4[4]);
    xnor g2011(n5579 ,n1354 ,n5205);
    nor g2012(n2263 ,n6 ,n1995);
    nand g2013(n4329 ,n2589 ,n3901);
    nand g2014(n3744 ,n6811 ,n3141);
    nand g2015(n3228 ,n1192 ,n2035);
    xnor g2016(n1339 ,n0[85] ,n7113);
    nand g2017(n4332 ,n2580 ,n3891);
    nor g2018(n1966 ,n7089 ,n1240);
    nand g2019(n4859 ,n3371 ,n4604);
    nor g2020(n3001 ,n2207 ,n2435);
    nand g2021(n619 ,n518 ,n618);
    or g2022(n3285 ,n1954 ,n2871);
    nand g2023(n7130 ,n6669 ,n6722);
    xnor g2024(n1556 ,n0[11] ,n1[11]);
    nand g2025(n6788 ,n1[127] ,n7088);
    nand g2026(n6778 ,n1[121] ,n7088);
    xnor g2027(n1598 ,n0[98] ,n1[98]);
    nor g2028(n2737 ,n1767 ,n2508);
    nor g2029(n4135 ,n1962 ,n3917);
    nand g2030(n1851 ,n0[22] ,n1221);
    nand g2031(n4109 ,n3040 ,n3573);
    nand g2032(n6057 ,n6016 ,n5778);
    nor g2033(n2639 ,n0[0] ,n1963);
    nor g2034(n2332 ,n1[61] ,n1956);
    nand g2035(n10[30] ,n4633 ,n4866);
    or g2036(n104 ,n72 ,n21);
    nand g2037(n2010 ,n0[120] ,n1009);
    nor g2038(n1842 ,n814 ,n11);
    nor g2039(n1946 ,n803 ,n1097);
    nand g2040(n3082 ,n11 ,n2396);
    nand g2041(n2432 ,n0[42] ,n718);
    xnor g2042(n1699 ,n1[119] ,n4[15]);
    nand g2043(n358 ,n7042 ,n7010);
    nor g2044(n2111 ,n1033 ,n1951);
    xnor g2045(n5075 ,n4806 ,n4426);
    or g2046(n3393 ,n1954 ,n2920);
    nand g2047(n1169 ,n6933 ,n797);
    xnor g2048(n2693 ,n0[55] ,n1970);
    nor g2049(n1734 ,n1032 ,n849);
    nor g2050(n2420 ,n1957 ,n1586);
    nand g2051(n10[5] ,n4617 ,n5317);
    nand g2052(n4822 ,n1966 ,n4439);
    nor g2053(n4852 ,n2325 ,n4683);
    nand g2054(n1224 ,n0[50] ,n822);
    nand g2055(n6821 ,n6581 ,n7093);
    nand g2056(n2778 ,n1555 ,n2623);
    nor g2057(n2364 ,n0[55] ,n719);
    or g2058(n329 ,n7048 ,n7016);
    nand g2059(n3542 ,n1953 ,n2960);
    nor g2060(n4191 ,n3980 ,n3789);
    or g2061(n1790 ,n725 ,n1231);
    nand g2062(n565 ,n525 ,n564);
    nor g2063(n3290 ,n1954 ,n2866);
    nand g2064(n1983 ,n1077 ,n1064);
    nor g2065(n2435 ,n1962 ,n1405);
    nand g2066(n624 ,n0[90] ,n622);
    nor g2067(n2191 ,n1963 ,n1520);
    nor g2068(n3798 ,n6825 ,n2804);
    nand g2069(n4677 ,n3888 ,n4528);
    nand g2070(n7084 ,n675 ,n640);
    not g2071(n6073 ,n6072);
    nand g2072(n6991 ,n6620 ,n6817);
    nor g2073(n4589 ,n2732 ,n4348);
    xnor g2074(n6857 ,n395 ,n419);
    nor g2075(n1838 ,n0[27] ,n1012);
    nor g2076(n3323 ,n1954 ,n2887);
    xnor g2077(n4479 ,n3944 ,n2839);
    nor g2078(n6716 ,n6826 ,n6583);
    nand g2079(n196 ,n0[60] ,n1[60]);
    xnor g2080(n1658 ,n6902 ,n6903);
    nand g2081(n7134 ,n6658 ,n6718);
    or g2082(n191 ,n0[46] ,n1[46]);
    or g2083(n6411 ,n6082 ,n6349);
    nand g2084(n4964 ,n3372 ,n4607);
    nor g2085(n2729 ,n724 ,n2041);
    nand g2086(n221 ,n0[35] ,n1[35]);
    not g2087(n5990 ,n5989);
    or g2088(n4719 ,n3500 ,n4562);
    nor g2089(n6252 ,n712 ,n6189);
    nor g2090(n2334 ,n0[43] ,n1957);
    nor g2091(n5405 ,n706 ,n5268);
    nand g2092(n4391 ,n787 ,n4234);
    nor g2093(n5745 ,n1954 ,n5588);
    nor g2094(n3462 ,n6823 ,n2822);
    not g2095(n6580 ,n6578);
    or g2096(n2040 ,n952 ,n2021);
    nand g2097(n6628 ,n0[106] ,n0[74]);
    nand g2098(n640 ,n0[92] ,n622);
    nand g2099(n3646 ,n2469 ,n2789);
    nand g2100(n3610 ,n1[36] ,n3095);
    not g2101(n6220 ,n6219);
    or g2102(n4066 ,n3667 ,n3796);
    nor g2103(n5658 ,n6 ,n5531);
    xnor g2104(n1646 ,n0[43] ,n1[59]);
    nor g2105(n3425 ,n710 ,n3250);
    nor g2106(n5011 ,n2719 ,n4778);
    nand g2107(n5558 ,n4823 ,n5236);
    xnor g2108(n5206 ,n4682 ,n5006);
    nand g2109(n6276 ,n6223 ,n6205);
    not g2110(n795 ,n6826);
    nand g2111(n7002 ,n6694 ,n6806);
    nand g2112(n1088 ,n0[87] ,n791);
    or g2113(n10[28] ,n4864 ,n4696);
    nand g2114(n1071 ,n0[95] ,n787);
    nand g2115(n4829 ,n1966 ,n4433);
    nor g2116(n5655 ,n4489 ,n5532);
    or g2117(n2331 ,n0[59] ,n1958);
    xnor g2118(n1532 ,n0[54] ,n4[14]);
    nand g2119(n5379 ,n3886 ,n5022);
    xnor g2120(n2920 ,n1669 ,n1505);
    not g2121(n5970 ,n5969);
    nor g2122(n2094 ,n1962 ,n1388);
    nand g2123(n5518 ,n3654 ,n5259);
    nand g2124(n9[121] ,n5118 ,n6396);
    not g2125(n4658 ,n4659);
    nor g2126(n4248 ,n1960 ,n3815);
    nand g2127(n5711 ,n4007 ,n5482);
    nand g2128(n3318 ,n1952 ,n2882);
    nor g2129(n2289 ,n1958 ,n1592);
    nand g2130(n4546 ,n1128 ,n4121);
    xnor g2131(n2922 ,n1611 ,n1543);
    nor g2132(n5231 ,n3445 ,n5186);
    nor g2133(n1022 ,n0[110] ,n715);
    nor g2134(n1731 ,n1050 ,n855);
    xnor g2135(n1296 ,n1[15] ,n4[15]);
    nand g2136(n3623 ,n1[47] ,n2795);
    nor g2137(n4946 ,n3510 ,n4733);
    xnor g2138(n2800 ,n0[111] ,n1302);
    nand g2139(n5826 ,n4184 ,n5714);
    nand g2140(n1836 ,n0[40] ,n916);
    xnor g2141(n6866 ,n245 ,n271);
    nand g2142(n4348 ,n2439 ,n4028);
    or g2143(n5083 ,n712 ,n4988);
    nand g2144(n3127 ,n1[41] ,n2612);
    nand g2145(n5142 ,n6827 ,n4910);
    xnor g2146(n1391 ,n1[53] ,n2[53]);
    nor g2147(n5872 ,n706 ,n5839);
    nand g2148(n2593 ,n0[1] ,n707);
    nand g2149(n663 ,n1[12] ,n621);
    nor g2150(n3518 ,n6825 ,n2828);
    nand g2151(n5860 ,n717 ,n5726);
    nor g2152(n5701 ,n5507 ,n5522);
    not g2153(n6068 ,n6067);
    nor g2154(n5648 ,n4785 ,n5562);
    not g2155(n820 ,n0[64]);
    nor g2156(n6319 ,n6254 ,n6253);
    nand g2157(n5095 ,n4240 ,n4869);
    nand g2158(n3650 ,n0[0] ,n3075);
    not g2159(n739 ,n0[74]);
    nor g2160(n2261 ,n1961 ,n1397);
    xor g2161(n7097 ,n0[37] ,n0[5]);
    or g2162(n9[58] ,n4503 ,n6296);
    nor g2163(n5104 ,n712 ,n4995);
    nand g2164(n668 ,n1[23] ,n621);
    nand g2165(n1213 ,n0[12] ,n791);
    nand g2166(n4351 ,n3600 ,n4014);
    nand g2167(n518 ,n0[126] ,n6983);
    nand g2168(n7034 ,n6645 ,n7139);
    nand g2169(n3760 ,n6805 ,n3065);
    nand g2170(n3196 ,n0[66] ,n2506);
    nand g2171(n1642 ,n1211 ,n973);
    nor g2172(n4751 ,n6 ,n4587);
    nor g2173(n3859 ,n2045 ,n3729);
    nand g2174(n6625 ,n0[83] ,n6580);
    or g2175(n6482 ,n6432 ,n6348);
    nand g2176(n1167 ,n6925 ,n795);
    nand g2177(n4764 ,n2560 ,n4457);
    nor g2178(n3344 ,n1954 ,n2897);
    nand g2179(n5520 ,n4178 ,n5370);
    nor g2180(n4680 ,n4527 ,n4376);
    or g2181(n3057 ,n0[32] ,n2205);
    nor g2182(n3712 ,n2219 ,n3193);
    nor g2183(n325 ,n7019 ,n6987);
    nand g2184(n1024 ,n0[25] ,n737);
    xnor g2185(n4466 ,n3947 ,n2814);
    nor g2186(n5237 ,n3544 ,n5176);
    nand g2187(n4713 ,n717 ,n4425);
    or g2188(n2066 ,n719 ,n1526);
    nand g2189(n1832 ,n0[58] ,n1221);
    nor g2190(n6259 ,n712 ,n6246);
    nand g2191(n654 ,n0[95] ,n622);
    xnor g2192(n6315 ,n6176 ,n5946);
    nand g2193(n5124 ,n4046 ,n4951);
    nand g2194(n2482 ,n0[115] ,n2021);
    nand g2195(n2431 ,n0[43] ,n718);
    nor g2196(n927 ,n0[47] ,n790);
    xnor g2197(n4403 ,n3811 ,n1974);
    nand g2198(n593 ,n504 ,n592);
    nand g2199(n6172 ,n5442 ,n6071);
    nand g2200(n4290 ,n3618 ,n4036);
    nor g2201(n3056 ,n1802 ,n2311);
    nand g2202(n699 ,n5893 ,n5975);
    nand g2203(n357 ,n7033 ,n7001);
    nand g2204(n119 ,n63 ,n118);
    nand g2205(n5779 ,n717 ,n5640);
    not g2206(n5485 ,n5433);
    nand g2207(n623 ,n0[71] ,n622);
    xnor g2208(n1639 ,n0[15] ,n1[15]);
    nor g2209(n3448 ,n1954 ,n2933);
    nor g2210(n5890 ,n712 ,n5834);
    nor g2211(n2241 ,n1959 ,n1399);
    or g2212(n4243 ,n1965 ,n3943);
    nand g2213(n590 ,n476 ,n589);
    nor g2214(n2153 ,n913 ,n1962);
    nand g2215(n2035 ,n718 ,n1483);
    nand g2216(n4006 ,n0[29] ,n3490);
    nand g2217(n1192 ,n6948 ,n796);
    or g2218(n2380 ,n1[40] ,n1958);
    nor g2219(n3534 ,n6825 ,n2846);
    or g2220(n184 ,n0[35] ,n1[35]);
    or g2221(n185 ,n0[40] ,n1[40]);
    nand g2222(n224 ,n0[32] ,n1[32]);
    nand g2223(n5647 ,n717 ,n5527);
    xnor g2224(n5573 ,n5209 ,n1537);
    xnor g2225(n2880 ,n1681 ,n1509);
    xnor g2226(n1706 ,n0[70] ,n1[86]);
    nand g2227(n7059 ,n678 ,n644);
    nand g2228(n6109 ,n4642 ,n5978);
    not g2229(n4891 ,n4890);
    nor g2230(n1735 ,n1226 ,n1003);
    xnor g2231(n2961 ,n1[124] ,n1553);
    nor g2232(n3853 ,n3242 ,n3679);
    or g2233(n2109 ,n719 ,n1508);
    nand g2234(n6274 ,n6181 ,n6197);
    nand g2235(n411 ,n361 ,n410);
    nand g2236(n4727 ,n2326 ,n4453);
    nand g2237(n4583 ,n2517 ,n4224);
    nand g2238(n3334 ,n1953 ,n2892);
    xnor g2239(n2653 ,n1693 ,n1564);
    nand g2240(n6699 ,n1[66] ,n6580);
    nand g2241(n7087 ,n686 ,n654);
    xnor g2242(n2896 ,n1258 ,n1359);
    or g2243(n480 ,n0[121] ,n6978);
    xnor g2244(n5985 ,n5270 ,n5841);
    xnor g2245(n1624 ,n0[113] ,n1[113]);
    nand g2246(n614 ,n474 ,n613);
    nor g2247(n2770 ,n1531 ,n2625);
    nor g2248(n2149 ,n6 ,n1738);
    xnor g2249(n4835 ,n4579 ,n2660);
    nand g2250(n4656 ,n792 ,n4459);
    nor g2251(n6306 ,n5649 ,n6192);
    or g2252(n2201 ,n1960 ,n1435);
    nor g2253(n4454 ,n2505 ,n4231);
    nand g2254(n935 ,n0[7] ,n709);
    nand g2255(n1199 ,n6839 ,n795);
    nand g2256(n6763 ,n0[38] ,n6737);
    xnor g2257(n5459 ,n4577 ,n5156);
    xnor g2258(n1458 ,n1[95] ,n2[31]);
    xnor g2259(n6846 ,n240 ,n261);
    nand g2260(n6452 ,n3343 ,n6334);
    nor g2261(n4151 ,n4047 ,n3770);
    nor g2262(n5053 ,n4889 ,n4885);
    nor g2263(n5837 ,n4199 ,n5718);
    nor g2264(n5966 ,n5930 ,n5885);
    xnor g2265(n1676 ,n0[106] ,n4[2]);
    or g2266(n1998 ,n0[9] ,n1246);
    nand g2267(n3934 ,n2151 ,n3633);
    nand g2268(n6780 ,n1[126] ,n7088);
    nand g2269(n508 ,n0[119] ,n6976);
    nor g2270(n4703 ,n6824 ,n4477);
    nor g2271(n2369 ,n0[49] ,n1956);
    xnor g2272(n2711 ,n1980 ,n1973);
    xnor g2273(n6878 ,n248 ,n277);
    nand g2274(n1238 ,n0[93] ,n715);
    nand g2275(n4307 ,n720 ,n3831);
    nor g2276(n5794 ,n5533 ,n5693);
    nand g2277(n3685 ,n1[50] ,n2978);
    nand g2278(n3307 ,n1952 ,n2879);
    xnor g2279(n4432 ,n2834 ,n3952);
    xnor g2280(n4927 ,n2846 ,n4463);
    nor g2281(n3143 ,n1568 ,n2565);
    xnor g2282(n1468 ,n1[66] ,n2[2]);
    nor g2283(n2026 ,n865 ,n1022);
    nor g2284(n973 ,n3[2] ,n3[1]);
    xnor g2285(n3835 ,n1[89] ,n2713);
    nand g2286(n3380 ,n2167 ,n3070);
    nand g2287(n6740 ,n0[42] ,n6737);
    nand g2288(n3711 ,n2213 ,n3192);
    xnor g2289(n4846 ,n4371 ,n4369);
    nor g2290(n4675 ,n793 ,n4410);
    nor g2291(n2265 ,n940 ,n1759);
    nor g2292(n3426 ,n1954 ,n2928);
    or g2293(n10[13] ,n4986 ,n5498);
    nor g2294(n3099 ,n1854 ,n2194);
    xnor g2295(n1295 ,n1[34] ,n4[26]);
    nor g2296(n2382 ,n0[63] ,n1956);
    nor g2297(n4664 ,n2260 ,n4471);
    or g2298(n2440 ,n816 ,n1544);
    or g2299(n10[14] ,n4985 ,n5436);
    or g2300(n6085 ,n3374 ,n5951);
    nor g2301(n5041 ,n727 ,n4905);
    or g2302(n3504 ,n6825 ,n2815);
    nor g2303(n5893 ,n711 ,n5846);
    nand g2304(n4390 ,n794 ,n4222);
    not g2305(n6107 ,n6108);
    nand g2306(n521 ,n0[116] ,n6973);
    nor g2307(n2659 ,n2422 ,n2202);
    nor g2308(n6589 ,n0[112] ,n0[80]);
    not g2309(n1045 ,n1044);
    nand g2310(n6634 ,n1[76] ,n6579);
    xnor g2311(n1345 ,n0[0] ,n4[16]);
    nor g2312(n3308 ,n1954 ,n2879);
    nand g2313(n6679 ,n0[112] ,n0[80]);
    nand g2314(n4075 ,n3643 ,n3637);
    nor g2315(n4015 ,n791 ,n3519);
    not g2316(n1540 ,n1539);
    nand g2317(n5213 ,n4952 ,n5078);
    xnor g2318(n1418 ,n1[0] ,n2[0]);
    or g2319(n4674 ,n794 ,n4403);
    not g2320(n2904 ,n2903);
    xnor g2321(n5732 ,n5460 ,n2709);
    nor g2322(n6390 ,n5093 ,n6358);
    xnor g2323(n1650 ,n0[105] ,n4[1]);
    or g2324(n5776 ,n713 ,n5640);
    xor g2325(n702 ,n6249 ,n6172);
    nand g2326(n7142 ,n6635 ,n6710);
    nor g2327(n2288 ,n1963 ,n1556);
    nand g2328(n936 ,n0[27] ,n805);
    nand g2329(n2031 ,n936 ,n2025);
    nor g2330(n2117 ,n1960 ,n1466);
    nor g2331(n6157 ,n4928 ,n6055);
    nand g2332(n1147 ,n6867 ,n797);
    nor g2333(n3044 ,n725 ,n2093);
    nand g2334(n6793 ,n1[123] ,n7088);
    not g2335(n1221 ,n11);
    nand g2336(n7129 ,n6680 ,n6723);
    nand g2337(n645 ,n0[81] ,n622);
    xnor g2338(n1349 ,n0[2] ,n4[18]);
    nor g2339(n1747 ,n0[122] ,n999);
    nor g2340(n3422 ,n2158 ,n3017);
    nor g2341(n3406 ,n1954 ,n2941);
    not g2342(n4814 ,n4813);
    xnor g2343(n1590 ,n0[79] ,n1[79]);
    nand g2344(n6777 ,n1[120] ,n7088);
    nand g2345(n3168 ,n2579 ,n2492);
    nor g2346(n6593 ,n0[114] ,n0[82]);
    nand g2347(n4148 ,n3469 ,n4045);
    nor g2348(n4855 ,n3400 ,n4707);
    nor g2349(n3523 ,n2138 ,n3124);
    nor g2350(n4991 ,n2513 ,n4678);
    or g2351(n4202 ,n2325 ,n3950);
    nor g2352(n2499 ,n1958 ,n1457);
    nand g2353(n2744 ,n1551 ,n2619);
    or g2354(n6486 ,n6375 ,n6415);
    not g2355(n1953 ,n1954);
    nor g2356(n5087 ,n6824 ,n4893);
    nor g2357(n910 ,n0[69] ,n0[13]);
    nor g2358(n5174 ,n6824 ,n4925);
    nor g2359(n2413 ,n0[53] ,n719);
    xnor g2360(n1720 ,n0[46] ,n0[30]);
    nand g2361(n7014 ,n6614 ,n7159);
    xnor g2362(n6868 ,n550 ,n577);
    nand g2363(n4820 ,n1966 ,n4440);
    xnor g2364(n3840 ,n1[95] ,n2657);
    not g2365(n734 ,n0[75]);
    xnor g2366(n1383 ,n6941 ,n6940);
    nor g2367(n2743 ,n718 ,n2350);
    nand g2368(n354 ,n7032 ,n7000);
    nand g2369(n6678 ,n0[104] ,n0[72]);
    nand g2370(n1210 ,n0[4] ,n709);
    nand g2371(n4757 ,n717 ,n4574);
    nand g2372(n7028 ,n6626 ,n7145);
    nand g2373(n2514 ,n1883 ,n1870);
    nor g2374(n3915 ,n2315 ,n3760);
    nor g2375(n4953 ,n4198 ,n4598);
    xnor g2376(n1469 ,n1[114] ,n2[50]);
    not g2377(n6344 ,n6343);
    nor g2378(n6521 ,n5548 ,n6476);
    nand g2379(n3243 ,n0[98] ,n2555);
    or g2380(n5426 ,n5105 ,n5276);
    or g2381(n4491 ,n2542 ,n4168);
    not g2382(n3942 ,n3941);
    nand g2383(n4753 ,n715 ,n4474);
    nor g2384(n1852 ,n821 ,n1220);
    nor g2385(n6515 ,n5094 ,n6470);
    nand g2386(n6239 ,n3995 ,n6134);
    nand g2387(n3662 ,n0[50] ,n2986);
    or g2388(n1766 ,n0[104] ,n885);
    nand g2389(n3022 ,n1220 ,n2349);
    xnor g2390(n538 ,n6982 ,n0[125]);
    nor g2391(n3904 ,n2252 ,n3686);
    xor g2392(n6828 ,n6953 ,n0[96]);
    nor g2393(n3366 ,n1954 ,n2913);
    nand g2394(n2549 ,n1127 ,n1896);
    nand g2395(n2475 ,n0[4] ,n1964);
    xnor g2396(n6842 ,n239 ,n259);
    nand g2397(n7013 ,n6677 ,n7160);
    nand g2398(n6958 ,n6761 ,n6794);
    nand g2399(n4772 ,n2560 ,n4440);
    nor g2400(n6027 ,n3356 ,n5876);
    nand g2401(n6287 ,n6010 ,n6209);
    nand g2402(n4001 ,n0[92] ,n3490);
    nand g2403(n9[30] ,n5045 ,n5663);
    xnor g2404(n1423 ,n1[16] ,n2[16]);
    nand g2405(n3702 ,n782 ,n3167);
    nand g2406(n6265 ,n717 ,n6245);
    nand g2407(n1879 ,n765 ,n980);
    nor g2408(n6150 ,n5562 ,n698);
    or g2409(n336 ,n7021 ,n6989);
    nor g2410(n6183 ,n5468 ,n6138);
    nor g2411(n5301 ,n3527 ,n5042);
    or g2412(n16 ,n7076 ,n0[20]);
    nor g2413(n6528 ,n4728 ,n6490);
    or g2414(n4057 ,n2572 ,n3764);
    nand g2415(n4524 ,n4319 ,n4158);
    nor g2416(n4177 ,n3222 ,n4075);
    or g2417(n9[18] ,n4524 ,n6237);
    xnor g2418(n1634 ,n0[106] ,n1[106]);
    nor g2419(n1816 ,n0[48] ,n969);
    nand g2420(n5130 ,n4026 ,n4849);
    nor g2421(n5714 ,n2551 ,n5505);
    or g2422(n4686 ,n711 ,n4429);
    nand g2423(n1068 ,n0[52] ,n792);
    xnor g2424(n5575 ,n5005 ,n5376);
    nor g2425(n5507 ,n4871 ,n5291);
    nand g2426(n4549 ,n1169 ,n4140);
    nand g2427(n3681 ,n3149 ,n2084);
    nor g2428(n3403 ,n1222 ,n2799);
    nor g2429(n6012 ,n3328 ,n5902);
    nor g2430(n2051 ,n1960 ,n1948);
    nor g2431(n4267 ,n3216 ,n3875);
    nor g2432(n4193 ,n6 ,n4104);
    xnor g2433(n2668 ,n1690 ,n1502);
    xnor g2434(n2836 ,n0[121] ,n1377);
    nor g2435(n2433 ,n989 ,n1775);
    nor g2436(n4863 ,n4150 ,n4709);
    nand g2437(n627 ,n0[73] ,n622);
    or g2438(n6557 ,n5383 ,n6527);
    nand g2439(n2603 ,n0[8] ,n707);
    xnor g2440(n1351 ,n0[44] ,n0[28]);
    nand g2441(n506 ,n0[110] ,n6967);
    nor g2442(n6548 ,n5561 ,n6516);
    nand g2443(n3407 ,n1953 ,n2926);
    nor g2444(n5870 ,n4651 ,n5760);
    nand g2445(n4324 ,n2603 ,n3885);
    xor g2446(n6034 ,n5940 ,n1507);
    or g2447(n2163 ,n719 ,n1584);
    nor g2448(n3294 ,n1954 ,n2856);
    nand g2449(n4264 ,n720 ,n3834);
    nand g2450(n3968 ,n0[6] ,n3490);
    or g2451(n9[69] ,n5676 ,n5923);
    not g2452(n5842 ,n5843);
    nor g2453(n4611 ,n727 ,n4479);
    not g2454(n2891 ,n2890);
    nor g2455(n6043 ,n713 ,n5971);
    xnor g2456(n6867 ,n93 ,n119);
    nor g2457(n4035 ,n3722 ,n3316);
    xnor g2458(n4465 ,n3938 ,n2820);
    nor g2459(n5900 ,n1954 ,n5752);
    nand g2460(n4823 ,n1966 ,n4468);
    nand g2461(n4683 ,n4131 ,n4379);
    nor g2462(n1054 ,n708 ,n0[5]);
    nand g2463(n5760 ,n5546 ,n5612);
    nor g2464(n4645 ,n711 ,n4467);
    xnor g2465(n1479 ,n1[73] ,n2[9]);
    nand g2466(n5382 ,n4822 ,n5145);
    or g2467(n3043 ,n2634 ,n2375);
    xnor g2468(n5207 ,n4882 ,n1501);
    nand g2469(n211 ,n0[50] ,n1[50]);
    nand g2470(n6519 ,n6485 ,n6495);
    nand g2471(n3133 ,n1493 ,n2602);
    nor g2472(n6582 ,n0[111] ,n0[79]);
    or g2473(n341 ,n7035 ,n7003);
    nor g2474(n3905 ,n6 ,n3492);
    nor g2475(n5788 ,n4053 ,n5682);
    nand g2476(n1162 ,n6844 ,n795);
    nor g2477(n6115 ,n706 ,n6068);
    nand g2478(n967 ,n790 ,n792);
    xnor g2479(n3944 ,n2687 ,n2836);
    not g2480(n712 ,n717);
    nand g2481(n9[65] ,n4038 ,n6488);
    xnor g2482(n4838 ,n4573 ,n4426);
    nand g2483(n6966 ,n6745 ,n6775);
    xnor g2484(n2660 ,n4[30] ,n1482);
    nand g2485(n133 ,n53 ,n132);
    not g2486(n814 ,n0[66]);
    xnor g2487(n1299 ,n1[59] ,n1[27]);
    xnor g2488(n89 ,n0[5] ,n7061);
    nand g2489(n3415 ,n1952 ,n2862);
    nor g2490(n6703 ,n6826 ,n6588);
    nor g2491(n6230 ,n3482 ,n6124);
    nor g2492(n5513 ,n5335 ,n5159);
    xnor g2493(n1267 ,n0[86] ,n7114);
    nor g2494(n4966 ,n3362 ,n4602);
    nor g2495(n2383 ,n0[27] ,n1963);
    nand g2496(n6222 ,n6149 ,n6072);
    xnor g2497(n1572 ,n0[4] ,n1[4]);
    nor g2498(n2133 ,n1961 ,n1468);
    xor g2499(n7108 ,n0[48] ,n0[16]);
    xnor g2500(n3943 ,n2691 ,n2802);
    nand g2501(n5539 ,n4705 ,n5312);
    nand g2502(n376 ,n7018 ,n6986);
    nand g2503(n4832 ,n1966 ,n4458);
    nor g2504(n5112 ,n4646 ,n5012);
    or g2505(n333 ,n7047 ,n7015);
    nor g2506(n5687 ,n3781 ,n5415);
    not g2507(n3503 ,n3502);
    nand g2508(n1206 ,n1[123] ,n2[59]);
    nor g2509(n2286 ,n1959 ,n1925);
    nand g2510(n6017 ,n4004 ,n5880);
    or g2511(n1737 ,n0[40] ,n991);
    nor g2512(n978 ,n724 ,n0[115]);
    nand g2513(n1148 ,n3[2] ,n783);
    nand g2514(n575 ,n519 ,n574);
    nor g2515(n5737 ,n711 ,n5587);
    nand g2516(n647 ,n0[89] ,n622);
    nand g2517(n6626 ,n1[74] ,n6579);
    nand g2518(n3282 ,n1952 ,n2871);
    nor g2519(n4012 ,n832 ,n3489);
    xnor g2520(n1290 ,n1[42] ,n4[2]);
    xnor g2521(n4410 ,n3810 ,n1968);
    or g2522(n3003 ,n2631 ,n2333);
    nor g2523(n3034 ,n2322 ,n2321);
    nor g2524(n5489 ,n4783 ,n5385);
    nand g2525(n10[7] ,n4615 ,n5319);
    nand g2526(n4940 ,n3542 ,n4725);
    xnor g2527(n3816 ,n1[91] ,n2708);
    nor g2528(n1749 ,n0[34] ,n1233);
    xnor g2529(n6849 ,n393 ,n415);
    nand g2530(n1796 ,n0[41] ,n1221);
    nand g2531(n3680 ,n3148 ,n2255);
    xnor g2532(n6930 ,n230 ,n303);
    nand g2533(n3602 ,n0[20] ,n2794);
    xnor g2534(n1366 ,n7092 ,n7050);
    or g2535(n2977 ,n2174 ,n2206);
    xnor g2536(n2940 ,n1609 ,n1573);
    nand g2537(n3349 ,n1952 ,n2902);
    xnor g2538(n2705 ,n0[52] ,n1967);
    nand g2539(n3767 ,n7131 ,n3068);
    nand g2540(n4517 ,n2009 ,n4362);
    nand g2541(n4268 ,n0[81] ,n3847);
    nor g2542(n5419 ,n706 ,n5244);
    nand g2543(n3325 ,n1953 ,n2887);
    nor g2544(n5522 ,n4966 ,n5292);
    not g2545(n1955 ,n711);
    nand g2546(n5045 ,n4691 ,n4872);
    or g2547(n7091 ,n3[3] ,n3[0]);
    xnor g2548(n252 ,n1[48] ,n0[48]);
    nor g2549(n2434 ,n721 ,n1508);
    nand g2550(n4519 ,n3677 ,n4300);
    nand g2551(n2028 ,n714 ,n998);
    nand g2552(n4110 ,n3243 ,n3575);
    nand g2553(n4155 ,n3483 ,n3925);
    nand g2554(n1066 ,n0[124] ,n709);
    nor g2555(n4944 ,n722 ,n4681);
    not g2556(n2008 ,n2007);
    nand g2557(n3277 ,n1953 ,n2860);
    not g2558(n5191 ,n5190);
    or g2559(n3316 ,n2746 ,n2218);
    not g2560(n768 ,n0[78]);
    nand g2561(n1133 ,n6951 ,n797);
    not g2562(n746 ,n0[114]);
    nor g2563(n1780 ,n0[45] ,n965);
    nand g2564(n7078 ,n664 ,n632);
    nor g2565(n5962 ,n5535 ,n5869);
    xnor g2566(n6510 ,n6413 ,n6306);
    nand g2567(n4281 ,n720 ,n3823);
    not g2568(n5976 ,n5977);
    nand g2569(n6467 ,n5779 ,n6431);
    nand g2570(n4067 ,n3604 ,n3636);
    nand g2571(n1975 ,n1080 ,n1210);
    nand g2572(n3591 ,n0[110] ,n2794);
    not g2573(n4895 ,n4894);
    or g2574(n3018 ,n2181 ,n2264);
    nand g2575(n6448 ,n3334 ,n6326);
    nor g2576(n2635 ,n0[23] ,n721);
    xnor g2577(n6217 ,n6032 ,n6109);
    nand g2578(n3987 ,n3591 ,n3097);
    nand g2579(n4541 ,n1156 ,n4137);
    or g2580(n2397 ,n1963 ,n1571);
    nand g2581(n4522 ,n4073 ,n4308);
    not g2582(n3263 ,n3234);
    or g2583(n5256 ,n4156 ,n5187);
    nand g2584(n7038 ,n6656 ,n7135);
    nand g2585(n4789 ,n845 ,n4433);
    nand g2586(n4347 ,n823 ,n4078);
    nand g2587(n4269 ,n2064 ,n3968);
    nor g2588(n1046 ,n725 ,n0[16]);
    nand g2589(n4017 ,n3622 ,n3491);
    xnor g2590(n1615 ,n0[71] ,n1[71]);
    nand g2591(n3720 ,n3172 ,n2748);
    nand g2592(n3467 ,n3117 ,n3118);
    nand g2593(n6613 ,n1[69] ,n6579);
    nor g2594(n2360 ,n0[116] ,n1956);
    nand g2595(n215 ,n0[40] ,n1[40]);
    xnor g2596(n6424 ,n6248 ,n6306);
    nand g2597(n3774 ,n1162 ,n3171);
    nand g2598(n3645 ,n0[55] ,n2796);
    nand g2599(n3769 ,n1219 ,n2741);
    nor g2600(n2322 ,n1961 ,n1392);
    or g2601(n2084 ,n1960 ,n1407);
    nor g2602(n5439 ,n5188 ,n5261);
    nand g2603(n1788 ,n1239 ,n1224);
    nor g2604(n2214 ,n1957 ,n1614);
    or g2605(n2784 ,n2196 ,n2118);
    nand g2606(n5035 ,n4964 ,n4887);
    nand g2607(n1942 ,n1227 ,n968);
    nand g2608(n4084 ,n3624 ,n3683);
    xnor g2609(n5057 ,n4590 ,n4452);
    nand g2610(n6809 ,n6581 ,n7105);
    nor g2611(n3253 ,n0[40] ,n2409);
    nand g2612(n9[35] ,n5113 ,n6547);
    nand g2613(n310 ,n170 ,n309);
    nor g2614(n4618 ,n4356 ,n4507);
    nand g2615(n608 ,n480 ,n607);
    or g2616(n5413 ,n706 ,n5374);
    xor g2617(n5285 ,n4670 ,n5004);
    not g2618(n4886 ,n4885);
    nor g2619(n2738 ,n1574 ,n2612);
    nor g2620(n3315 ,n1748 ,n3028);
    nor g2621(n4653 ,n6 ,n4452);
    nand g2622(n5789 ,n3625 ,n5647);
    nand g2623(n3647 ,n3133 ,n2762);
    or g2624(n2129 ,n719 ,n1563);
    nor g2625(n6523 ,n1954 ,n6463);
    not g2626(n838 ,n1[43]);
    xnor g2627(n6863 ,n92 ,n117);
    or g2628(n4740 ,n3532 ,n4555);
    nand g2629(n4930 ,n1955 ,n4658);
    xnor g2630(n5431 ,n4843 ,n5015);
    nand g2631(n4285 ,n2132 ,n4006);
    nand g2632(n3603 ,n0[21] ,n2794);
    nand g2633(n3783 ,n6818 ,n3235);
    nand g2634(n415 ,n362 ,n414);
    nor g2635(n2272 ,n1959 ,n1433);
    nand g2636(n1237 ,n0[70] ,n715);
    xnor g2637(n559 ,n6972 ,n0[115]);
    not g2638(n822 ,n0[49]);
    or g2639(n6036 ,n706 ,n5970);
    nand g2640(n3758 ,n7139 ,n3055);
    nor g2641(n4218 ,n3562 ,n3907);
    nand g2642(n6987 ,n6695 ,n6821);
    nand g2643(n43 ,n7085 ,n0[29]);
    nor g2644(n5176 ,n6824 ,n4901);
    xnor g2645(n4455 ,n3940 ,n2806);
    xnor g2646(n1489 ,n0[29] ,n1[29]);
    xnor g2647(n545 ,n6958 ,n0[101]);
    nor g2648(n3333 ,n1954 ,n2870);
    nor g2649(n2613 ,n0[4] ,n721);
    nand g2650(n3235 ,n1205 ,n2294);
    nand g2651(n5486 ,n5129 ,n5298);
    nand g2652(n4765 ,n2560 ,n4439);
    not g2653(n1245 ,n1244);
    nand g2654(n3268 ,n1952 ,n2855);
    nand g2655(n1910 ,n1095 ,n1016);
    xnor g2656(n1516 ,n0[83] ,n4[27]);
    not g2657(n2025 ,n2024);
    nand g2658(n5829 ,n5554 ,n5701);
    xnor g2659(n3838 ,n2688 ,n2683);
    nand g2660(n2607 ,n0[17] ,n1964);
    nor g2661(n5697 ,n5504 ,n5506);
    nand g2662(n3402 ,n1953 ,n2922);
    xnor g2663(n1491 ,n0[18] ,n1[18]);
    nand g2664(n3222 ,n1131 ,n2190);
    nand g2665(n6357 ,n6270 ,n6276);
    nor g2666(n1854 ,n755 ,n1220);
    xnor g2667(n1485 ,n0[31] ,n1[31]);
    or g2668(n481 ,n0[126] ,n6983);
    not g2669(n5835 ,n5836);
    nand g2670(n2509 ,n794 ,n2000);
    nor g2671(n6706 ,n6826 ,n6597);
    nor g2672(n4807 ,n2267 ,n4472);
    nor g2673(n4786 ,n4027 ,n4515);
    xor g2674(n7118 ,n0[58] ,n0[26]);
    nand g2675(n5022 ,n715 ,n5013);
    nor g2676(n5967 ,n1954 ,n5866);
    nor g2677(n6047 ,n5892 ,n5979);
    nor g2678(n4314 ,n4057 ,n3693);
    nor g2679(n2171 ,n1961 ,n1400);
    nor g2680(n3563 ,n709 ,n3258);
    nand g2681(n9[32] ,n4647 ,n6515);
    nand g2682(n5529 ,n4391 ,n5305);
    xnor g2683(n1707 ,n6906 ,n6907);
    nand g2684(n3302 ,n1952 ,n2874);
    nor g2685(n2291 ,n1961 ,n1924);
    nor g2686(n2781 ,n1728 ,n2510);
    nor g2687(n6134 ,n5883 ,n6059);
    or g2688(n2211 ,n719 ,n1629);
    nor g2689(n2324 ,n1961 ,n1389);
    nor g2690(n6286 ,n6227 ,n6199);
    nand g2691(n1145 ,n6873 ,n797);
    nand g2692(n3998 ,n710 ,n3799);
    nand g2693(n5361 ,n3807 ,n5142);
    nand g2694(n6098 ,n3375 ,n5952);
    nor g2695(n5229 ,n3284 ,n5090);
    nor g2696(n3087 ,n1221 ,n2391);
    nand g2697(n499 ,n0[125] ,n6982);
    nor g2698(n4987 ,n3271 ,n4703);
    nor g2699(n3475 ,n1954 ,n2943);
    nand g2700(n1187 ,n6857 ,n795);
    nor g2701(n1781 ,n0[41] ,n1017);
    nand g2702(n1911 ,n750 ,n1247);
    nor g2703(n1865 ,n809 ,n971);
    nand g2704(n4693 ,n717 ,n4579);
    not g2705(n813 ,n0[99]);
    nand g2706(n3709 ,n2079 ,n3183);
    not g2707(n747 ,n0[35]);
    nor g2708(n3781 ,n1954 ,n2952);
    nor g2709(n4984 ,n3567 ,n4710);
    nor g2710(n4203 ,n2325 ,n4101);
    nor g2711(n4523 ,n3692 ,n4305);
    xnor g2712(n2909 ,n1648 ,n1532);
    xnor g2713(n1407 ,n1[23] ,n2[23]);
    xnor g2714(n1585 ,n0[101] ,n1[101]);
    nand g2715(n5193 ,n4241 ,n4934);
    nor g2716(n1991 ,n871 ,n932);
    nor g2717(n3454 ,n789 ,n3259);
    not g2718(n844 ,n0[44]);
    nand g2719(n3237 ,n1207 ,n2144);
    nand g2720(n6677 ,n0[91] ,n6580);
    nand g2721(n3343 ,n1952 ,n2954);
    nand g2722(n6820 ,n6581 ,n7094);
    or g2723(n322 ,n7046 ,n7014);
    nor g2724(n3317 ,n1954 ,n2882);
    nand g2725(n4102 ,n3690 ,n3430);
    nor g2726(n3559 ,n3125 ,n3130);
    xnor g2727(n1380 ,n0[1] ,n4[17]);
    nand g2728(n3166 ,n1974 ,n2326);
    or g2729(n3908 ,n2377 ,n3490);
    not g2730(n1553 ,n1552);
    nor g2731(n3482 ,n1954 ,n2949);
    nand g2732(n3113 ,n1561 ,n2584);
    nand g2733(n3754 ,n7145 ,n3062);
    xnor g2734(n1948 ,n1[96] ,n2[32]);
    nor g2735(n3382 ,n2383 ,n3119);
    nand g2736(n279 ,n197 ,n278);
    nor g2737(n5800 ,n5190 ,n5626);
    xnor g2738(n1413 ,n1[19] ,n2[19]);
    nand g2739(n3234 ,n1126 ,n2183);
    nor g2740(n3801 ,n0[83] ,n3103);
    nand g2741(n6790 ,n1[115] ,n7088);
    or g2742(n3095 ,n2613 ,n2381);
    nand g2743(n3160 ,n2573 ,n2447);
    nand g2744(n5913 ,n5815 ,n5486);
    nor g2745(n1797 ,n733 ,n11);
    nand g2746(n5252 ,n708 ,n5074);
    nand g2747(n4393 ,n793 ,n4223);
    nand g2748(n6756 ,n0[34] ,n6737);
    nand g2749(n3713 ,n2222 ,n3194);
    nor g2750(n4302 ,n2757 ,n3928);
    nor g2751(n2384 ,n0[54] ,n719);
    nand g2752(n9[47] ,n5763 ,n5795);
    nor g2753(n6088 ,n3478 ,n5957);
    nand g2754(n1853 ,n0[33] ,n1221);
    nor g2755(n3892 ,n715 ,n3520);
    nor g2756(n3572 ,n2325 ,n3249);
    or g2757(n3861 ,n2320 ,n3706);
    nand g2758(n7067 ,n662 ,n630);
    nand g2759(n4585 ,n2523 ,n4232);
    nand g2760(n603 ,n502 ,n602);
    nor g2761(n6587 ,n0[110] ,n0[78]);
    xnor g2762(n5851 ,n5572 ,n1725);
    xnor g2763(n1350 ,n0[5] ,n4[21]);
    nand g2764(n6493 ,n6448 ,n6421);
    nor g2765(n5042 ,n727 ,n4902);
    xnor g2766(n1928 ,n1[122] ,n2[58]);
    nand g2767(n9[31] ,n5331 ,n5399);
    xnor g2768(n1408 ,n1[22] ,n2[22]);
    or g2769(n6298 ,n6155 ,n6210);
    xnor g2770(n5578 ,n1291 ,n5204);
    nand g2771(n10[19] ,n4767 ,n5339);
    or g2772(n24 ,n7081 ,n0[25]);
    xnor g2773(n2708 ,n1[123] ,n1299);
    nor g2774(n5299 ,n3531 ,n5041);
    xnor g2775(n1256 ,n6938 ,n6937);
    nand g2776(n10[10] ,n4769 ,n5346);
    xnor g2777(n82 ,n0[29] ,n7085);
    nand g2778(n3092 ,n11 ,n2395);
    nor g2779(n1051 ,n0[111] ,n715);
    nand g2780(n4088 ,n7149 ,n3422);
    nand g2781(n5630 ,n3270 ,n693);
    nand g2782(n143 ,n65 ,n142);
    nand g2783(n5400 ,n5102 ,n5264);
    not g2784(n793 ,n6);
    nand g2785(n423 ,n367 ,n422);
    xnor g2786(n1341 ,n6922 ,n6923);
    nand g2787(n454 ,n323 ,n453);
    nand g2788(n4095 ,n7135 ,n3668);
    not g2789(n3249 ,n3248);
    nor g2790(n4780 ,n726 ,n4438);
    nor g2791(n6169 ,n5797 ,n6039);
    not g2792(n818 ,n0[19]);
    nor g2793(n3305 ,n1954 ,n2876);
    or g2794(n3521 ,n6825 ,n2854);
    nor g2795(n4236 ,n2722 ,n3986);
    nor g2796(n2237 ,n1959 ,n1385);
    nor g2797(n1783 ,n0[32] ,n947);
    nor g2798(n861 ,n709 ,n0[39]);
    not g2799(n6802 ,n7156);
    xnor g2800(n1447 ,n1[112] ,n2[48]);
    nor g2801(n5811 ,n4758 ,n5696);
    nand g2802(n4065 ,n2752 ,n3665);
    or g2803(n6066 ,n4385 ,n5981);
    nand g2804(n6526 ,n6482 ,n6497);
    nand g2805(n6394 ,n5550 ,n6319);
    nand g2806(n3777 ,n7124 ,n2761);
    nor g2807(n6170 ,n5658 ,n6069);
    nand g2808(n592 ,n493 ,n591);
    nor g2809(n3272 ,n2330 ,n2796);
    nor g2810(n3291 ,n0[48] ,n3252);
    nor g2811(n5998 ,n3305 ,n5861);
    not g2812(n4462 ,n4461);
    or g2813(n5665 ,n4397 ,n5477);
    nor g2814(n2742 ,n2108 ,n2188);
    nor g2815(n5957 ,n713 ,n5935);
    nand g2816(n5982 ,n717 ,n5934);
    xnor g2817(n6044 ,n5848 ,n4101);
    nor g2818(n5883 ,n712 ,n5751);
    nand g2819(n633 ,n0[76] ,n622);
    nor g2820(n5462 ,n4192 ,n5272);
    nand g2821(n6745 ,n0[45] ,n6737);
    nor g2822(n5275 ,n4086 ,n5047);
    nand g2823(n433 ,n351 ,n432);
    xnor g2824(n405 ,n7003 ,n7035);
    xor g2825(n2688 ,n0[54] ,n1972);
    nand g2826(n6132 ,n6053 ,n6057);
    nand g2827(n10[20] ,n4761 ,n5340);
    nand g2828(n2749 ,n1562 ,n2638);
    nand g2829(n6566 ,n4153 ,n6548);
    nor g2830(n3100 ,n1858 ,n2226);
    nand g2831(n869 ,n801 ,n742);
    nor g2832(n5029 ,n722 ,n5010);
    nand g2833(n3129 ,n1[49] ,n2632);
    nor g2834(n3901 ,n2246 ,n3749);
    nor g2835(n5143 ,n727 ,n4912);
    nand g2836(n6471 ,n6290 ,n6417);
    nor g2837(n6029 ,n4487 ,n5886);
    nand g2838(n3986 ,n2468 ,n3543);
    nor g2839(n905 ,n1[65] ,n2[1]);
    nand g2840(n5384 ,n5131 ,n4759);
    nand g2841(n44 ,n7084 ,n0[28]);
    nor g2842(n2108 ,n1960 ,n1412);
    xnor g2843(n5392 ,n1273 ,n5065);
    nor g2844(n2751 ,n2071 ,n2070);
    nand g2845(n200 ,n0[49] ,n1[49]);
    not g2846(n6111 ,n6110);
    nor g2847(n6299 ,n6230 ,n6201);
    nor g2848(n5503 ,n722 ,n5375);
    nor g2849(n6242 ,n4200 ,n6144);
    or g2850(n469 ,n0[115] ,n6972);
    or g2851(n4969 ,n4306 ,n4800);
    or g2852(n168 ,n0[52] ,n1[52]);
    or g2853(n2465 ,n1961 ,n1444);
    or g2854(n2208 ,n1961 ,n1936);
    nor g2855(n3350 ,n1954 ,n2901);
    nand g2856(n992 ,n0[58] ,n714);
    nor g2857(n6171 ,n4751 ,n6070);
    nand g2858(n2511 ,n794 ,n1985);
    xnor g2859(n3960 ,n2824 ,n2842);
    or g2860(n9[11] ,n5344 ,n6577);
    nor g2861(n3429 ,n2266 ,n3018);
    nor g2862(n5136 ,n4969 ,n5012);
    nand g2863(n7128 ,n6675 ,n6724);
    nor g2864(n2095 ,n789 ,n1461);
    nand g2865(n6772 ,n1[107] ,n7088);
    not g2866(n6423 ,n6422);
    nand g2867(n6504 ,n6460 ,n6435);
    xnor g2868(n5204 ,n1360 ,n4838);
    or g2869(n6328 ,n713 ,n6307);
    xnor g2870(n6877 ,n400 ,n429);
    nor g2871(n6041 ,n712 ,n5972);
    nand g2872(n6696 ,n0[120] ,n0[88]);
    nor g2873(n6438 ,n3547 ,n6347);
    xnor g2874(n2684 ,n1[102] ,n1514);
    nor g2875(n1778 ,n0[13] ,n967);
    not g2876(n1566 ,n1565);
    nand g2877(n5432 ,n3287 ,n5287);
    nand g2878(n3558 ,n787 ,n2924);
    or g2879(n6046 ,n5891 ,n5980);
    nand g2880(n9[119] ,n5875 ,n6147);
    xnor g2881(n6312 ,n1580 ,n6195);
    nand g2882(n3208 ,n1171 ,n2129);
    nor g2883(n6609 ,n0[104] ,n0[72]);
    nor g2884(n1821 ,n738 ,n1220);
    nand g2885(n10[17] ,n4760 ,n5337);
    not g2886(n1483 ,n1482);
    nand g2887(n6450 ,n3786 ,n6329);
    nor g2888(n5651 ,n4870 ,n5539);
    nand g2889(n916 ,n0[41] ,n743);
    nor g2890(n6173 ,n4652 ,n6070);
    nand g2891(n2557 ,n1153 ,n1840);
    nand g2892(n6030 ,n4011 ,n5865);
    not g2893(n5261 ,n5262);
    nor g2894(n1757 ,n0[25] ,n1228);
    nand g2895(n3069 ,n714 ,n2139);
    nor g2896(n3613 ,n772 ,n2972);
    nor g2897(n5514 ,n4714 ,n5381);
    nand g2898(n7017 ,n6668 ,n7156);
    xnor g2899(n77 ,n0[24] ,n7080);
    xnor g2900(n1302 ,n0[79] ,n7107);
    nor g2901(n3051 ,n1797 ,n2150);
    or g2902(n4400 ,n0[24] ,n4233);
    xnor g2903(n2822 ,n1664 ,n1381);
    nor g2904(n3457 ,n1954 ,n2936);
    nor g2905(n2715 ,n2619 ,n2338);
    nor g2906(n6097 ,n6000 ,n5990);
    or g2907(n475 ,n0[120] ,n6977);
    or g2908(n3046 ,n1237 ,n2325);
    xor g2909(n7110 ,n0[50] ,n0[18]);
    nand g2910(n674 ,n1[1] ,n621);
    or g2911(n2130 ,n719 ,n1500);
    nand g2912(n5128 ,n715 ,n5011);
    nor g2913(n2723 ,n1963 ,n2441);
    or g2914(n316 ,n7029 ,n6997);
    nor g2915(n1771 ,n725 ,n1037);
    nor g2916(n3731 ,n3262 ,n3212);
    nand g2917(n4343 ,n3714 ,n3899);
    nand g2918(n71 ,n7067 ,n0[11]);
    nor g2919(n5656 ,n3273 ,n693);
    nor g2920(n2631 ,n0[29] ,n721);
    or g2921(n4133 ,n1960 ,n3921);
    nor g2922(n6585 ,n0[107] ,n0[75]);
    or g2923(n3918 ,n2342 ,n3490);
    xnor g2924(n5271 ,n4664 ,n4874);
    xnor g2925(n1687 ,n0[42] ,n0[26]);
    nand g2926(n4051 ,n715 ,n3523);
    nand g2927(n1183 ,n6920 ,n795);
    nand g2928(n6554 ,n4407 ,n6524);
    nor g2929(n4633 ,n3508 ,n4553);
    nand g2930(n4241 ,n1966 ,n3940);
    nand g2931(n4257 ,n715 ,n3965);
    nor g2932(n2393 ,n0[58] ,n1958);
    or g2933(n256 ,n224 ,n173);
    nand g2934(n132 ,n22 ,n131);
    nor g2935(n6370 ,n3295 ,n6258);
    nor g2936(n1761 ,n998 ,n873);
    nor g2937(n3089 ,n1221 ,n2361);
    nand g2938(n4342 ,n3601 ,n3977);
    nor g2939(n5138 ,n727 ,n4901);
    nor g2940(n5028 ,n6 ,n5005);
    not g2941(n1531 ,n1530);
    nand g2942(n4563 ,n7133 ,n4353);
    xnor g2943(n2697 ,n0[125] ,n1520);
    nand g2944(n889 ,n0[17] ,n801);
    nand g2945(n7072 ,n670 ,n643);
    xnor g2946(n6889 ,n403 ,n435);
    xnor g2947(n5567 ,n4844 ,n5379);
    nand g2948(n7069 ,n666 ,n634);
    nor g2949(n2981 ,n724 ,n2243);
    xnor g2950(n1441 ,n1[71] ,n2[7]);
    nand g2951(n9[24] ,n6529 ,n6392);
    or g2952(n5905 ,n4519 ,n5793);
    or g2953(n4617 ,n2561 ,n4464);
    nand g2954(n4955 ,n3319 ,n4755);
    nand g2955(n7023 ,n6613 ,n7150);
    nor g2956(n2157 ,n986 ,n1742);
    nand g2957(n4971 ,n4042 ,n4754);
    nor g2958(n2218 ,n1961 ,n1475);
    xnor g2959(n1276 ,n6858 ,n6859);
    nand g2960(n5749 ,n717 ,n5639);
    nor g2961(n2299 ,n1959 ,n1478);
    nand g2962(n373 ,n7021 ,n6989);
    nand g2963(n3122 ,n828 ,n2577);
    nor g2964(n2619 ,n0[2] ,n721);
    nand g2965(n6379 ,n3277 ,n6264);
    xnor g2966(n2843 ,n1379 ,n1712);
    xnor g2967(n5723 ,n5455 ,n1607);
    or g2968(n321 ,n7045 ,n7013);
    nor g2969(n2387 ,n0[31] ,n721);
    nor g2970(n4804 ,n3495 ,n4496);
    or g2971(n317 ,n7037 ,n7005);
    nor g2972(n2166 ,n949 ,n1961);
    nor g2973(n4613 ,n727 ,n4478);
    nor g2974(n3021 ,n2275 ,n2274);
    xnor g2975(n4596 ,n4108 ,n4219);
    nand g2976(n199 ,n0[45] ,n1[45]);
    nand g2977(n111 ,n58 ,n110);
    nand g2978(n515 ,n0[114] ,n6971);
    nand g2979(n4071 ,n3134 ,n3712);
    nand g2980(n5601 ,n3376 ,n5411);
    nor g2981(n2424 ,n1958 ,n1626);
    nor g2982(n2430 ,n1[63] ,n1484);
    nor g2983(n864 ,n708 ,n0[63]);
    or g2984(n2170 ,n1962 ,n1426);
    nand g2985(n522 ,n0[105] ,n6962);
    nor g2986(n2104 ,n1959 ,n1404);
    or g2987(n692 ,n4697 ,n5050);
    nand g2988(n348 ,n7046 ,n7014);
    nand g2989(n1846 ,n0[126] ,n966);
    xnor g2990(n2654 ,n1264 ,n1594);
    or g2991(n4616 ,n2561 ,n4463);
    nand g2992(n3184 ,n2563 ,n2494);
    or g2993(n4723 ,n712 ,n4568);
    nor g2994(n5873 ,n706 ,n5841);
    xnor g2995(n1454 ,n1[98] ,n2[34]);
    or g2996(n2113 ,n1960 ,n1928);
    nor g2997(n3852 ,n1776 ,n3363);
    nor g2998(n5479 ,n4645 ,n5289);
    nor g2999(n2013 ,n0[96] ,n1042);
    nand g3000(n1194 ,n6856 ,n795);
    nor g3001(n2282 ,n1963 ,n1523);
    not g3002(n5292 ,n5291);
    nand g3003(n4580 ,n2511 ,n4216);
    nand g3004(n420 ,n339 ,n419);
    nand g3005(n9[74] ,n5680 ,n6133);
    xnor g3006(n1336 ,n0[78] ,n4[6]);
    xnor g3007(n537 ,n6981 ,n0[124]);
    nor g3008(n6077 ,n6011 ,n5985);
    or g3009(n4622 ,n2561 ,n4451);
    nor g3010(n3884 ,n2341 ,n3490);
    or g3011(n175 ,n0[45] ,n1[45]);
    xnor g3012(n1552 ,n1[28] ,n828);
    nor g3013(n4299 ,n2325 ,n4100);
    nor g3014(n6262 ,n711 ,n6242);
    nor g3015(n3513 ,n6825 ,n2851);
    xnor g3016(n1287 ,n0[123] ,n4[11]);
    nor g3017(n3642 ,n777 ,n3039);
    or g3018(n34 ,n7066 ,n0[10]);
    nand g3019(n4013 ,n0[70] ,n3490);
    or g3020(n2119 ,n719 ,n1489);
    nand g3021(n7020 ,n6699 ,n7153);
    nand g3022(n440 ,n341 ,n439);
    nor g3023(n3331 ,n1[41] ,n3142);
    nor g3024(n6596 ,n0[119] ,n0[87]);
    nor g3025(n6375 ,n3554 ,n6262);
    nor g3026(n851 ,n0[43] ,n0[42]);
    nand g3027(n5740 ,n1953 ,n5578);
    xnor g3028(n2663 ,n1[106] ,n1512);
    nand g3029(n3983 ,n1965 ,n3589);
    or g3030(n4687 ,n1965 ,n4449);
    or g3031(n9[63] ,n4343 ,n5813);
    xor g3032(n7051 ,n0[97] ,n0[65]);
    nor g3033(n941 ,n822 ,n723);
    nor g3034(n5233 ,n3473 ,n5194);
    nor g3035(n4247 ,n1960 ,n3833);
    nor g3036(n3672 ,n3143 ,n2996);
    nand g3037(n4048 ,n3630 ,n2211);
    or g3038(n4168 ,n2136 ,n3872);
    xnor g3039(n3813 ,n0[76] ,n2659);
    nand g3040(n4650 ,n1041 ,n4400);
    xnor g3041(n381 ,n7010 ,n7042);
    or g3042(n3303 ,n2740 ,n2734);
    nand g3043(n5825 ,n4389 ,n5657);
    nor g3044(n6234 ,n3481 ,n6128);
    nand g3045(n275 ,n222 ,n274);
    or g3046(n4142 ,n3367 ,n4080);
    nand g3047(n3967 ,n0[69] ,n3490);
    nor g3048(n2651 ,n2233 ,n2112);
    nand g3049(n6664 ,n0[93] ,n6579);
    xnor g3050(n1417 ,n1[18] ,n2[18]);
    nand g3051(n601 ,n498 ,n600);
    nand g3052(n6461 ,n5123 ,n6378);
    xnor g3053(n1445 ,n0[84] ,n0[68]);
    nand g3054(n887 ,n0[90] ,n724);
    xnor g3055(n5471 ,n4665 ,n5157);
    xnor g3056(n6876 ,n552 ,n581);
    nand g3057(n3375 ,n1953 ,n2912);
    nand g3058(n7075 ,n685 ,n652);
    nand g3059(n445 ,n368 ,n444);
    nand g3060(n6800 ,n1[105] ,n7088);
    or g3061(n2763 ,n1557 ,n2616);
    nor g3062(n3348 ,n1954 ,n2884);
    nand g3063(n4105 ,n3578 ,n3662);
    nand g3064(n4761 ,n2560 ,n4446);
    or g3065(n3012 ,n2249 ,n2248);
    not g3066(n5058 ,n5059);
    not g3067(n6203 ,n6202);
    nor g3068(n3553 ,n1954 ,n2898);
    xnor g3069(n2913 ,n1726 ,n1634);
    xnor g3070(n4594 ,n4222 ,n2808);
    nor g3071(n863 ,n791 ,n0[12]);
    xnor g3072(n3819 ,n2705 ,n2669);
    nand g3073(n1205 ,n1[4] ,n2[4]);
    or g3074(n3314 ,n1954 ,n2881);
    nand g3075(n360 ,n7034 ,n7002);
    not g3076(n2598 ,n2597);
    or g3077(n18 ,n7084 ,n0[28]);
    not g3078(n745 ,n0[88]);
    nor g3079(n2139 ,n0[107] ,n1730);
    nor g3080(n6331 ,n6255 ,n6256);
    nand g3081(n5187 ,n4241 ,n4987);
    nor g3082(n5671 ,n3366 ,n5429);
    nand g3083(n3378 ,n1953 ,n2872);
    nand g3084(n7164 ,n6581 ,n7115);
    nand g3085(n3588 ,n0[37] ,n2794);
    nand g3086(n2456 ,n0[75] ,n2020);
    nor g3087(n4847 ,n722 ,n4809);
    or g3088(n9[15] ,n5739 ,n6008);
    xnor g3089(n2694 ,n1[116] ,n1531);
    nor g3090(n5680 ,n4313 ,n5564);
    nand g3091(n573 ,n517 ,n572);
    nor g3092(n3362 ,n1954 ,n2905);
    or g3093(n6483 ,n5987 ,n6403);
    nand g3094(n5704 ,n4154 ,n5565);
    nand g3095(n1901 ,n0[41] ,n991);
    nand g3096(n6167 ,n6091 ,n6100);
    nor g3097(n5938 ,n4418 ,n5772);
    not g3098(n3954 ,n3953);
    nand g3099(n6813 ,n6581 ,n7101);
    nor g3100(n5337 ,n4743 ,n5165);
    nor g3101(n2411 ,n725 ,n1829);
    nor g3102(n2243 ,n903 ,n1747);
    nor g3103(n6704 ,n6826 ,n6590);
    nand g3104(n306 ,n193 ,n305);
    nand g3105(n5746 ,n5607 ,n5606);
    nand g3106(n2506 ,n1106 ,n1992);
    nor g3107(n2281 ,n1962 ,n1401);
    xnor g3108(n1941 ,n1[45] ,n2[45]);
    xnor g3109(n5069 ,n4661 ,n4579);
    nand g3110(n7153 ,n6581 ,n7052);
    not g3111(n4911 ,n4910);
    xnor g3112(n6421 ,n6311 ,n6243);
    nor g3113(n2412 ,n0[104] ,n1760);
    nand g3114(n7085 ,n656 ,n638);
    xnor g3115(n3959 ,n2838 ,n2829);
    nor g3116(n880 ,n0[119] ,n6);
    nor g3117(n2098 ,n1956 ,n1578);
    not g3118(n4227 ,n4226);
    nand g3119(n2523 ,n794 ,n1973);
    or g3120(n5672 ,n3744 ,n5545);
    nor g3121(n2103 ,n1957 ,n1641);
    nand g3122(n5099 ,n717 ,n4989);
    not g3123(n4990 ,n4989);
    nor g3124(n4154 ,n3773 ,n4065);
    nor g3125(n5350 ,n4719 ,n5162);
    xnor g3126(n1406 ,n1[63] ,n2[63]);
    xnor g3127(n1917 ,n1[100] ,n2[36]);
    not g3128(n3490 ,n3489);
    nand g3129(n4028 ,n991 ,n3265);
    nand g3130(n3723 ,n1161 ,n3046);
    nor g3131(n3891 ,n2244 ,n3741);
    nor g3132(n2787 ,n2146 ,n2131);
    nand g3133(n2078 ,n792 ,n2002);
    xnor g3134(n1384 ,n6837 ,n6836);
    nand g3135(n5364 ,n3504 ,n5146);
    nor g3136(n3377 ,n1954 ,n2872);
    nand g3137(n5556 ,n4817 ,n5234);
    nand g3138(n7160 ,n6581 ,n7119);
    nor g3139(n1727 ,n791 ,n910);
    xnor g3140(n2709 ,n1343 ,n1570);
    nand g3141(n261 ,n221 ,n260);
    nor g3142(n5156 ,n2283 ,n4883);
    xnor g3143(n231 ,n1[58] ,n0[58]);
    xnor g3144(n1477 ,n1[69] ,n2[5]);
    not g3145(n761 ,n0[20]);
    nor g3146(n1756 ,n1054 ,n945);
    nor g3147(n2045 ,n1961 ,n1418);
    xnor g3148(n1353 ,n0[17] ,n4[25]);
    nand g3149(n4363 ,n4019 ,n3923);
    nor g3150(n5342 ,n4626 ,n5176);
    nor g3151(n6289 ,n6228 ,n6198);
    nand g3152(n6449 ,n3379 ,n6327);
    nand g3153(n2003 ,n962 ,n924);
    nand g3154(n6618 ,n0[82] ,n6579);
    not g3155(n1006 ,n1005);
    nor g3156(n3488 ,n1222 ,n2804);
    xnor g3157(n5430 ,n5059 ,n4210);
    nor g3158(n5182 ,n3428 ,n4880);
    xnor g3159(n4433 ,n2831 ,n3956);
    nor g3160(n2154 ,n1961 ,n1479);
    nor g3161(n4271 ,n2325 ,n4107);
    not g3162(n708 ,n715);
    nor g3163(n5705 ,n5371 ,n5473);
    not g3164(n2938 ,n2937);
    xnor g3165(n6413 ,n6308 ,n6174);
    not g3166(n4828 ,n4827);
    nor g3167(n4598 ,n722 ,n4456);
    nor g3168(n3053 ,n1800 ,n2195);
    nor g3169(n3058 ,n1823 ,n2161);
    xnor g3170(n1563 ,n0[14] ,n1[14]);
    not g3171(n841 ,n1[53]);
    nor g3172(n6607 ,n0[120] ,n0[88]);
    nor g3173(n5546 ,n4834 ,n5363);
    nor g3174(n4691 ,n713 ,n4579);
    nand g3175(n9[67] ,n4040 ,n6570);
    nand g3176(n1247 ,n0[10] ,n0[8]);
    nor g3177(n2485 ,n1956 ,n1439);
    nor g3178(n4262 ,n710 ,n4110);
    nor g3179(n1856 ,n757 ,n1220);
    nand g3180(n5247 ,n4956 ,n5067);
    xnor g3181(n2646 ,n768 ,n1977);
    xor g3182(n6176 ,n6066 ,n1538);
    xnor g3183(n242 ,n1[38] ,n0[38]);
    xnor g3184(n5055 ,n4370 ,n4592);
    nor g3185(n2174 ,n1956 ,n1627);
    nand g3186(n4016 ,n3621 ,n3491);
    or g3187(n492 ,n0[108] ,n6965);
    nor g3188(n3108 ,n1875 ,n2319);
    xnor g3189(n1370 ,n6921 ,n6920);
    nand g3190(n6688 ,n0[79] ,n6580);
    nand g3191(n3604 ,n0[52] ,n2796);
    nor g3192(n2183 ,n860 ,n1960);
    nor g3193(n5340 ,n4625 ,n5174);
    nor g3194(n6432 ,n3408 ,n6333);
    nor g3195(n3550 ,n1[67] ,n2910);
    nor g3196(n2426 ,n807 ,n2012);
    nand g3197(n3204 ,n1154 ,n2239);
    or g3198(n5498 ,n4247 ,n5384);
    nor g3199(n5802 ,n5104 ,n5681);
    nor g3200(n2138 ,n874 ,n1998);
    xnor g3201(n6119 ,n5943 ,n4109);
    xnor g3202(n406 ,n7004 ,n7036);
    nand g3203(n1146 ,n6916 ,n797);
    nand g3204(n1170 ,n6833 ,n797);
    nand g3205(n145 ,n42 ,n144);
    xnor g3206(n1508 ,n0[25] ,n1[25]);
    nor g3207(n5867 ,n5802 ,n5764);
    nor g3208(n2972 ,n2637 ,n2340);
    nand g3209(n2538 ,n1113 ,n1834);
    nor g3210(n2760 ,n2082 ,n2081);
    nand g3211(n456 ,n328 ,n455);
    nor g3212(n5254 ,n3299 ,n5051);
    nand g3213(n444 ,n317 ,n443);
    nand g3214(n1229 ,n0[104] ,n714);
    xnor g3215(n1272 ,n6929 ,n6928);
    xnor g3216(n1861 ,n0[43] ,n743);
    nor g3217(n4402 ,n3787 ,n4274);
    or g3218(n172 ,n0[48] ,n1[48]);
    xnor g3219(n4209 ,n3541 ,n1981);
    nor g3220(n3806 ,n1222 ,n2840);
    nor g3221(n2177 ,n850 ,n2011);
    nand g3222(n10[27] ,n4621 ,n5324);
    nand g3223(n634 ,n0[77] ,n622);
    nand g3224(n658 ,n1[9] ,n621);
    nand g3225(n4000 ,n0[116] ,n3335);
    nor g3226(n3102 ,n1862 ,n2438);
    nor g3227(n2462 ,n892 ,n1751);
    not g3228(n2626 ,n2625);
    nand g3229(n7025 ,n6619 ,n7148);
    nand g3230(n6351 ,n717 ,n6311);
    xnor g3231(n1355 ,n1[62] ,n1[30]);
    nand g3232(n6494 ,n6449 ,n6424);
    nor g3233(n2212 ,n1957 ,n1594);
    nor g3234(n911 ,n0[15] ,n0[7]);
    nand g3235(n5151 ,n6827 ,n4924);
    nand g3236(n3994 ,n0[14] ,n3491);
    nor g3237(n6712 ,n6826 ,n6582);
    nand g3238(n3345 ,n1952 ,n2897);
    xnor g3239(n6951 ,n83 ,n161);
    nor g3240(n5524 ,n4030 ,n5372);
    nand g3241(n5220 ,n4930 ,n5046);
    xnor g3242(n1637 ,n0[77] ,n1[77]);
    nor g3243(n4600 ,n712 ,n4577);
    nor g3244(n2375 ,n0[40] ,n1957);
    not g3245(n6340 ,n6339);
    xnor g3246(n6035 ,n4[8] ,n5932);
    nand g3247(n3684 ,n3150 ,n2421);
    nand g3248(n426 ,n338 ,n425);
    or g3249(n6441 ,n5381 ,n6356);
    nand g3250(n4758 ,n3614 ,n4509);
    xnor g3251(n384 ,n7013 ,n7045);
    nand g3252(n127 ,n45 ,n126);
    or g3253(n327 ,n7031 ,n6999);
    nand g3254(n4076 ,n3644 ,n3638);
    nand g3255(n4562 ,n1123 ,n4187);
    or g3256(n164 ,n0[43] ,n1[43]);
    nor g3257(n4222 ,n3560 ,n3902);
    nand g3258(n431 ,n349 ,n430);
    xnor g3259(n228 ,n1[55] ,n0[55]);
    nor g3260(n4119 ,n2798 ,n3938);
    xnor g3261(n4442 ,n2811 ,n3959);
    not g3262(n5721 ,n5698);
    nand g3263(n262 ,n166 ,n261);
    nand g3264(n6670 ,n0[86] ,n6579);
    not g3265(n6579 ,n6578);
    or g3266(n4306 ,n2541 ,n3871);
    or g3267(n4137 ,n1960 ,n3855);
    not g3268(n787 ,n710);
    nor g3269(n968 ,n725 ,n0[105]);
    nand g3270(n6492 ,n6447 ,n6416);
    nand g3271(n300 ,n190 ,n299);
    xnor g3272(n5202 ,n4425 ,n4836);
    nor g3273(n6082 ,n3323 ,n5958);
    nand g3274(n374 ,n7028 ,n6996);
    nor g3275(n3526 ,n6825 ,n2843);
    nand g3276(n3433 ,n1953 ,n2931);
    nand g3277(n5845 ,n4405 ,n5642);
    nor g3278(n4776 ,n727 ,n688);
    or g3279(n5436 ,n4248 ,n5389);
    nand g3280(n6329 ,n1955 ,n6280);
    or g3281(n496 ,n0[102] ,n6959);
    or g3282(n5110 ,n3730 ,n4950);
    nand g3283(n4999 ,n2060 ,n4673);
    nor g3284(n1037 ,n810 ,n0[75]);
    nor g3285(n4217 ,n3979 ,n3924);
    or g3286(n4167 ,n1961 ,n3910);
    nand g3287(n3585 ,n0[40] ,n2967);
    nand g3288(n2504 ,n1881 ,n1830);
    or g3289(n2999 ,n2622 ,n2393);
    nand g3290(n4157 ,n793 ,n4109);
    nor g3291(n6377 ,n5192 ,n6272);
    nand g3292(n3785 ,n6816 ,n3238);
    or g3293(n2754 ,n2094 ,n2214);
    nand g3294(n6159 ,n6092 ,n6080);
    nor g3295(n3874 ,n3215 ,n3661);
    nand g3296(n5225 ,n4713 ,n5120);
    xnor g3297(n1450 ,n1[104] ,n2[40]);
    nand g3298(n1859 ,n0[32] ,n1221);
    nand g3299(n582 ,n492 ,n581);
    nand g3300(n6101 ,n6028 ,n5991);
    xnor g3301(n1425 ,n1[10] ,n2[10]);
    xnor g3302(n549 ,n6962 ,n0[105]);
    nor g3303(n4866 ,n4145 ,n4703);
    not g3304(n780 ,n0[46]);
    xnor g3305(n2919 ,n1654 ,n1541);
    nor g3306(n2342 ,n1[85] ,n1956);
    nand g3307(n10[22] ,n4763 ,n5342);
    nor g3308(n6604 ,n0[127] ,n0[95]);
    nor g3309(n4418 ,n6 ,n4225);
    nand g3310(n1161 ,n6855 ,n796);
    xnor g3311(n1543 ,n0[49] ,n4[9]);
    nor g3312(n6369 ,n3276 ,n6257);
    nor g3313(n6094 ,n4520 ,n6024);
    nand g3314(n4783 ,n4041 ,n4486);
    nand g3315(n4571 ,n2525 ,n4224);
    nand g3316(n574 ,n489 ,n573);
    nor g3317(n3495 ,n6825 ,n2818);
    nor g3318(n1977 ,n878 ,n1086);
    nand g3319(n3200 ,n2005 ,n2124);
    nand g3320(n1158 ,n6945 ,n795);
    xnor g3321(n5979 ,n5845 ,n5463);
    nor g3322(n2748 ,n2104 ,n2103);
    nor g3323(n2146 ,n719 ,n1527);
    nor g3324(n5236 ,n3579 ,n5175);
    or g3325(n5807 ,n5602 ,n5560);
    not g3326(n809 ,n0[89]);
    not g3327(n4438 ,n4437);
    nand g3328(n4124 ,n3737 ,n3851);
    xnor g3329(n6881 ,n401 ,n431);
    nor g3330(n5178 ,n6824 ,n4927);
    nand g3331(n2428 ,n742 ,n1849);
    or g3332(n3032 ,n2305 ,n2304);
    nand g3333(n5817 ,n5707 ,n5667);
    xnor g3334(n1362 ,n6838 ,n6839);
    xnor g3335(n6865 ,n397 ,n423);
    not g3336(n621 ,n620);
    nand g3337(n6642 ,n1[79] ,n6580);
    or g3338(n4701 ,n1965 ,n4451);
    not g3339(n2596 ,n2595);
    nor g3340(n2161 ,n1957 ,n1616);
    nor g3341(n4132 ,n2445 ,n4097);
    or g3342(n3451 ,n791 ,n3259);
    nor g3343(n6725 ,n6826 ,n6601);
    nor g3344(n2248 ,n1962 ,n1398);
    xnor g3345(n80 ,n0[27] ,n7083);
    nand g3346(n5020 ,n3423 ,n4880);
    not g3347(n5480 ,n5479);
    or g3348(n4414 ,n4350 ,n4088);
    nor g3349(n3907 ,n789 ,n3794);
    nor g3350(n2105 ,n1962 ,n1464);
    xnor g3351(n2849 ,n1265 ,n1718);
    nand g3352(n7037 ,n6653 ,n7136);
    not g3353(n4367 ,n4366);
    nand g3354(n3576 ,n0[69] ,n2794);
    nand g3355(n563 ,n513 ,n562);
    nand g3356(n9[81] ,n5915 ,n6364);
    xnor g3357(n1248 ,n0[116] ,n4[4]);
    nor g3358(n6724 ,n6826 ,n6600);
    xnor g3359(n2928 ,n1615 ,n1510);
    not g3360(n796 ,n6826);
    nand g3361(n4337 ,n3653 ,n3863);
    or g3362(n3048 ,n1238 ,n2325);
    xnor g3363(n1511 ,n0[48] ,n4[8]);
    nand g3364(n1830 ,n0[6] ,n964);
    xnor g3365(n5725 ,n4683 ,n5528);
    nand g3366(n218 ,n0[41] ,n1[41]);
    nand g3367(n1105 ,n0[39] ,n708);
    xnor g3368(n1715 ,n1[6] ,n4[6]);
    xnor g3369(n1526 ,n0[7] ,n1[7]);
    nor g3370(n3101 ,n1856 ,n2250);
    or g3371(n706 ,n1232 ,n974);
    nand g3372(n6630 ,n0[107] ,n0[75]);
    nor g3373(n4965 ,n3369 ,n4606);
    nor g3374(n2089 ,n719 ,n1631);
    nand g3375(n6791 ,n1[124] ,n7088);
    or g3376(n4165 ,n3228 ,n3971);
    xnor g3377(n5594 ,n5199 ,n1307);
    xnor g3378(n2860 ,n1593 ,n1494);
    nor g3379(n2346 ,n0[87] ,n1956);
    xnor g3380(n4591 ,n4227 ,n3492);
    nand g3381(n3221 ,n1142 ,n2187);
    nand g3382(n4298 ,n720 ,n3822);
    nor g3383(n5339 ,n4649 ,n5159);
    xnor g3384(n5781 ,n5269 ,n5527);
    nand g3385(n3548 ,n1953 ,n2962);
    nand g3386(n153 ,n67 ,n152);
    nand g3387(n3148 ,n1[118] ,n2376);
    nor g3388(n5315 ,n4807 ,n5182);
    nor g3389(n4497 ,n3932 ,n4312);
    xnor g3390(n2921 ,n1599 ,n1511);
    nor g3391(n2629 ,n0[14] ,n721);
    nand g3392(n161 ,n43 ,n160);
    xnor g3393(n2713 ,n1[121] ,n1528);
    nand g3394(n2500 ,n0[91] ,n2018);
    nor g3395(n4192 ,n6 ,n3950);
    nor g3396(n3881 ,n715 ,n3517);
    nand g3397(n453 ,n356 ,n452);
    or g3398(n3401 ,n1954 ,n2922);
    nor g3399(n5490 ,n4691 ,n5355);
    nand g3400(n4798 ,n4499 ,n4488);
    nand g3401(n6627 ,n0[70] ,n6580);
    xnor g3402(n3812 ,n0[53] ,n2965);
    or g3403(n1904 ,n730 ,n983);
    or g3404(n9[50] ,n4522 ,n6185);
    xor g3405(n5286 ,n4669 ,n5008);
    nor g3406(n4661 ,n959 ,n4472);
    nor g3407(n4472 ,n793 ,n4212);
    xnor g3408(n4659 ,n4118 ,n1986);
    xor g3409(n695 ,n2670 ,n5271);
    nand g3410(n3654 ,n3136 ,n2774);
    not g3411(n2901 ,n2900);
    nor g3412(n5935 ,n4749 ,n5774);
    nor g3413(n3667 ,n818 ,n3087);
    or g3414(n4030 ,n3709 ,n3275);
    nor g3415(n2176 ,n872 ,n1871);
    nand g3416(n3386 ,n2088 ,n2765);
    nor g3417(n6575 ,n6542 ,n6572);
    nand g3418(n149 ,n52 ,n148);
    nand g3419(n2353 ,n1964 ,n1557);
    nand g3420(n2516 ,n794 ,n1989);
    nor g3421(n5101 ,n713 ,n4996);
    nor g3422(n5756 ,n5470 ,n5615);
    or g3423(n177 ,n0[62] ,n1[62]);
    nor g3424(n3697 ,n1[39] ,n3162);
    or g3425(n5929 ,n4337 ,n5807);
    nand g3426(n6264 ,n1955 ,n6249);
    xnor g3427(n5059 ,n4671 ,n4569);
    nand g3428(n4122 ,n2560 ,n3945);
    nand g3429(n2968 ,n938 ,n2276);
    nor g3430(n4398 ,n722 ,n4227);
    nand g3431(n417 ,n359 ,n416);
    nor g3432(n3259 ,n904 ,n2608);
    nand g3433(n359 ,n7023 ,n6991);
    nand g3434(n3763 ,n7136 ,n3067);
    or g3435(n2080 ,n719 ,n1538);
    nand g3436(n4996 ,n1069 ,n4679);
    xnor g3437(n1294 ,n0[12] ,n4[28]);
    nand g3438(n4320 ,n2607 ,n3915);
    nor g3439(n4994 ,n2514 ,n4675);
    nor g3440(n2724 ,n1241 ,n2606);
    xnor g3441(n2888 ,n1485 ,n1323);
    nand g3442(n3598 ,n0[101] ,n2794);
    nor g3443(n2296 ,n1961 ,n1919);
    nand g3444(n4520 ,n3674 ,n4302);
    nand g3445(n10[15] ,n4772 ,n5349);
    or g3446(n4301 ,n3718 ,n3854);
    nand g3447(n631 ,n0[91] ,n622);
    nand g3448(n7047 ,n6686 ,n7126);
    nor g3449(n2135 ,n1957 ,n1932);
    nand g3450(n3136 ,n1506 ,n2566);
    xnor g3451(n5730 ,n4665 ,n5454);
    xnor g3452(n6946 ,n234 ,n311);
    xnor g3453(n1399 ,n1[34] ,n2[34]);
    not g3454(n5642 ,n5641);
    nor g3455(n3267 ,n1954 ,n2857);
    nor g3456(n2193 ,n970 ,n1785);
    xnor g3457(n5581 ,n5262 ,n2679);
    nand g3458(n2510 ,n979 ,n1923);
    xnor g3459(n1262 ,n0[120] ,n0[88]);
    nand g3460(n6522 ,n6481 ,n6494);
    nand g3461(n6466 ,n6428 ,n6422);
    xnor g3462(n5850 ,n5573 ,n1294);
    nand g3463(n7042 ,n6667 ,n7131);
    nor g3464(n2722 ,n1007 ,n2450);
    nand g3465(n6302 ,n6160 ,n6210);
    nand g3466(n4275 ,n791 ,n4114);
    nand g3467(n5806 ,n5686 ,n5699);
    nand g3468(n6549 ,n1952 ,n705);
    nor g3469(n4024 ,n3210 ,n3386);
    xor g3470(n7117 ,n0[57] ,n0[25]);
    nand g3471(n6335 ,n1955 ,n6305);
    not g3472(n5980 ,n5979);
    xnor g3473(n5947 ,n5725 ,n4808);
    nand g3474(n3691 ,n843 ,n3157);
    nand g3475(n3695 ,n781 ,n3160);
    nand g3476(n295 ,n217 ,n294);
    xor g3477(n3823 ,n2684 ,n1[70]);
    nand g3478(n4782 ,n1799 ,n4518);
    nand g3479(n4961 ,n3389 ,n4777);
    nand g3480(n4956 ,n3565 ,n4756);
    nand g3481(n3199 ,n1968 ,n2326);
    xnor g3482(n1388 ,n1[57] ,n2[57]);
    nor g3483(n6567 ,n5920 ,n6544);
    or g3484(n560 ,n528 ,n477);
    nor g3485(n6037 ,n5735 ,n5949);
    nand g3486(n7004 ,n6618 ,n6804);
    nand g3487(n5268 ,n4161 ,n5063);
    nor g3488(n2127 ,n1960 ,n1443);
    nand g3489(n4797 ,n1835 ,n4526);
    nor g3490(n6251 ,n712 ,n6190);
    nor g3491(n6547 ,n5091 ,n6531);
    nand g3492(n5612 ,n5480 ,n5478);
    nand g3493(n3206 ,n1174 ,n2069);
    nor g3494(n6490 ,n6439 ,n6426);
    nand g3495(n146 ,n26 ,n145);
    xnor g3496(n1323 ,n0[15] ,n4[31]);
    nand g3497(n1179 ,n6900 ,n796);
    nor g3498(n5313 ,n3426 ,n5072);
    not g3499(n823 ,n0[11]);
    nor g3500(n6059 ,n1954 ,n5953);
    nand g3501(n4952 ,n3390 ,n4722);
    nand g3502(n5886 ,n5191 ,n5743);
    not g3503(n755 ,n0[104]);
    not g3504(n5986 ,n5985);
    not g3505(n966 ,n967);
    xor g3506(n687 ,n3946 ,n2849);
    nor g3507(n944 ,n747 ,n0[33]);
    nor g3508(n5677 ,n4414 ,n5539);
    nor g3509(n1785 ,n0[51] ,n1239);
    xnor g3510(n2683 ,n1990 ,n1987);
    or g3511(n4605 ,n706 ,n4570);
    xnor g3512(n6348 ,n6170 ,n6248);
    nand g3513(n5171 ,n4238 ,n4978);
    nand g3514(n638 ,n0[93] ,n622);
    nor g3515(n4731 ,n2325 ,n4460);
    nand g3516(n4621 ,n2560 ,n4450);
    not g3517(n2644 ,n2538);
    nand g3518(n9[127] ,n5052 ,n5812);
    xnor g3519(n2710 ,n1[97] ,n1260);
    xnor g3520(n6387 ,n6305 ,n2695);
    xnor g3521(n3855 ,n1[87] ,n2699);
    nand g3522(n4494 ,n794 ,n4360);
    nand g3523(n6633 ,n0[71] ,n6579);
    nand g3524(n7166 ,n6581 ,n7113);
    nor g3525(n4179 ,n3224 ,n4077);
    nor g3526(n5895 ,n711 ,n5837);
    nand g3527(n6973 ,n6762 ,n6796);
    not g3528(n719 ,n718);
    xnor g3529(n3947 ,n1334 ,n2827);
    not g3530(n749 ,n0[7]);
    nor g3531(n5115 ,n6 ,n5007);
    xnor g3532(n386 ,n7015 ,n7047);
    nand g3533(n2507 ,n792 ,n1969);
    nand g3534(n6782 ,n1[122] ,n7088);
    nand g3535(n3665 ,n0[10] ,n3080);
    xnor g3536(n2884 ,n1327 ,n1492);
    xnor g3537(n2801 ,n1371 ,n1707);
    xnor g3538(n380 ,n7009 ,n7041);
    nor g3539(n6142 ,n792 ,n6045);
    xnor g3540(n2858 ,n1697 ,n1632);
    nand g3541(n3327 ,n1952 ,n2884);
    nand g3542(n7077 ,n661 ,n628);
    nand g3543(n455 ,n358 ,n454);
    nand g3544(n10[16] ,n4773 ,n5350);
    nand g3545(n1117 ,n6868 ,n796);
    nor g3546(n2721 ,n931 ,n2107);
    nor g3547(n4662 ,n2232 ,n4471);
    xnor g3548(n1308 ,n6833 ,n6832);
    xnor g3549(n6879 ,n96 ,n125);
    nand g3550(n5383 ,n4690 ,n5133);
    nand g3551(n3717 ,n3166 ,n2787);
    nor g3552(n5662 ,n722 ,n5531);
    nand g3553(n3794 ,n933 ,n3163);
    nor g3554(n2643 ,n801 ,n1873);
    nor g3555(n5795 ,n4655 ,n5609);
    not g3556(n807 ,n0[107]);
    nand g3557(n3287 ,n1952 ,n2858);
    nor g3558(n4385 ,n6 ,n4226);
    nor g3559(n2337 ,n0[68] ,n1958);
    nand g3560(n5564 ,n4827 ,n5231);
    nand g3561(n6693 ,n0[64] ,n6580);
    xnor g3562(n1310 ,n6873 ,n6872);
    nor g3563(n3060 ,n1820 ,n2240);
    nand g3564(n6747 ,n0[46] ,n6737);
    xnor g3565(n6888 ,n555 ,n587);
    nand g3566(n6620 ,n0[69] ,n6579);
    or g3567(n182 ,n0[53] ,n1[53]);
    nor g3568(n6000 ,n3333 ,n5862);
    nor g3569(n1083 ,n842 ,n790);
    nor g3570(n5798 ,n4092 ,n5710);
    nand g3571(n4514 ,n4001 ,n4151);
    nand g3572(n4865 ,n4143 ,n4632);
    or g3573(n3006 ,n2387 ,n2382);
    or g3574(n5819 ,n5543 ,n5706);
    nand g3575(n2501 ,n0[123] ,n2016);
    nor g3576(n6707 ,n6826 ,n6592);
    xor g3577(n7105 ,n0[45] ,n0[13]);
    nand g3578(n3886 ,n710 ,n3525);
    xnor g3579(n2824 ,n0[117] ,n1339);
    nand g3580(n2551 ,n1136 ,n1898);
    nor g3581(n3346 ,n1954 ,n2900);
    nor g3582(n3449 ,n1954 ,n2888);
    nor g3583(n5415 ,n713 ,n5373);
    or g3584(n2520 ,n6 ,n1977);
    nand g3585(n568 ,n483 ,n567);
    not g3586(n707 ,n721);
    xnor g3587(n2661 ,n1[108] ,n1499);
    nor g3588(n4377 ,n709 ,n4366);
    not g3589(n5264 ,n5263);
    xnor g3590(n6938 ,n232 ,n307);
    xnor g3591(n4918 ,n2812 ,n4442);
    nor g3592(n5322 ,n4750 ,n5085);
    nand g3593(n3483 ,n798 ,n2798);
    nand g3594(n606 ,n475 ,n605);
    nand g3595(n3371 ,n1953 ,n2909);
    xnor g3596(n1691 ,n6898 ,n6899);
    nor g3597(n3671 ,n823 ,n3081);
    nand g3598(n7016 ,n6611 ,n7157);
    or g3599(n2151 ,n1959 ,n1441);
    xnor g3600(n2687 ,n0[125] ,n1259);
    nand g3601(n5481 ,n4705 ,n5299);
    nand g3602(n527 ,n0[107] ,n6964);
    nor g3603(n6723 ,n6826 ,n6599);
    nand g3604(n370 ,n7027 ,n6995);
    xnor g3605(n6896 ,n557 ,n591);
    xnor g3606(n1517 ,n0[82] ,n4[26]);
    xnor g3607(n233 ,n1[60] ,n0[60]);
    nand g3608(n5525 ,n4490 ,n5352);
    nand g3609(n6327 ,n1955 ,n6310);
    not g3610(n4428 ,n4427);
    nor g3611(n4424 ,n2504 ,n4231);
    not g3612(n3264 ,n3236);
    nor g3613(n2335 ,n0[35] ,n1958);
    nor g3614(n6022 ,n4286 ,n5879);
    nand g3615(n4315 ,n3556 ,n3870);
    nor g3616(n2641 ,n0[6] ,n721);
    nand g3617(n466 ,n329 ,n465);
    nand g3618(n4698 ,n717 ,n4431);
    nand g3619(n1104 ,n0[78] ,n792);
    nand g3620(n2474 ,n1997 ,n2030);
    nor g3621(n4231 ,n793 ,n3814);
    nor g3622(n5861 ,n712 ,n5843);
    nor g3623(n2001 ,n863 ,n958);
    nand g3624(n3705 ,n2467 ,n3123);
    xnor g3625(n2813 ,n1262 ,n7116);
    xnor g3626(n1364 ,n0[104] ,n4[0]);
    nor g3627(n5032 ,n3480 ,n4890);
    nor g3628(n2301 ,n1957 ,n1590);
    nor g3629(n5791 ,n5662 ,n5563);
    nand g3630(n2543 ,n1147 ,n1796);
    xnor g3631(n1333 ,n0[119] ,n4[7]);
    nand g3632(n6139 ,n717 ,n6105);
    xnor g3633(n379 ,n7008 ,n7040);
    nor g3634(n3324 ,n1954 ,n2918);
    nand g3635(n4081 ,n720 ,n3699);
    nand g3636(n5131 ,n1039 ,n5014);
    xnor g3637(n3921 ,n1[82] ,n2712);
    xnor g3638(n1594 ,n0[125] ,n1[125]);
    nor g3639(n6056 ,n5631 ,n5976);
    xnor g3640(n2658 ,n1486 ,n1363);
    nand g3641(n6565 ,n6546 ,n6541);
    xnor g3642(n1525 ,n0[9] ,n1[9]);
    nand g3643(n2556 ,n1125 ,n1804);
    or g3644(n3274 ,n2758 ,n3207);
    xnor g3645(n2933 ,n1619 ,n1518);
    nand g3646(n2534 ,n1223 ,n1908);
    not g3647(n792 ,n6);
    nand g3648(n3936 ,n2182 ,n3635);
    nor g3649(n5123 ,n4055 ,n4973);
    nor g3650(n5772 ,n794 ,n5639);
    xnor g3651(n6952 ,n540 ,n619);
    xnor g3652(n6908 ,n529 ,n597);
    nor g3653(n5916 ,n5560 ,n5796);
    nand g3654(n2585 ,n1075 ,n1857);
    or g3655(n6091 ,n6003 ,n5783);
    not g3656(n826 ,n0[39]);
    xnor g3657(n6880 ,n553 ,n583);
    nand g3658(n5921 ,n5426 ,n5798);
    nor g3659(n6433 ,n3431 ,n6342);
    nor g3660(n2081 ,n1958 ,n1639);
    nand g3661(n5119 ,n798 ,n4908);
    nand g3662(n6403 ,n3433 ,n6342);
    or g3663(n2253 ,n709 ,n1456);
    nor g3664(n5270 ,n4195 ,n5062);
    not g3665(n839 ,n1[32]);
    or g3666(n2731 ,n944 ,n2576);
    nor g3667(n6103 ,n4291 ,n6005);
    or g3668(n3805 ,n6825 ,n2845);
    not g3669(n770 ,n1[47]);
    not g3670(n6243 ,n6242);
    xnor g3671(n1524 ,n0[58] ,n4[18]);
    nor g3672(n4292 ,n824 ,n4016);
    or g3673(n9[61] ,n5911 ,n5967);
    not g3674(n1225 ,n1224);
    nand g3675(n5716 ,n4002 ,n5403);
    or g3676(n4629 ,n3509 ,n4549);
    nor g3677(n4317 ,n780 ,n3914);
    nand g3678(n5769 ,n4388 ,n5643);
    not g3679(n1568 ,n1567);
    nor g3680(n4164 ,n789 ,n4112);
    nor g3681(n6153 ,n5814 ,n6079);
    nand g3682(n277 ,n223 ,n276);
    nor g3683(n3620 ,n771 ,n2794);
    nor g3684(n2096 ,n1956 ,n1521);
    nand g3685(n5857 ,n1955 ,n5769);
    nor g3686(n6231 ,n5468 ,n6168);
    xnor g3687(n557 ,n6970 ,n0[113]);
    nand g3688(n4578 ,n2518 ,n4215);
    nor g3689(n6718 ,n6826 ,n6594);
    nand g3690(n655 ,n1[7] ,n621);
    nand g3691(n268 ,n187 ,n267);
    not g3692(n6197 ,n6196);
    xor g3693(n7122 ,n0[62] ,n0[30]);
    nor g3694(n6321 ,n711 ,n6309);
    or g3695(n320 ,n7038 ,n7006);
    nand g3696(n1005 ,n0[32] ,n747);
    xnor g3697(n5576 ,n1346 ,n5202);
    nand g3698(n4276 ,n0[68] ,n3903);
    nand g3699(n3759 ,n7161 ,n3056);
    nor g3700(n718 ,n3[1] ,n1148);
    nor g3701(n6600 ,n0[123] ,n0[91]);
    nand g3702(n2481 ,n0[64] ,n1764);
    nor g3703(n3413 ,n1954 ,n2862);
    nor g3704(n1741 ,n977 ,n1056);
    or g3705(n4216 ,n792 ,n3819);
    not g3706(n5086 ,n5085);
    nand g3707(n1130 ,n6896 ,n797);
    xnor g3708(n3931 ,n2964 ,n1976);
    xnor g3709(n5586 ,n4988 ,n5208);
    nand g3710(n6151 ,n3327 ,n6036);
    xnor g3711(n2695 ,n4[19] ,n1521);
    nand g3712(n6181 ,n3268 ,n6137);
    nand g3713(n1060 ,n0[29] ,n709);
    nand g3714(n3561 ,n787 ,n3257);
    xnor g3715(n1326 ,n0[32] ,n1[48]);
    or g3716(n3025 ,n2287 ,n2286);
    xnor g3717(n1320 ,n0[78] ,n7106);
    xor g3718(n7050 ,n0[96] ,n0[64]);
    nor g3719(n3796 ,n1222 ,n2801);
    nor g3720(n2112 ,n787 ,n1462);
    not g3721(n772 ,n1[45]);
    nand g3722(n346 ,n7039 ,n7007);
    nor g3723(n1074 ,n775 ,n710);
    xnor g3724(n5585 ,n4669 ,n5265);
    nand g3725(n584 ,n479 ,n583);
    not g3726(n4888 ,n4887);
    nand g3727(n5700 ,n4523 ,n5418);
    nor g3728(n4373 ,n4294 ,n4284);
    nand g3729(n434 ,n343 ,n433);
    xnor g3730(n391 ,n6989 ,n7021);
    or g3731(n3903 ,n2336 ,n3490);
    nand g3732(n6004 ,n3302 ,n5858);
    nand g3733(n304 ,n176 ,n303);
    nand g3734(n6428 ,n3359 ,n6330);
    xnor g3735(n1435 ,n1[89] ,n2[25]);
    nor g3736(n3498 ,n6825 ,n2821);
    nand g3737(n3215 ,n1137 ,n2145);
    nand g3738(n6629 ,n0[72] ,n6580);
    nand g3739(n3489 ,n2795 ,n2796);
    xnor g3740(n1369 ,n6869 ,n6868);
    nand g3741(n3765 ,n6804 ,n3074);
    nand g3742(n2455 ,n0[8] ,n1773);
    nor g3743(n2735 ,n2047 ,n2110);
    xnor g3744(n1402 ,n1[32] ,n2[32]);
    nor g3745(n3354 ,n1954 ,n2903);
    not g3746(n5278 ,n5277);
    xnor g3747(n2897 ,n1326 ,n1511);
    nand g3748(n5675 ,n4189 ,n5521);
    nand g3749(n7005 ,n6625 ,n7168);
    nand g3750(n1032 ,n0[1] ,n804);
    or g3751(n178 ,n0[54] ,n1[54]);
    nor g3752(n1779 ,n0[37] ,n965);
    xnor g3753(n2645 ,n1991 ,n2004);
    nor g3754(n2788 ,n2038 ,n2123);
    nor g3755(n2090 ,n6 ,n1976);
    xnor g3756(n6341 ,n6188 ,n6141);
    nor g3757(n3071 ,n1837 ,n2039);
    nor g3758(n2408 ,n0[52] ,n1957);
    or g3759(n3545 ,n1954 ,n2960);
    nand g3760(n6674 ,n1[64] ,n6580);
    nand g3761(n6785 ,n1[106] ,n7088);
    or g3762(n4149 ,n6 ,n4098);
    nor g3763(n1826 ,n744 ,n11);
    or g3764(n2298 ,n1961 ,n1886);
    xnor g3765(n2819 ,n1369 ,n1677);
    nand g3766(n7132 ,n6663 ,n6720);
    or g3767(n2780 ,n2127 ,n2126);
    nor g3768(n6737 ,n3[0] ,n6736);
    xnor g3769(n5727 ,n4662 ,n5456);
    nand g3770(n4781 ,n1794 ,n4517);
    nand g3771(n3779 ,n1129 ,n3164);
    nand g3772(n3183 ,n1973 ,n2326);
    nor g3773(n4376 ,n788 ,n4366);
    or g3774(n4206 ,n4049 ,n3777);
    nand g3775(n2610 ,n884 ,n1809);
    nand g3776(n375 ,n7029 ,n6997);
    nor g3777(n6437 ,n3719 ,n6324);
    not g3778(n835 ,n0[93]);
    nand g3779(n52 ,n7079 ,n0[23]);
    nand g3780(n6275 ,n6233 ,n6217);
    nor g3781(n991 ,n725 ,n0[43]);
    nor g3782(n3114 ,n2452 ,n2247);
    xnor g3783(n1249 ,n0[94] ,n7122);
    nand g3784(n4113 ,n2455 ,n3439);
    or g3785(n4394 ,n2790 ,n4336);
    not g3786(n5070 ,n5069);
    nand g3787(n643 ,n0[80] ,n622);
    nand g3788(n6995 ,n6647 ,n6813);
    nor g3789(n4509 ,n4295 ,n4317);
    nor g3790(n2185 ,n1956 ,n1630);
    nor g3791(n4183 ,n715 ,n4110);
    nand g3792(n684 ,n1[6] ,n621);
    xnor g3793(n3836 ,n2706 ,n2649);
    nand g3794(n441 ,n352 ,n440);
    nor g3795(n5621 ,n5084 ,n5394);
    nand g3796(n3555 ,n1953 ,n2880);
    nand g3797(n6270 ,n6186 ,n6204);
    xor g3798(n701 ,n5838 ,n6195);
    nand g3799(n6616 ,n0[111] ,n0[79]);
    xnor g3800(n6337 ,n6249 ,n5931);
    xnor g3801(n1301 ,n1[41] ,n4[1]);
    nand g3802(n950 ,n0[22] ,n791);
    nor g3803(n5597 ,n4695 ,n5455);
    nand g3804(n6978 ,n6750 ,n6778);
    nand g3805(n3351 ,n1952 ,n2895);
    nand g3806(n1089 ,n0[63] ,n791);
    xnor g3807(n6385 ,n6306 ,n6308);
    nor g3808(n3919 ,n2466 ,n3765);
    xnor g3809(n6884 ,n554 ,n585);
    nand g3810(n3347 ,n1952 ,n2856);
    xnor g3811(n1576 ,n1[43] ,n1[11]);
    nor g3812(n6361 ,n1954 ,n6250);
    nor g3813(n2144 ,n899 ,n1961);
    nand g3814(n3280 ,n852 ,n3096);
    nor g3815(n3330 ,n2374 ,n3127);
    nand g3816(n1103 ,n0[21] ,n708);
    nand g3817(n274 ,n186 ,n273);
    nand g3818(n2533 ,n793 ,n1968);
    or g3819(n5611 ,n5535 ,n5216);
    nand g3820(n6102 ,n3996 ,n5966);
    nor g3821(n2444 ,n0[66] ,n1992);
    nand g3822(n3486 ,n1953 ,n2952);
    nor g3823(n6038 ,n711 ,n5974);
    xnor g3824(n556 ,n6969 ,n0[112]);
    nand g3825(n3075 ,n1220 ,n2351);
    xnor g3826(n398 ,n6996 ,n7028);
    nand g3827(n2205 ,n1790 ,n2022);
    or g3828(n4630 ,n3498 ,n4557);
    nor g3829(n2338 ,n0[34] ,n1957);
    nor g3830(n1823 ,n736 ,n1220);
    nor g3831(n1097 ,n807 ,n731);
    nor g3832(n4005 ,n833 ,n3279);
    nand g3833(n1198 ,n6843 ,n796);
    xnor g3834(n1518 ,n0[59] ,n4[19]);
    nor g3835(n2991 ,n1741 ,n2501);
    nand g3836(n2496 ,n0[63] ,n718);
    nand g3837(n6468 ,n6451 ,n6429);
    nor g3838(n2437 ,n1961 ,n1413);
    nand g3839(n3410 ,n3122 ,n3120);
    xnor g3840(n1373 ,n0[83] ,n7111);
    nor g3841(n2739 ,n725 ,n2462);
    xnor g3842(n2825 ,n1272 ,n1659);
    nand g3843(n1153 ,n6848 ,n795);
    nor g3844(n5314 ,n3427 ,n5181);
    nor g3845(n1754 ,n724 ,n1006);
    or g3846(n4172 ,n2154 ,n3876);
    not g3847(n827 ,n0[45]);
    nand g3848(n995 ,n0[48] ,n714);
    xnor g3849(n5019 ,n4596 ,n4099);
    nor g3850(n3055 ,n1803 ,n2486);
    nor g3851(n2733 ,n725 ,n2043);
    nand g3852(n609 ,n523 ,n608);
    nand g3853(n5326 ,n790 ,n5082);
    nor g3854(n2741 ,n2061 ,n2051);
    nand g3855(n5801 ,n4044 ,n5703);
    or g3856(n2238 ,n1962 ,n1427);
    nand g3857(n5833 ,n4494 ,n5643);
    nand g3858(n6812 ,n6581 ,n7102);
    nand g3859(n156 ,n17 ,n155);
    nor g3860(n4419 ,n4166 ,n4320);
    xnor g3861(n2675 ,n1660 ,n1608);
    nand g3862(n579 ,n526 ,n578);
    nand g3863(n3190 ,n740 ,n2530);
    nand g3864(n890 ,n0[106] ,n724);
    xnor g3865(n6907 ,n103 ,n139);
    nand g3866(n9[96] ,n5258 ,n6528);
    nand g3867(n424 ,n335 ,n423);
    nand g3868(n5425 ,n5102 ,n5276);
    nand g3869(n607 ,n510 ,n606);
    nor g3870(n1772 ,n725 ,n900);
    nand g3871(n3594 ,n0[56] ,n2989);
    xor g3872(n4912 ,n4435 ,n2828);
    nand g3873(n5557 ,n4825 ,n5235);
    nor g3874(n2348 ,n0[46] ,n1956);
    xnor g3875(n2871 ,n1604 ,n1522);
    nand g3876(n514 ,n0[100] ,n6957);
    nand g3877(n106 ,n28 ,n105);
    nand g3878(n4335 ,n2579 ,n3922);
    or g3879(n2064 ,n1959 ,n1476);
    nand g3880(n3635 ,n1[51] ,n2979);
    nor g3881(n5352 ,n5187 ,n5048);
    nand g3882(n7036 ,n6650 ,n7137);
    xnor g3883(n6859 ,n91 ,n115);
    nand g3884(n4007 ,n0[102] ,n3490);
    nor g3885(n3509 ,n6825 ,n2809);
    nor g3886(n3627 ,n3241 ,n3023);
    xnor g3887(n5197 ,n4997 ,n1489);
    nor g3888(n3062 ,n1824 ,n2280);
    or g3889(n2190 ,n1960 ,n1940);
    nand g3890(n3084 ,n1220 ,n2397);
    nand g3891(n5473 ,n4701 ,n5333);
    xnor g3892(n1570 ,n0[116] ,n0[100]);
    nor g3893(n2356 ,n721 ,n1577);
    xnor g3894(n1352 ,n0[88] ,n4[16]);
    nand g3895(n2448 ,n0[35] ,n718);
    xnor g3896(n4213 ,n3539 ,n1988);
    or g3897(n3027 ,n2191 ,n2292);
    nor g3898(n6155 ,n3388 ,n6038);
    nand g3899(n9[82] ,n5688 ,n6167);
    nor g3900(n4663 ,n946 ,n4471);
    nand g3901(n1110 ,n6840 ,n795);
    nand g3902(n4817 ,n1966 ,n4444);
    nor g3903(n1801 ,n730 ,n11);
    nand g3904(n10[1] ,n4744 ,n4863);
    nand g3905(n5501 ,n4685 ,n5351);
    nor g3906(n3894 ,n3383 ,n3382);
    nor g3907(n5461 ,n4162 ,n5272);
    nor g3908(n2996 ,n1567 ,n2631);
    nand g3909(n2498 ,n1907 ,n1782);
    nand g3910(n4131 ,n708 ,n3963);
    nor g3911(n3418 ,n788 ,n3254);
    not g3912(n1551 ,n1550);
    nand g3913(n2602 ,n0[15] ,n1964);
    nor g3914(n6374 ,n3457 ,n6261);
    or g3915(n9[104] ,n5303 ,n6532);
    nand g3916(n2492 ,n0[51] ,n718);
    xnor g3917(n4212 ,n3540 ,n2003);
    or g3918(n9[43] ,n4498 ,n6568);
    nor g3919(n3367 ,n1[92] ,n2961);
    or g3920(n4058 ,n3655 ,n3516);
    or g3921(n3014 ,n2638 ,n2368);
    nor g3922(n2367 ,n0[50] ,n1956);
    nand g3923(n5540 ,n4706 ,n5314);
    not g3924(n5460 ,n5459);
    nor g3925(n5194 ,n6824 ,n4917);
    nand g3926(n5212 ,n4980 ,n5075);
    nand g3927(n5463 ,n4406 ,n5273);
    nand g3928(n6516 ,n6466 ,n6465);
    nand g3929(n6541 ,n717 ,n6512);
    nor g3930(n1745 ,n788 ,n911);
    nor g3931(n3153 ,n837 ,n2344);
    nand g3932(n462 ,n322 ,n461);
    xnor g3933(n4476 ,n3941 ,n2816);
    nand g3934(n4572 ,n1084 ,n4224);
    xnor g3935(n5293 ,n4211 ,n4994);
    nand g3936(n5609 ,n5547 ,n5412);
    or g3937(n3864 ,n787 ,n3795);
    xnor g3938(n544 ,n6957 ,n0[100]);
    nand g3939(n4483 ,n3616 ,n4180);
    or g3940(n5060 ,n2460 ,n4884);
    nand g3941(n6383 ,n6284 ,n6287);
    nand g3942(n4646 ,n4032 ,n4534);
    not g3943(n4232 ,n4231);
    nand g3944(n2005 ,n0[56] ,n992);
    nand g3945(n6990 ,n6615 ,n6818);
    xnor g3946(n5722 ,n5007 ,n5530);
    nand g3947(n6429 ,n6085 ,n6337);
    xnor g3948(n3952 ,n2826 ,n2811);
    nand g3949(n61 ,n7063 ,n0[7]);
    not g3950(n815 ,n0[111]);
    xnor g3951(n1925 ,n1[43] ,n2[43]);
    xnor g3952(n542 ,n6955 ,n0[98]);
    nand g3953(n4769 ,n2560 ,n4434);
    xor g3954(n2914 ,n1[96] ,n1569);
    nand g3955(n5164 ,n798 ,n4920);
    nand g3956(n2536 ,n1146 ,n1851);
    or g3957(n2757 ,n2425 ,n2076);
    or g3958(n722 ,n3[0] ,n1950);
    nand g3959(n4575 ,n2520 ,n4230);
    nand g3960(n4770 ,n2560 ,n4435);
    nor g3961(n5116 ,n6 ,n5006);
    nor g3962(n6373 ,n3342 ,n6259);
    nand g3963(n5420 ,n4981 ,n5279);
    not g3964(n3962 ,n3961);
    or g3965(n2245 ,n719 ,n1622);
    nand g3966(n6619 ,n1[71] ,n6580);
    nand g3967(n2230 ,n793 ,n2001);
    nand g3968(n2114 ,n794 ,n1999);
    nand g3969(n6653 ,n1[83] ,n6579);
    or g3970(n15 ,n7074 ,n0[18]);
    nor g3971(n4775 ,n727 ,n689);
    xnor g3972(n2810 ,n1305 ,n1682);
    nor g3973(n2354 ,n0[57] ,n1957);
    nor g3974(n5623 ,n5100 ,n5459);
    or g3975(n3359 ,n1954 ,n2878);
    xor g3976(n7092 ,n0[32] ,n0[0]);
    not g3977(n5482 ,n5481);
    nand g3978(n3690 ,n787 ,n3261);
    nand g3979(n1126 ,n1[64] ,n2[0]);
    nor g3980(n2305 ,n1961 ,n1421);
    nor g3981(n2415 ,n0[119] ,n1957);
    or g3982(n4053 ,n3649 ,n3533);
    not g3983(n759 ,n0[115]);
    nor g3984(n2328 ,n725 ,n1844);
    xnor g3985(n2831 ,n0[101] ,n1283);
    nand g3986(n208 ,n0[48] ,n1[48]);
    or g3987(n5328 ,n3532 ,n5040);
    nand g3988(n5509 ,n794 ,n5379);
    xnor g3989(n1702 ,n0[68] ,n1[84]);
    nand g3990(n3883 ,n709 ,n3523);
    nor g3991(n1755 ,n859 ,n1027);
    xnor g3992(n2823 ,n0[105] ,n1288);
    nor g3993(n2358 ,n721 ,n1534);
    or g3994(n9[124] ,n5618 ,n5926);
    xnor g3995(n6511 ,n6188 ,n6413);
    nand g3996(n4640 ,n717 ,n4467);
    nor g3997(n3707 ,n1[54] ,n3176);
    nand g3998(n2007 ,n1228 ,n1012);
    nor g3999(n1850 ,n754 ,n11);
    not g4000(n6730 ,n3[3]);
    nor g4001(n6063 ,n5737 ,n5964);
    or g4002(n2069 ,n719 ,n1490);
    nand g4003(n1197 ,n6924 ,n795);
    not g4004(n805 ,n0[25]);
    nand g4005(n2471 ,n0[38] ,n718);
    nor g4006(n3655 ,n811 ,n3076);
    nand g4007(n1134 ,n6845 ,n795);
    xnor g4008(n6902 ,n254 ,n289);
    nand g4009(n6186 ,n3322 ,n6126);
    nor g4010(n3428 ,n1954 ,n2930);
    nand g4011(n4815 ,n1966 ,n4445);
    xnor g4012(n1597 ,n0[32] ,n1[32]);
    nor g4013(n2309 ,n1956 ,n1922);
    nand g4014(n6762 ,n0[52] ,n6737);
    nor g4015(n4525 ,n4163 ,n4338);
    nand g4016(n3716 ,n2458 ,n3186);
    nor g4017(n6108 ,n4942 ,n5981);
    xnor g4018(n2882 ,n1348 ,n1602);
    xnor g4019(n1340 ,n0[79] ,n4[7]);
    xnor g4020(n1601 ,n0[67] ,n1[67]);
    nand g4021(n7168 ,n6581 ,n7111);
    nand g4022(n948 ,n0[26] ,n725);
    not g4023(n1043 ,n1042);
    nand g4024(n269 ,n213 ,n268);
    xnor g4025(n1430 ,n1[24] ,n2[24]);
    not g4026(n1029 ,n1028);
    not g4027(n4816 ,n4815);
    nor g4028(n2283 ,n6 ,n1971);
    not g4029(n4220 ,n4219);
    or g4030(n9[1] ,n4148 ,n6506);
    nor g4031(n5622 ,n5193 ,n5424);
    nand g4032(n4080 ,n720 ,n3700);
    nand g4033(n1131 ,n6915 ,n796);
    nor g4034(n6446 ,n6088 ,n6344);
    nor g4035(n5928 ,n4322 ,n5787);
    or g4036(n3300 ,n1954 ,n2873);
    nand g4037(n3461 ,n798 ,n2822);
    not g4038(n5972 ,n5971);
    xnor g4039(n1586 ,n0[110] ,n1[110]);
    nor g4040(n5255 ,n4301 ,n5185);
    not g4041(n4210 ,n4209);
    nor g4042(n2624 ,n0[21] ,n1963);
    or g4043(n6123 ,n706 ,n6106);
    xnor g4044(n1403 ,n1[126] ,n2[62]);
    nand g4045(n3112 ,n0[35] ,n2576);
    xnor g4046(n4845 ,n4587 ,n4453);
    nand g4047(n7162 ,n6581 ,n7117);
    nand g4048(n3244 ,n1214 ,n2453);
    nand g4049(n9[97] ,n4974 ,n6390);
    nand g4050(n6621 ,n1[72] ,n6579);
    or g4051(n3854 ,n2254 ,n3756);
    xnor g4052(n1933 ,n1[94] ,n2[30]);
    nand g4053(n7029 ,n6631 ,n7144);
    nor g4054(n4214 ,n3586 ,n3852);
    nand g4055(n3173 ,n1980 ,n2326);
    nand g4056(n5767 ,n5566 ,n5697);
    nand g4057(n3270 ,n1952 ,n2923);
    nor g4058(n2628 ,n0[18] ,n721);
    nand g4059(n6655 ,n0[116] ,n0[84]);
    nand g4060(n937 ,n0[17] ,n818);
    nand g4061(n3238 ,n1208 ,n2153);
    nand g4062(n7140 ,n6616 ,n6712);
    nand g4063(n3677 ,n0[4] ,n3078);
    nor g4064(n4794 ,n3642 ,n4566);
    nand g4065(n4638 ,n2791 ,n4386);
    or g4066(n2975 ,n2324 ,n2173);
    nand g4067(n6994 ,n6629 ,n6814);
    xor g4068(n7053 ,n0[99] ,n0[67]);
    xnor g4069(n4451 ,n3945 ,n2824);
    nand g4070(n6525 ,n6464 ,n6467);
    not g4071(n830 ,n1[63]);
    nand g4072(n4360 ,n3890 ,n4051);
    or g4073(n3897 ,n2212 ,n3743);
    xnor g4074(n2887 ,n1275 ,n1656);
    xnor g4075(n2877 ,n1487 ,n1711);
    or g4076(n4849 ,n2325 ,n4677);
    nand g4077(n135 ,n56 ,n134);
    nor g4078(n4688 ,n706 ,n4426);
    nor g4079(n5135 ,n727 ,n4897);
    nor g4080(n5323 ,n4629 ,n5090);
    nor g4081(n5311 ,n3419 ,n5077);
    nand g4082(n4092 ,n7142 ,n3460);
    nand g4083(n4346 ,n3602 ,n3982);
    nand g4084(n5027 ,n710 ,n5013);
    nor g4085(n4020 ,n3203 ,n3404);
    or g4086(n4706 ,n1965 ,n4466);
    nor g4087(n6310 ,n5650 ,n6194);
    nor g4088(n6545 ,n5159 ,n6519);
    nor g4089(n3460 ,n2293 ,n3027);
    xnor g4090(n1664 ,n6883 ,n6880);
    nand g4091(n3250 ,n894 ,n2032);
    xnor g4092(n4443 ,n2805 ,n3960);
    xnor g4093(n1616 ,n0[120] ,n1[120]);
    xnor g4094(n1599 ,n0[64] ,n1[64]);
    nand g4095(n6646 ,n0[113] ,n0[81]);
    nand g4096(n4487 ,n3410 ,n4310);
    nand g4097(n894 ,n0[2] ,n725);
    nand g4098(n6631 ,n1[75] ,n6579);
    xnor g4099(n5458 ,n4580 ,n5155);
    xnor g4100(n1329 ,n6946 ,n6947);
    nor g4101(n3341 ,n1954 ,n2895);
    nand g4102(n2493 ,n0[55] ,n718);
    nand g4103(n3606 ,n0[77] ,n2796);
    nand g4104(n4205 ,n3738 ,n3869);
    not g4105(n736 ,n0[120]);
    nand g4106(n3145 ,n2587 ,n2448);
    xnor g4107(n2706 ,n0[79] ,n1979);
    nor g4108(n5338 ,n4623 ,n5166);
    nand g4109(n2552 ,n1122 ,n1895);
    not g4110(n2796 ,n2797);
    nand g4111(n142 ,n16 ,n141);
    or g4112(n187 ,n0[39] ,n1[39]);
    nand g4113(n9[39] ,n5666 ,n5742);
    or g4114(n3519 ,n2984 ,n2730);
    nand g4115(n6090 ,n3345 ,n5955);
    not g4116(n725 ,n7);
    nand g4117(n7044 ,n6673 ,n7129);
    xnor g4118(n76 ,n0[23] ,n7079);
    xnor g4119(n1501 ,n0[86] ,n4[30]);
    nand g4120(n6531 ,n6478 ,n6492);
    nor g4121(n6477 ,n6370 ,n6419);
    nand g4122(n2011 ,n0[17] ,n1046);
    not g4123(n989 ,n988);
    xnor g4124(n1655 ,n6874 ,n6875);
    nand g4125(n447 ,n369 ,n446);
    nand g4126(n294 ,n168 ,n293);
    nand g4127(n3847 ,n723 ,n3802);
    or g4128(n4025 ,n3213 ,n3385);
    xnor g4129(n5274 ,n4669 ,n5000);
    nand g4130(n442 ,n319 ,n441);
    nand g4131(n1920 ,n1230 ,n918);
    not g4132(n5565 ,n5564);
    nand g4133(n3138 ,n1[37] ,n2378);
    or g4134(n2115 ,n719 ,n1588);
    nor g4135(n954 ,n1[117] ,n2[53]);
    xnor g4136(n5228 ,n4872 ,n4212);
    nand g4137(n2262 ,n792 ,n1987);
    xnor g4138(n2816 ,n1383 ,n1721);
    nand g4139(n3972 ,n0[7] ,n3490);
    nand g4140(n372 ,n7044 ,n7012);
    nand g4141(n151 ,n54 ,n150);
    xnor g4142(n6279 ,n6114 ,n2704);
    nand g4143(n6657 ,n0[85] ,n6579);
    xnor g4144(n103 ,n0[19] ,n7075);
    nor g4145(n6475 ,n5388 ,n6389);
    nor g4146(n2463 ,n1961 ,n1391);
    not g4147(n5373 ,n5374);
    nor g4148(n3499 ,n6825 ,n2810);
    nand g4149(n3996 ,n0[100] ,n3490);
    nand g4150(n897 ,n0[82] ,n724);
    nor g4151(n4495 ,n2559 ,n4174);
    nor g4152(n5362 ,n3518 ,n5143);
    nand g4153(n6779 ,n1[111] ,n7088);
    nand g4154(n686 ,n1[31] ,n621);
    nand g4155(n3699 ,n1[93] ,n2959);
    nand g4156(n7001 ,n6688 ,n6807);
    or g4157(n6003 ,n3485 ,n5895);
    nor g4158(n4744 ,n3536 ,n4564);
    not g4159(n6731 ,n3[2]);
    nand g4160(n6695 ,n0[65] ,n6580);
    nand g4161(n6453 ,n3407 ,n6335);
    nand g4162(n367 ,n7026 ,n6994);
    nand g4163(n920 ,n0[65] ,n814);
    nor g4164(n6508 ,n6446 ,n6436);
    xnor g4165(n1647 ,n0[91] ,n4[19]);
    nor g4166(n2217 ,n719 ,n1537);
    nor g4167(n3965 ,n2329 ,n3590);
    nand g4168(n6376 ,n6298 ,n6302);
    nand g4169(n918 ,n813 ,n754);
    nand g4170(n3701 ,n1[64] ,n2914);
    nand g4171(n4949 ,n3393 ,n4736);
    nand g4172(n6735 ,n3[2] ,n6732);
    nor g4173(n2082 ,n1961 ,n1448);
    nor g4174(n3041 ,n1553 ,n2640);
    nand g4175(n2019 ,n723 ,n1019);
    or g4176(n4399 ,n3785 ,n4270);
    or g4177(n5404 ,n5103 ,n5260);
    nand g4178(n4767 ,n2560 ,n4445);
    xnor g4179(n2701 ,n1[120] ,n1554);
    nor g4180(n5981 ,n793 ,n5853);
    nand g4181(n960 ,n6825 ,n727);
    nand g4182(n3313 ,n1952 ,n2859);
    nor g4183(n1878 ,n767 ,n11);
    xnor g4184(n2809 ,n1266 ,n1688);
    xnor g4185(n4371 ,n3246 ,n3961);
    or g4186(n6498 ,n5993 ,n6457);
    nand g4187(n258 ,n180 ,n257);
    xnor g4188(n6950 ,n235 ,n313);
    nand g4189(n4404 ,n875 ,n4268);
    not g4190(n6803 ,n7159);
    nand g4191(n2547 ,n1182 ,n1822);
    xnor g4192(n1533 ,n1[49] ,n1[17]);
    xnor g4193(n382 ,n7011 ,n7043);
    nor g4194(n926 ,n0[95] ,n789);
    nand g4195(n5927 ,n5524 ,n5786);
    xnor g4196(n1259 ,n0[93] ,n7121);
    not g4197(n5294 ,n5293);
    nand g4198(n5668 ,n4402 ,n5484);
    nand g4199(n3622 ,n1[45] ,n2795);
    nor g4200(n3374 ,n1954 ,n2912);
    nand g4201(n2558 ,n1140 ,n1859);
    nor g4202(n1877 ,n766 ,n11);
    xnor g4203(n1573 ,n0[50] ,n4[10]);
    nor g4204(n1828 ,n806 ,n11);
    nand g4205(n7155 ,n6581 ,n7050);
    xnor g4206(n1620 ,n0[72] ,n1[72]);
    or g4207(n26 ,n7078 ,n0[22]);
    nor g4208(n6540 ,n5561 ,n6536);
    xnor g4209(n6887 ,n98 ,n129);
    nand g4210(n313 ,n195 ,n312);
    nand g4211(n6997 ,n6659 ,n6811);
    nand g4212(n439 ,n360 ,n438);
    nor g4213(n2584 ,n749 ,n721);
    nand g4214(n65 ,n7076 ,n0[20]);
    nor g4215(n2059 ,n1961 ,n1917);
    nor g4216(n5758 ,n713 ,n5584);
    nor g4217(n3878 ,n2373 ,n3490);
    nand g4218(n3772 ,n1186 ,n2751);
    xnor g4219(n5263 ,n4997 ,n5004);
    nand g4220(n3192 ,n1967 ,n2326);
    nor g4221(n5149 ,n727 ,n4922);
    or g4222(n4714 ,n3524 ,n4558);
    nand g4223(n1035 ,n0[113] ,n738);
    nor g4224(n3365 ,n1954 ,n2907);
    nand g4225(n4161 ,n792 ,n3961);
    nand g4226(n650 ,n0[68] ,n622);
    xnor g4227(n1548 ,n0[26] ,n1[26]);
    nand g4228(n3706 ,n2102 ,n3173);
    nor g4229(n3668 ,n2484 ,n3036);
    xnor g4230(n1929 ,n1[101] ,n2[37]);
    xnor g4231(n4844 ,n4359 ,n4441);
    nor g4232(n2067 ,n1961 ,n1437);
    nand g4233(n4319 ,n2326 ,n4102);
    xnor g4234(n3849 ,n1[88] ,n2701);
    or g4235(n2983 ,n2624 ,n2413);
    nand g4236(n3179 ,n1983 ,n2326);
    nand g4237(n10[24] ,n4619 ,n5321);
    xnor g4238(n6215 ,n6106 ,n5972);
    nor g4239(n2290 ,n721 ,n1542);
    xnor g4240(n5583 ,n4670 ,n5260);
    nor g4241(n2164 ,n1961 ,n1386);
    nor g4242(n1052 ,n709 ,n0[6]);
    not g4243(n6825 ,n6734);
    or g4244(n7088 ,n6734 ,n6827);
    nand g4245(n3443 ,n1952 ,n2955);
    nor g4246(n4136 ,n1959 ,n3817);
    nand g4247(n9[62] ,n4277 ,n5635);
    nand g4248(n4734 ,n6827 ,n4473);
    nand g4249(n3764 ,n7157 ,n3073);
    nor g4250(n2180 ,n1959 ,n1943);
    nand g4251(n443 ,n363 ,n442);
    or g4252(n337 ,n7026 ,n6994);
    not g4253(n5891 ,n5890);
    nand g4254(n4425 ,n2308 ,n4230);
    nand g4255(n4526 ,n2005 ,n4367);
    xnor g4256(n1394 ,n1[49] ,n2[49]);
    xnor g4257(n1625 ,n0[102] ,n1[102]);
    nand g4258(n270 ,n185 ,n269);
    nand g4259(n2505 ,n1846 ,n1868);
    nor g4260(n1762 ,n1038 ,n853);
    xnor g4261(n555 ,n6968 ,n0[111]);
    nand g4262(n3080 ,n11 ,n2379);
    nand g4263(n5408 ,n5248 ,n5251);
    not g4264(n620 ,n7088);
    nand g4265(n2020 ,n714 ,n1038);
    xnor g4266(n1429 ,n0[45] ,n0[37]);
    nand g4267(n6058 ,n6018 ,n5782);
    nor g4268(n1837 ,n812 ,n11);
    nand g4269(n3630 ,n0[62] ,n2794);
    nand g4270(n6133 ,n700 ,n6058);
    nor g4271(n2486 ,n721 ,n1500);
    xnor g4272(n1629 ,n0[94] ,n1[94]);
    nor g4273(n3562 ,n710 ,n3254);
    xnor g4274(n6281 ,n5932 ,n6173);
    not g4275(n2886 ,n2885);
    xnor g4276(n6072 ,n5639 ,n5935);
    nand g4277(n3950 ,n3444 ,n3558);
    nand g4278(n6267 ,n717 ,n6244);
    nand g4279(n6476 ,n6445 ,n6427);
    nor g4280(n4871 ,n3364 ,n4600);
    or g4281(n5952 ,n712 ,n5940);
    nand g4282(n3643 ,n0[53] ,n2796);
    or g4283(n4197 ,n2325 ,n3957);
    nor g4284(n4221 ,n3418 ,n3984);
    xnor g4285(n1578 ,n0[20] ,n1[20]);
    xnor g4286(n5584 ,n5264 ,n4211);
    nand g4287(n6296 ,n4252 ,n6231);
    not g4288(n760 ,n0[91]);
    or g4289(n4027 ,n3214 ,n3380);
    nand g4290(n2530 ,n977 ,n1903);
    nand g4291(n9[120] ,n5669 ,n6538);
    nor g4292(n5309 ,n3412 ,n5178);
    not g4293(n773 ,n0[28]);
    nor g4294(n2049 ,n0[73] ,n1733);
    xnor g4295(n2932 ,n1635 ,n1580);
    nand g4296(n6742 ,n0[55] ,n6737);
    nand g4297(n6352 ,n6265 ,n6282);
    nor g4298(n4176 ,n3221 ,n4067);
    nor g4299(n4534 ,n3497 ,n4250);
    xor g4300(n7101 ,n0[41] ,n0[9]);
    nand g4301(n1127 ,n6907 ,n795);
    nand g4302(n1191 ,n6897 ,n795);
    nor g4303(n3137 ,n1845 ,n2588);
    xnor g4304(n1623 ,n0[112] ,n1[112]);
    xnor g4305(n1611 ,n0[65] ,n1[65]);
    xnor g4306(n2807 ,n1378 ,n1691);
    nand g4307(n6643 ,n0[88] ,n6580);
    xnor g4308(n3820 ,n1[65] ,n2710);
    not g4309(n5888 ,n5887);
    nand g4310(n1155 ,n6875 ,n796);
    nand g4311(n1044 ,n821 ,n769);
    nor g4312(n3658 ,n737 ,n3089);
    or g4313(n183 ,n0[41] ,n1[41]);
    nor g4314(n5368 ,n3808 ,n5150);
    nand g4315(n5380 ,n4170 ,n5128);
    or g4316(n3030 ,n2300 ,n2296);
    nand g4317(n122 ,n34 ,n121);
    nor g4318(n4225 ,n2781 ,n3865);
    or g4319(n3896 ,n2122 ,n3711);
    not g4320(n2560 ,n2561);
    nand g4321(n273 ,n218 ,n272);
    nand g4322(n6367 ,n6285 ,n6288);
    nor g4323(n3337 ,n1222 ,n2821);
    nand g4324(n3721 ,n3180 ,n2788);
    nor g4325(n4023 ,n3209 ,n3392);
    nand g4326(n1848 ,n0[68] ,n964);
    xnor g4327(n6890 ,n251 ,n283);
    nor g4328(n4453 ,n4258 ,n4160);
    nor g4329(n913 ,n1[6] ,n2[6]);
    nand g4330(n921 ,n0[34] ,n725);
    nand g4331(n1795 ,n0[80] ,n1023);
    nand g4332(n3618 ,n1[61] ,n3003);
    nor g4333(n1767 ,n1223 ,n1242);
    nand g4334(n6827 ,n6824 ,n6823);
    nand g4335(n1807 ,n0[1] ,n1221);
    nand g4336(n4396 ,n709 ,n4234);
    xnor g4337(n2717 ,n1[59] ,n1486);
    nor g4338(n958 ,n0[44] ,n790);
    nand g4339(n10[3] ,n4932 ,n4712);
    xnor g4340(n1297 ,n0[64] ,n1[80]);
    nor g4341(n6583 ,n0[115] ,n0[83]);
    nand g4342(n6400 ,n5910 ,n6340);
    or g4343(n6479 ,n6393 ,n6421);
    xnor g4344(n4924 ,n2845 ,n4446);
    nor g4345(n1751 ,n0[90] ,n1018);
    xnor g4346(n547 ,n6960 ,n0[103]);
    nand g4347(n6499 ,n6366 ,n703);
    xnor g4348(n5016 ,n4098 ,n4809);
    xnor g4349(n5960 ,n5723 ,n1674);
    nor g4350(n5654 ,n4868 ,n5540);
    nor g4351(n862 ,n710 ,n0[60]);
    nor g4352(n2361 ,n721 ,n1555);
    nor g4353(n6069 ,n793 ,n5956);
    nand g4354(n1087 ,n0[60] ,n708);
    not g4355(n4821 ,n4820);
    nand g4356(n4083 ,n720 ,n3698);
    nand g4357(n2582 ,n0[10] ,n707);
    nand g4358(n1218 ,n1[55] ,n2[55]);
    nand g4359(n3619 ,n0[36] ,n2794);
    or g4360(n5954 ,n713 ,n5932);
    nand g4361(n9[4] ,n5821 ,n6007);
    not g4362(n2866 ,n2865);
    nand g4363(n3169 ,n2581 ,n2497);
    nor g4364(n6364 ,n6299 ,n6293);
    nand g4365(n5920 ,n4159 ,n5791);
    xnor g4366(n1303 ,n1[35] ,n4[27]);
    nand g4367(n6671 ,n1[67] ,n6580);
    nor g4368(n2195 ,n1958 ,n1634);
    nand g4369(n605 ,n508 ,n604);
    nor g4370(n4539 ,n1176 ,n4135);
    nor g4371(n4480 ,n3030 ,n4297);
    nand g4372(n1185 ,n6912 ,n795);
    nand g4373(n3477 ,n1964 ,n2717);
    nor g4374(n5678 ,n4415 ,n5540);
    not g4375(n5552 ,n5551);
    nand g4376(n5822 ,n5652 ,n5712);
    nand g4377(n3862 ,n2208 ,n3640);
    nor g4378(n3902 ,n789 ,n3800);
    nor g4379(n5114 ,n4667 ,n4881);
    or g4380(n4739 ,n3531 ,n4551);
    nand g4381(n7079 ,n668 ,n635);
    nand g4382(n7163 ,n6581 ,n7116);
    nor g4383(n3517 ,n2401 ,n3005);
    nand g4384(n4261 ,n720 ,n3826);
    xnor g4385(n5289 ,n4663 ,n4996);
    nor g4386(n4042 ,n3755 ,n3025);
    or g4387(n6049 ,n711 ,n6032);
    nand g4388(n5877 ,n717 ,n5839);
    nand g4389(n641 ,n0[88] ,n622);
    xnor g4390(n2679 ,n1666 ,n1622);
    nand g4391(n285 ,n205 ,n284);
    nand g4392(n3233 ,n1206 ,n2062);
    xnor g4393(n399 ,n6997 ,n7029);
    nand g4394(n1091 ,n0[44] ,n789);
    nor g4395(n3505 ,n6825 ,n2816);
    nor g4396(n5804 ,n5518 ,n5702);
    not g4397(n6581 ,n6826);
    nand g4398(n4970 ,n3008 ,n4627);
    xnor g4399(n1434 ,n1[76] ,n2[12]);
    xnor g4400(n1476 ,n1[102] ,n2[38]);
    xnor g4401(n6844 ,n544 ,n565);
    nand g4402(n139 ,n59 ,n138);
    nand g4403(n567 ,n514 ,n566);
    xnor g4404(n1261 ,n0[107] ,n7103);
    xnor g4405(n2915 ,n1646 ,n1518);
    or g4406(n2985 ,n2621 ,n2384);
    xnor g4407(n5244 ,n4424 ,n4879);
    nand g4408(n51 ,n7057 ,n0[1]);
    or g4409(n2979 ,n2627 ,n2386);
    nor g4410(n2969 ,n2618 ,n2390);
    nor g4411(n972 ,n724 ,n0[3]);
    xnor g4412(n1690 ,n1[118] ,n4[14]);
    nand g4413(n2522 ,n1101 ,n1727);
    nor g4414(n5930 ,n1954 ,n5747);
    nor g4415(n5493 ,n5122 ,n5387);
    nand g4416(n7133 ,n6661 ,n6719);
    nand g4417(n1230 ,n0[97] ,n0[96]);
    or g4418(n39 ,n7070 ,n0[14]);
    nor g4419(n6320 ,n1954 ,n6279);
    nor g4420(n3676 ,n761 ,n3088);
    nand g4421(n6953 ,n6753 ,n6784);
    xnor g4422(n1713 ,n0[37] ,n1[53]);
    nand g4423(n1232 ,n3[3] ,n3[0]);
    or g4424(n3040 ,n1816 ,n2491);
    nor g4425(n4159 ,n3735 ,n3846);
    nor g4426(n2147 ,n1956 ,n1572);
    or g4427(n2046 ,n1959 ,n1414);
    nand g4428(n5629 ,n5106 ,n5458);
    not g4429(n810 ,n0[72]);
    nor g4430(n2228 ,n6 ,n1978);
    nand g4431(n6783 ,n1[113] ,n7088);
    nand g4432(n4715 ,n3807 ,n4559);
    or g4433(n4388 ,n6 ,n4358);
    xnor g4434(n5588 ,n5201 ,n2650);
    nand g4435(n672 ,n1[20] ,n621);
    nor g4436(n3511 ,n1819 ,n3009);
    xnor g4437(n6943 ,n81 ,n157);
    nor g4438(n5753 ,n1954 ,n5595);
    xnor g4439(n2689 ,n1[112] ,n1566);
    nand g4440(n5396 ,n5240 ,n5239);
    nand g4441(n1058 ,n0[45] ,n788);
    not g4442(n1497 ,n1496);
    xnor g4443(n1652 ,n0[67] ,n1[83]);
    xnor g4444(n2814 ,n0[75] ,n1261);
    nor g4445(n5521 ,n4012 ,n5386);
    nand g4446(n6381 ,n3452 ,n6267);
    xnor g4447(n2853 ,n1309 ,n1332);
    nor g4448(n4505 ,n3577 ,n4325);
    nor g4449(n3860 ,n2770 ,n3779);
    xor g4450(n7104 ,n0[44] ,n0[12]);
    xnor g4451(n1289 ,n0[4] ,n4[20]);
    nand g4452(n3373 ,n1953 ,n2911);
    nor g4453(n6594 ,n0[117] ,n0[85]);
    nand g4454(n5397 ,n717 ,n5269);
    nand g4455(n9[113] ,n4419 ,n6397);
    or g4456(n2531 ,n1229 ,n1946);
    nand g4457(n6112 ,n5509 ,n5978);
    xnor g4458(n1474 ,n1[67] ,n2[3]);
    nand g4459(n2554 ,n1109 ,n1899);
    or g4460(n2774 ,n1506 ,n2621);
    xnor g4461(n3910 ,n1[86] ,n2714);
    nand g4462(n1069 ,n0[76] ,n793);
    nand g4463(n4325 ,n2601 ,n3919);
    nand g4464(n2472 ,n0[50] ,n718);
    nand g4465(n4456 ,n4255 ,n4208);
    nand g4466(n6062 ,n5790 ,n5994);
    nand g4467(n2419 ,n0[41] ,n718);
    nand g4468(n1139 ,n6941 ,n795);
    or g4469(n6149 ,n3348 ,n6042);
    or g4470(n2970 ,n2633 ,n2334);
    nand g4471(n3205 ,n1194 ,n2066);
    nor g4472(n3626 ,n2547 ,n2975);
    xnor g4473(n5943 ,n5722 ,n4810);
    nand g4474(n3890 ,n709 ,n3522);
    nor g4475(n5799 ,n5720 ,n5683);
    nand g4476(n4957 ,n3545 ,n4757);
    nand g4477(n5385 ,n4830 ,n5183);
    nor g4478(n3963 ,n3580 ,n3801);
    xnor g4479(n6873 ,n399 ,n427);
    nand g4480(n3786 ,n1953 ,n2953);
    nor g4481(n4386 ,n3204 ,n4269);
    nand g4482(n2573 ,n0[26] ,n707);
    or g4483(n4255 ,n710 ,n4116);
    xnor g4484(n1628 ,n0[90] ,n1[90]);
    nand g4485(n3675 ,n0[14] ,n3083);
    xnor g4486(n1251 ,n0[71] ,n7099);
    xnor g4487(n1684 ,n6866 ,n6867);
    nand g4488(n1896 ,n0[51] ,n1221);
    nor g4489(n6389 ,n1954 ,n6315);
    or g4490(n4716 ,n3518 ,n4560);
    or g4491(n5125 ,n722 ,n5006);
    nor g4492(n1750 ,n971 ,n1031);
    xor g4493(n7109 ,n0[49] ,n0[17]);
    xnor g4494(n4436 ,n2829 ,n3952);
    nor g4495(n4521 ,n3676 ,n4303);
    nand g4496(n3172 ,n1976 ,n2326);
    nand g4497(n6967 ,n6747 ,n6776);
    not g4498(n846 ,n6889);
    nand g4499(n1181 ,n6937 ,n796);
    xnor g4500(n1662 ,n0[40] ,n1[56]);
    xnor g4501(n1331 ,n0[39] ,n0[23]);
    nand g4502(n1121 ,n6887 ,n795);
    nand g4503(n7156 ,n6581 ,n7123);
    nor g4504(n3409 ,n1222 ,n2847);
    xor g4505(n7120 ,n0[60] ,n0[28]);
    nand g4506(n5249 ,n3313 ,n5054);
    nor g4507(n2173 ,n1958 ,n1947);
    not g4508(n6578 ,n7088);
    xnor g4509(n532 ,n6976 ,n0[119]);
    or g4510(n6141 ,n4597 ,n6069);
    xor g4511(n6833 ,n389 ,n376);
    nand g4512(n1889 ,n0[31] ,n1221);
    nor g4513(n1004 ,n820 ,n0[66]);
    or g4514(n188 ,n0[44] ,n1[44]);
    nand g4515(n4726 ,n2326 ,n4441);
    not g4516(n779 ,n1[51]);
    nand g4517(n2544 ,n1149 ,n1812);
    nor g4518(n3408 ,n1954 ,n2926);
    nand g4519(n3993 ,n0[39] ,n3490);
    nand g4520(n7015 ,n6664 ,n7158);
    nor g4521(n6020 ,n5900 ,n5919);
    or g4522(n338 ,n7028 ,n6996);
    nand g4523(n7138 ,n6646 ,n6714);
    xnor g4524(n1401 ,n1[42] ,n2[42]);
    not g4525(n782 ,n1[52]);
    nand g4526(n1171 ,n6884 ,n795);
    xnor g4527(n6911 ,n73 ,n141);
    nand g4528(n9[73] ,n4497 ,n6443);
    not g4529(n832 ,n0[109]);
    nor g4530(n6266 ,n713 ,n6248);
    nand g4531(n5533 ,n4702 ,n5309);
    nand g4532(n2036 ,n707 ,n1484);
    nand g4533(n5634 ,n3486 ,n5413);
    nand g4534(n292 ,n165 ,n291);
    nand g4535(n9[27] ,n6549 ,n6567);
    nand g4536(n3242 ,n7166 ,n2563);
    nand g4537(n3732 ,n6821 ,n3098);
    or g4538(n2765 ,n1533 ,n2632);
    nand g4539(n6130 ,n717 ,n6109);
    nor g4540(n868 ,n0[9] ,n0[8]);
    xnor g4541(n540 ,n0[127] ,n6984);
    nand g4542(n6536 ,n6486 ,n6503);
    nand g4543(n3670 ,n0[26] ,n3084);
    nand g4544(n1108 ,n6880 ,n796);
    nand g4545(n7145 ,n6628 ,n6707);
    nor g4546(n2377 ,n1[37] ,n719);
    xnor g4547(n4881 ,n4583 ,n4424);
    nand g4548(n1883 ,n0[21] ,n966);
    nor g4549(n6021 ,n3324 ,n5890);
    nand g4550(n5551 ,n4817 ,n5367);
    nor g4551(n5410 ,n713 ,n5269);
    nand g4552(n1063 ,n0[31] ,n708);
    nand g4553(n5163 ,n4242 ,n4856);
    nand g4554(n6355 ,n6295 ,n6294);
    nand g4555(n516 ,n0[102] ,n6959);
    nand g4556(n1214 ,n1[54] ,n2[54]);
    nand g4557(n7026 ,n6621 ,n7147);
    nor g4558(n3090 ,n1221 ,n2394);
    xnor g4559(n5889 ,n5640 ,n1500);
    xnor g4560(n3946 ,n1366 ,n2834);
    nor g4561(n2532 ,n1963 ,n1521);
    nor g4562(n4277 ,n4037 ,n4071);
    xnor g4563(n377 ,n7006 ,n7038);
    nand g4564(n4266 ,n720 ,n3830);
    or g4565(n3464 ,n1954 ,n2937);
    nand g4566(n6489 ,n6462 ,n6411);
    nand g4567(n6781 ,n1[112] ,n7088);
    not g4568(n741 ,n0[82]);
    nor g4569(n4251 ,n2325 ,n4108);
    xnor g4570(n1412 ,n1[59] ,n2[59]);
    xnor g4571(n1456 ,n0[111] ,n0[47]);
    nor g4572(n6258 ,n712 ,n6247);
    xnor g4573(n6944 ,n538 ,n615);
    nand g4574(n6226 ,n3402 ,n6118);
    nand g4575(n5892 ,n1955 ,n5834);
    or g4576(n3306 ,n1[34] ,n3146);
    nand g4577(n2599 ,n0[6] ,n707);
    xnor g4578(n4444 ,n2803 ,n3949);
    nand g4579(n5433 ,n3415 ,n5285);
    xnor g4580(n1498 ,n1[36] ,n1[4]);
    nand g4581(n1918 ,n714 ,n1228);
    not g4582(n4708 ,n4707);
    nand g4583(n3236 ,n1217 ,n2128);
    nand g4584(n666 ,n1[13] ,n621);
    nand g4585(n4939 ,n3551 ,n4724);
    not g4586(n4573 ,n4572);
    xnor g4587(n1365 ,n1[36] ,n4[28]);
    nand g4588(n5898 ,n3576 ,n5792);
    nand g4589(n5282 ,n4608 ,n5071);
    nand g4590(n9[71] ,n5678 ,n5692);
    xnor g4591(n1622 ,n0[109] ,n1[109]);
    nor g4592(n21 ,n7057 ,n0[1]);
    or g4593(n487 ,n0[105] ,n6962);
    nand g4594(n3700 ,n1[92] ,n2961);
    nor g4595(n6247 ,n5444 ,n6144);
    xnor g4596(n1312 ,n0[90] ,n7118);
    nand g4597(n154 ,n41 ,n153);
    nor g4598(n4975 ,n4332 ,n4731);
    nor g4599(n855 ,n0[100] ,n788);
    nand g4600(n5707 ,n2893 ,n5478);
    or g4601(n1786 ,n995 ,n1225);
    xnor g4602(n2677 ,n0[124] ,n1269);
    nand g4603(n3231 ,n1215 ,n2097);
    nor g4604(n4696 ,n6824 ,n4476);
    nand g4605(n3980 ,n3588 ,n2257);
    xnor g4606(n1924 ,n1[44] ,n2[44]);
    nand g4607(n4979 ,n4023 ,n4791);
    nand g4608(n4506 ,n3603 ,n4279);
    nand g4609(n3152 ,n1[85] ,n2343);
    nand g4610(n1106 ,n0[67] ,n0[64]);
    nor g4611(n4606 ,n713 ,n4573);
    or g4612(n3858 ,n787 ,n3519);
    nor g4613(n2378 ,n0[37] ,n719);
    xnor g4614(n378 ,n7007 ,n7039);
    nor g4615(n5812 ,n5519 ,n5613);
    nand g4616(n6666 ,n0[76] ,n6579);
    not g4617(n845 ,n6823);
    nand g4618(n214 ,n0[62] ,n1[62]);
    nand g4619(n4537 ,n1191 ,n4186);
    nand g4620(n673 ,n1[8] ,n621);
    nand g4621(n6662 ,n1[86] ,n6579);
    nor g4622(n4670 ,n2134 ,n4469);
    xnor g4623(n5596 ,n4845 ,n5275);
    nor g4624(n6409 ,n5153 ,n6360);
    nor g4625(n6606 ,n0[116] ,n0[84]);
    nand g4626(n6307 ,n4157 ,n6193);
    nand g4627(n1235 ,n0[9] ,n0[8]);
    nand g4628(n3593 ,n0[125] ,n2794);
    nor g4629(n2359 ,n1963 ,n1530);
    nor g4630(n2215 ,n2024 ,n1757);
    or g4631(n2306 ,n1961 ,n1477);
    nand g4632(n5224 ,n717 ,n5060);
    nor g4633(n4341 ,n3608 ,n4094);
    nand g4634(n2355 ,n707 ,n1503);
    nand g4635(n6638 ,n0[110] ,n0[78]);
    nand g4636(n5679 ,n3627 ,n5547);
    xnor g4637(n1306 ,n6913 ,n6912);
    xnor g4638(n6942 ,n233 ,n309);
    nand g4639(n7090 ,n3[1] ,n6731);
    nor g4640(n5620 ,n5083 ,n5460);
    nand g4641(n1093 ,n0[87] ,n788);
    nand g4642(n7065 ,n658 ,n627);
    nor g4643(n859 ,n709 ,n0[100]);
    nor g4644(n6147 ,n3230 ,n6095);
    nor g4645(n3447 ,n1954 ,n2954);
    nand g4646(n4976 ,n4022 ,n4813);
    nor g4647(n6572 ,n1954 ,n6563);
    nor g4648(n1730 ,n0[105] ,n1227);
    nor g4649(n3453 ,n1954 ,n2935);
    nand g4650(n1764 ,n723 ,n920);
    nor g4651(n4146 ,n1960 ,n3840);
    nand g4652(n3312 ,n1953 ,n2881);
    nor g4653(n2982 ,n1749 ,n2416);
    xnor g4654(n1379 ,n6861 ,n6860);
    xnor g4655(n6282 ,n5940 ,n6172);
    nand g4656(n6799 ,n1[104] ,n7088);
    nand g4657(n4972 ,n4031 ,n4746);
    nor g4658(n2785 ,n2444 ,n2498);
    xnor g4659(n2820 ,n0[106] ,n1252);
    nor g4660(n3899 ,n2554 ,n3713);
    xnor g4661(n2835 ,n1271 ,n1684);
    xnor g4662(n531 ,n6975 ,n0[118]);
    nor g4663(n4678 ,n794 ,n4422);
    nor g4664(n3607 ,n768 ,n2797);
    nand g4665(n9[93] ,n5255 ,n5822);
    nor g4666(n6014 ,n3354 ,n5871);
    nand g4667(n7031 ,n6636 ,n7142);
    xnor g4668(n5729 ,n4663 ,n5459);
    xnor g4669(n2680 ,n1699 ,n1582);
    nand g4670(n266 ,n192 ,n265);
    nor g4671(n2370 ,n0[47] ,n1958);
    nand g4672(n4762 ,n2560 ,n4468);
    xnor g4673(n2959 ,n1[125] ,n1567);
    nand g4674(n6612 ,n0[101] ,n0[69]);
    nand g4675(n6543 ,n1952 ,n704);
    nor g4676(n5717 ,n4091 ,n5553);
    nor g4677(n2340 ,n0[45] ,n1957);
    nor g4678(n3652 ,n729 ,n3079);
    nand g4679(n3118 ,n1[48] ,n2617);
    nor g4680(n6011 ,n3304 ,n5863);
    nor g4681(n3445 ,n1222 ,n2819);
    xnor g4682(n1610 ,n0[114] ,n1[114]);
    nand g4683(n3188 ,n1906 ,n2457);
    nand g4684(n7045 ,n6676 ,n7128);
    not g4685(n742 ,n0[16]);
    nand g4686(n6051 ,n1955 ,n6032);
    nor g4687(n4416 ,n6 ,n4214);
    nor g4688(n2648 ,n2277 ,n2095);
    nor g4689(n4997 ,n2116 ,n4672);
    not g4690(n5267 ,n5268);
    xnor g4691(n3948 ,n1719 ,n2831);
    nor g4692(n2155 ,n6 ,n1739);
    not g4693(n6338 ,n6337);
    nand g4694(n4802 ,n710 ,n4588);
    nand g4695(n875 ,n714 ,n728);
    nand g4696(n5628 ,n5536 ,n5406);
    nand g4697(n4096 ,n3244 ,n3688);
    nor g4698(n5738 ,n1954 ,n5576);
    xor g4699(n703 ,n6170 ,n6310);
    nor g4700(n3535 ,n6825 ,n2847);
    nand g4701(n7131 ,n6696 ,n6721);
    nand g4702(n204 ,n0[55] ,n1[55]);
    nand g4703(n3751 ,n7152 ,n3101);
    not g4704(n763 ,n1[48]);
    xnor g4705(n1567 ,n1[61] ,n1[29]);
    not g4706(n1957 ,n718);
    nand g4707(n5910 ,n3300 ,n5749);
    nor g4708(n1050 ,n708 ,n0[4]);
    or g4709(n2200 ,n1960 ,n1451);
    nor g4710(n1994 ,n861 ,n914);
    not g4711(n4694 ,n4693);
    nor g4712(n4793 ,n3641 ,n4563);
    nor g4713(n3002 ,n1[61] ,n2564);
    nand g4714(n2581 ,n0[27] ,n1964);
    nand g4715(n679 ,n1[30] ,n621);
    nand g4716(n4992 ,n2533 ,n4676);
    xnor g4717(n6872 ,n551 ,n579);
    not g4718(n726 ,n6825);
    or g4719(n2032 ,n912 ,n2029);
    xnor g4720(n1592 ,n0[76] ,n1[76]);
    not g4721(n5719 ,n5718);
    xnor g4722(n5456 ,n5154 ,n4467);
    nor g4723(n6551 ,n5545 ,n6518);
    nor g4724(n2374 ,n0[41] ,n719);
    nand g4725(n3210 ,n1130 ,n2080);
    nand g4726(n5226 ,n5104 ,n5059);
    nand g4727(n1149 ,n6871 ,n795);
    nand g4728(n5859 ,n1955 ,n5727);
    nand g4729(n6811 ,n6581 ,n7103);
    xnor g4730(n4477 ,n3939 ,n2817);
    nand g4731(n9[91] ,n5694 ,n6562);
    nand g4732(n6667 ,n1[88] ,n6580);
    nor g4733(n6078 ,n6013 ,n5989);
    not g4734(n799 ,n0[17]);
    not g4735(n775 ,n0[94]);
    xnor g4736(n2664 ,n1[104] ,n1539);
    nor g4737(n2158 ,n719 ,n1606);
    xnor g4738(n1666 ,n0[93] ,n4[21]);
    nand g4739(n4558 ,n1152 ,n4264);
    nand g4740(n6976 ,n6742 ,n6773);
    nand g4741(n6972 ,n6758 ,n6790);
    or g4742(n489 ,n0[104] ,n6961);
    nand g4743(n6002 ,n3443 ,n5894);
    nand g4744(n962 ,n0[30] ,n789);
    nand g4745(n265 ,n207 ,n264);
    nor g4746(n5346 ,n4715 ,n5186);
    nand g4747(n10[23] ,n4764 ,n5343);
    nand g4748(n1099 ,n0[15] ,n0[7]);
    nand g4749(n6506 ,n4726 ,n6440);
    not g4750(n819 ,n0[10]);
    not g4751(n4919 ,n4918);
    or g4752(n328 ,n7043 ,n7011);
    nand g4753(n4018 ,n3623 ,n3491);
    nor g4754(n5334 ,n3509 ,n5135);
    nand g4755(n3660 ,n2482 ,n2968);
    nand g4756(n4655 ,n4010 ,n4373);
    nor g4757(n6099 ,n6027 ,n5983);
    nand g4758(n9[28] ,n5227 ,n6061);
    xnor g4759(n2850 ,n0[115] ,n1373);
    nand g4760(n4642 ,n794 ,n4441);
    nand g4761(n566 ,n470 ,n565);
    xnor g4762(n3818 ,n2693 ,n2676);
    nand g4763(n4861 ,n3470 ,n4601);
    xnor g4764(n5731 ,n5390 ,n4461);
    nand g4765(n1010 ,n0[40] ,n808);
    nor g4766(n2271 ,n721 ,n1490);
    nor g4767(n3478 ,n1954 ,n2947);
    or g4768(n6117 ,n706 ,n6066);
    nand g4769(n366 ,n7048 ,n7016);
    nand g4770(n3761 ,n7138 ,n3045);
    nand g4771(n4278 ,n0[37] ,n3908);
    nor g4772(n1770 ,n724 ,n1001);
    nor g4773(n5786 ,n5049 ,n5720);
    xnor g4774(n2649 ,n2002 ,n1994);
    xnor g4775(n2937 ,n1676 ,n1636);
    nor g4776(n5179 ,n6824 ,n4926);
    nand g4777(n418 ,n344 ,n417);
    nor g4778(n6009 ,n5604 ,n5929);
    or g4779(n3049 ,n1236 ,n2325);
    nor g4780(n1866 ,n740 ,n977);
    nand g4781(n3708 ,n776 ,n3177);
    nor g4782(n6584 ,n0[108] ,n0[76]);
    or g4783(n5423 ,n4998 ,n5277);
    nor g4784(n907 ,n1[123] ,n2[59]);
    nand g4785(n4056 ,n2767 ,n3651);
    nand g4786(n6694 ,n0[80] ,n6580);
    not g4787(n730 ,n0[73]);
    xnor g4788(n1307 ,n0[118] ,n0[6]);
    xnor g4789(n383 ,n7012 ,n7044);
    nand g4790(n2542 ,n1198 ,n1833);
    nor g4791(n4805 ,n2285 ,n4470);
    xnor g4792(n2841 ,n1372 ,n1701);
    nand g4793(n3780 ,n1196 ,n3179);
    xnor g4794(n6855 ,n90 ,n113);
    nand g4795(n2625 ,n761 ,n707);
    nor g4796(n3468 ,n2299 ,n3029);
    xnor g4797(n1487 ,n0[1] ,n1[1]);
    xnor g4798(n1886 ,n1[86] ,n2[22]);
    nand g4799(n3741 ,n6813 ,n3052);
    nand g4800(n3632 ,n1[38] ,n2775);
    or g4801(n1743 ,n0[113] ,n987);
    not g4802(n4914 ,n4913);
    xnor g4803(n2912 ,n1662 ,n1560);
    or g4804(n3275 ,n2759 ,n3208);
    nand g4805(n3340 ,n1952 ,n2894);
    xnor g4806(n2672 ,n1[111] ,n1493);
    nor g4807(n2454 ,n721 ,n1640);
    xnor g4808(n1709 ,n0[72] ,n4[0]);
    nor g4809(n5297 ,n794 ,n5056);
    nand g4810(n9[75] ,n5109 ,n6550);
    nand g4811(n9[88] ,n5496 ,n6530);
    nor g4812(n2394 ,n1963 ,n1529);
    nand g4813(n1228 ,n0[26] ,n0[24]);
    nor g4814(n4858 ,n3266 ,n4700);
    xnor g4815(n6927 ,n77 ,n149);
    nor g4816(n4709 ,n6824 ,n689);
    nand g4817(n2494 ,n0[53] ,n718);
    xnor g4818(n2842 ,n0[81] ,n1274);
    xnor g4819(n1885 ,n1[127] ,n2[63]);
    nand g4820(n3973 ,n0[5] ,n3491);
    nor g4821(n4200 ,n6 ,n4101);
    nand g4822(n3459 ,n710 ,n2963);
    not g4823(n2794 ,n2795);
    nand g4824(n3689 ,n838 ,n3155);
    nor g4825(n5511 ,n722 ,n5378);
    or g4826(n3319 ,n1954 ,n2883);
    xnor g4827(n1541 ,n0[62] ,n4[22]);
    nor g4828(n3530 ,n6825 ,n2849);
    nand g4829(n4548 ,n1143 ,n4167);
    xnor g4830(n1253 ,n6925 ,n6924);
    nand g4831(n68 ,n7082 ,n0[26]);
    nand g4832(n1978 ,n1091 ,n1213);
    nand g4833(n1135 ,n6932 ,n796);
    nand g4834(n5211 ,n4949 ,n5080);
    nand g4835(n635 ,n0[87] ,n622);
    or g4836(n3010 ,n2164 ,n2236);
    not g4837(n786 ,n6913);
    nor g4838(n2987 ,n0[48] ,n2193);
    xnor g4839(n2905 ,n1286 ,n1325);
    nand g4840(n5169 ,n717 ,n4992);
    nor g4841(n6311 ,n4416 ,n6192);
    xnor g4842(n1927 ,n1[14] ,n2[14]);
    nand g4843(n3933 ,n2148 ,n3632);
    or g4844(n3437 ,n1954 ,n2932);
    xnor g4845(n1605 ,n0[92] ,n1[92]);
    xnor g4846(n1252 ,n0[74] ,n7102);
    nor g4847(n5907 ,n5419 ,n5785);
    xnor g4848(n5201 ,n4994 ,n4999);
    nand g4849(n1101 ,n0[69] ,n0[13]);
    xnor g4850(n1686 ,n0[89] ,n4[17]);
    nand g4851(n4928 ,n4239 ,n4609);
    xnor g4852(n552 ,n6965 ,n0[108]);
    xnor g4853(n2652 ,n1588 ,n1549);
    nand g4854(n1811 ,n0[43] ,n1221);
    nor g4855(n1047 ,n725 ,n0[35]);
    nand g4856(n4049 ,n3631 ,n2036);
    nand g4857(n3198 ,n1246 ,n2578);
    nand g4858(n3787 ,n6815 ,n3240);
    nand g4859(n4929 ,n3013 ,n4650);
    nand g4860(n7008 ,n6670 ,n7165);
    or g4861(n2148 ,n1962 ,n1416);
    xnor g4862(n6914 ,n226 ,n295);
    xnor g4863(n2960 ,n1708 ,n1581);
    nand g4864(n4557 ,n1181 ,n4141);
    nor g4865(n2233 ,n708 ,n1608);
    nand g4866(n1969 ,n1058 ,n928);
    nand g4867(n3379 ,n1953 ,n2915);
    nand g4868(n7061 ,n683 ,n651);
    nand g4869(n5500 ,n4684 ,n5311);
    nand g4870(n4511 ,n3708 ,n4179);
    nor g4871(n6255 ,n5999 ,n6216);
    xnor g4872(n1546 ,n0[60] ,n4[20]);
    nor g4873(n4038 ,n3747 ,n3010);
    nor g4874(n1819 ,n0[24] ,n1040);
    not g4875(n5550 ,n5549);
    nor g4876(n6380 ,n3293 ,n6266);
    xnor g4877(n244 ,n1[40] ,n0[40]);
    nand g4878(n3569 ,n1952 ,n2957);
    nand g4879(n1002 ,n0[98] ,n754);
    nand g4880(n4538 ,n1163 ,n4134);
    nand g4881(n5561 ,n4815 ,n5368);
    xnor g4882(n388 ,n7049 ,n7017);
    nor g4883(n5836 ,n3487 ,n5641);
    xnor g4884(n248 ,n1[44] ,n0[44]);
    xnor g4885(n4408 ,n3812 ,n1993);
    nor g4886(n2125 ,n1963 ,n1638);
    nor g4887(n5097 ,n712 ,n4993);
    nand g4888(n1078 ,n0[14] ,n708);
    nand g4889(n278 ,n188 ,n277);
    nor g4890(n4171 ,n3724 ,n3934);
    nor g4891(n2386 ,n0[51] ,n719);
    xnor g4892(n2665 ,n1[103] ,n1561);
    xnor g4893(n5210 ,n5000 ,n1347);
    nand g4894(n6682 ,n0[87] ,n6580);
    nand g4895(n2436 ,n919 ,n1787);
    nor g4896(n923 ,n0[70] ,n715);
    xnor g4897(n395 ,n6993 ,n7025);
    xnor g4898(n1264 ,n0[109] ,n4[5]);
    nor g4899(n5958 ,n706 ,n5933);
    nand g4900(n611 ,n524 ,n610);
    xnor g4901(n1437 ,n1[8] ,n2[8]);
    nor g4902(n4120 ,n715 ,n4115);
    nand g4903(n138 ,n15 ,n137);
    nand g4904(n6760 ,n0[59] ,n6737);
    nor g4905(n6154 ,n6104 ,n6077);
    nor g4906(n2620 ,n0[15] ,n1963);
    or g4907(n2050 ,n909 ,n2020);
    nor g4908(n2627 ,n0[19] ,n1963);
    xnor g4909(n2833 ,n0[122] ,n1312);
    nor g4910(n3866 ,n3041 ,n3780);
    nand g4911(n895 ,n0[73] ,n739);
    or g4912(n4745 ,n3530 ,n4536);
    nand g4913(n4801 ,n4326 ,n4495);
    nand g4914(n3170 ,n1996 ,n2326);
    nor g4915(n3510 ,n1222 ,n2812);
    xnor g4916(n1674 ,n0[95] ,n4[23]);
    nand g4917(n524 ,n0[122] ,n6979);
    nor g4918(n3115 ,n754 ,n2328);
    nand g4919(n3636 ,n1[52] ,n2736);
    nor g4920(n3015 ,n2141 ,n2256);
    nor g4921(n5839 ,n4193 ,n5641);
    nor g4922(n3332 ,n1954 ,n2869);
    or g4923(n1012 ,n0[26] ,n0[24]);
    nor g4924(n5657 ,n5558 ,n5428);
    nor g4925(n3578 ,n941 ,n2987);
    nor g4926(n2362 ,n721 ,n1552);
    nand g4927(n1773 ,n714 ,n1015);
    nor g4928(n6410 ,n3308 ,n6321);
    not g4929(n4673 ,n4672);
    or g4930(n2074 ,n719 ,n1556);
    xnor g4931(n1397 ,n1[38] ,n2[38]);
    or g4932(n4620 ,n2561 ,n4455);
    xnor g4933(n5592 ,n5263 ,n2654);
    or g4934(n3035 ,n2532 ,n2175);
    not g4935(n767 ,n0[125]);
    xnor g4936(n6935 ,n79 ,n153);
    nor g4937(n4336 ,n821 ,n4110);
    nand g4938(n9[2] ,n6054 ,n6407);
    or g4939(n3245 ,n1[40] ,n2603);
    nor g4940(n6720 ,n6826 ,n6596);
    nand g4941(n5037 ,n960 ,n5014);
    nand g4942(n451 ,n350 ,n450);
    nand g4943(n3119 ,n1[59] ,n2331);
    nor g4944(n1893 ,n765 ,n1223);
    nor g4945(n5495 ,n3566 ,n5286);
    nand g4946(n352 ,n7035 ,n7003);
    xnor g4947(n1455 ,n1[97] ,n2[33]);
    xnor g4948(n6897 ,n405 ,n439);
    not g4949(n843 ,n1[38]);
    nor g4950(n881 ,n0[107] ,n0[106]);
    nand g4951(n3634 ,n1[43] ,n2970);
    xnor g4952(n87 ,n0[3] ,n7059);
    or g4953(n41 ,n7082 ,n0[26]);
    nand g4954(n2357 ,n1964 ,n1495);
    xnor g4955(n1416 ,n1[70] ,n2[6]);
    nand g4956(n7082 ,n657 ,n624);
    not g4957(n1963 ,n1964);
    or g4958(n3360 ,n2052 ,n3106);
    nand g4959(n4482 ,n3611 ,n4267);
    nor g4960(n3050 ,n2027 ,n2325);
    nand g4961(n2966 ,n1218 ,n2449);
    or g4962(n4724 ,n713 ,n4575);
    nor g4963(n5443 ,n5217 ,n5290);
    or g4964(n3543 ,n0[65] ,n3196);
    nor g4965(n1818 ,n810 ,n11);
    or g4966(n5667 ,n2893 ,n5479);
    nor g4967(n2294 ,n901 ,n1959);
    nor g4968(n2321 ,n1957 ,n1913);
    xnor g4969(n1584 ,n0[103] ,n1[103]);
    or g4970(n9[56] ,n4483 ,n6554);
    xnor g4971(n403 ,n7001 ,n7033);
    or g4972(n2142 ,n719 ,n1585);
    nand g4973(n4730 ,n2326 ,n4452);
    xnor g4974(n4440 ,n2850 ,n3955);
    xnor g4975(n2712 ,n1[114] ,n1503);
    nor g4976(n5139 ,n727 ,n4904);
    nor g4977(n4175 ,n2549 ,n3936);
    nor g4978(n3193 ,n1972 ,n722);
    xnor g4979(n2945 ,n1689 ,n1583);
    xnor g4980(n1682 ,n7054 ,n7055);
    xnor g4981(n243 ,n1[39] ,n0[39]);
    xor g4982(n7107 ,n0[47] ,n0[15]);
    nand g4983(n4654 ,n4009 ,n4374);
    xnor g4984(n5215 ,n4661 ,n4878);
    xnor g4985(n387 ,n7016 ,n7048);
    not g4986(n2899 ,n2898);
    nor g4987(n4032 ,n3734 ,n2780);
    xnor g4988(n1459 ,n1[62] ,n2[62]);
    nor g4989(n4204 ,n715 ,n3964);
    nor g4990(n3869 ,n2179 ,n3303);
    nand g4991(n4063 ,n787 ,n3795);
    nor g4992(n3927 ,n3104 ,n3684);
    nand g4993(n4763 ,n2560 ,n4458);
    nand g4994(n3683 ,n1[42] ,n2969);
    nand g4995(n3725 ,n1202 ,n3048);
    nand g4996(n1200 ,n6919 ,n795);
    not g4997(n5184 ,n5183);
    nor g4998(n3876 ,n3331 ,n3330);
    nand g4999(n6241 ,n4786 ,n6150);
    nor g5000(n6227 ,n3289 ,n6115);
    nor g5001(n2366 ,n721 ,n1565);
    nor g5002(n5792 ,n5477 ,n5709);
    nand g5003(n6539 ,n6472 ,n6496);
    nand g5004(n1950 ,n3[3] ,n973);
    xnor g5005(n4595 ,n4106 ,n4217);
    nor g5006(n4486 ,n4271 ,n3506);
    nor g5007(n4420 ,n4346 ,n4095);
    nand g5008(n4259 ,n715 ,n4117);
    nor g5009(n1758 ,n725 ,n1011);
    nand g5010(n3171 ,n1975 ,n2326);
    nand g5011(n7058 ,n676 ,n646);
    nand g5012(n1174 ,n6860 ,n795);
    nand g5013(n290 ,n167 ,n289);
    nand g5014(n586 ,n495 ,n585);
    xnor g5015(n1677 ,n6870 ,n6871);
    not g5016(n762 ,n0[47]);
    nand g5017(n2550 ,n1116 ,n1832);
    not g5018(n2642 ,n2641);
    nand g5019(n3246 ,n925 ,n2040);
    xnor g5020(n4439 ,n2852 ,n3958);
    or g5021(n3455 ,n1954 ,n2934);
    nand g5022(n1119 ,n6829 ,n796);
    nand g5023(n2427 ,n0[113] ,n1736);
    nand g5024(n355 ,n7019 ,n6987);
    nand g5025(n595 ,n515 ,n594);
    nand g5026(n5874 ,n1952 ,n5732);
    xnor g5027(n2946 ,n1297 ,n1494);
    xnor g5028(n1499 ,n1[44] ,n1[12]);
    nand g5029(n1072 ,n0[38] ,n710);
    nor g5030(n4219 ,n3278 ,n3978);
    nor g5031(n3782 ,n1954 ,n2899);
    nor g5032(n6714 ,n6826 ,n6591);
    not g5033(n740 ,n0[121]);
    nor g5034(n4641 ,n6 ,n4584);
    nand g5035(n1976 ,n1093 ,n943);
    nor g5036(n6597 ,n0[105] ,n0[73]);
    nand g5037(n1138 ,n6837 ,n796);
    nor g5038(n3005 ,n724 ,n2210);
    nand g5039(n4054 ,n3020 ,n3650);
    nor g5040(n5566 ,n4824 ,n5356);
    nand g5041(n311 ,n196 ,n310);
    nand g5042(n107 ,n57 ,n106);
    nand g5043(n123 ,n70 ,n122);
    xor g5044(n6831 ,n0[0] ,n7056);
    nand g5045(n7068 ,n663 ,n633);
    xnor g5046(n1283 ,n0[69] ,n7097);
    nand g5047(n578 ,n490 ,n577);
    nor g5048(n5331 ,n4344 ,n5167);
    nor g5049(n2206 ,n1960 ,n1463);
    nand g5050(n1080 ,n0[108] ,n790);
    nor g5051(n3098 ,n1850 ,n2099);
    xnor g5052(n1453 ,n0[5] ,n1[37]);
    nand g5053(n108 ,n32 ,n107);
    nand g5054(n120 ,n31 ,n119);
    nor g5055(n2451 ,n1956 ,n1609);
    nand g5056(n3227 ,n1193 ,n2074);
    nand g5057(n6537 ,n5788 ,n6475);
    nand g5058(n7167 ,n6581 ,n7112);
    nand g5059(n10[31] ,n4634 ,n4867);
    nand g5060(n3609 ,n1229 ,n2998);
    nand g5061(n6095 ,n4288 ,n5962);
    not g5062(n764 ,n0[76]);
    xnor g5063(n6339 ,n5640 ,n6190);
    nor g5064(n949 ,n1[7] ,n2[7]);
    xnor g5065(n1670 ,n6950 ,n6951);
    nand g5066(n5468 ,n4692 ,n5334);
    or g5067(n36 ,n7068 ,n0[12]);
    not g5068(n744 ,n0[113]);
    nor g5069(n6569 ,n5503 ,n6553);
    nand g5070(n4556 ,n1187 ,n4266);
    nand g5071(n9[109] ,n5744 ,n5912);
    nand g5072(n4756 ,n717 ,n4575);
    nand g5073(n5190 ,n4240 ,n4933);
    not g5074(n4882 ,n4881);
    nand g5075(n1128 ,n6985 ,n796);
    nand g5076(n257 ,n203 ,n256);
    nand g5077(n2517 ,n793 ,n1990);
    or g5078(n167 ,n0[50] ,n1[50]);
    nor g5079(n5048 ,n4693 ,n4872);
    nand g5080(n1223 ,n0[56] ,n714);
    nand g5081(n3446 ,n1953 ,n2933);
    nor g5082(n5429 ,n706 ,n5270);
    nand g5083(n124 ,n12 ,n123);
    nor g5084(n3879 ,n2371 ,n3490);
    xnor g5085(n6883 ,n97 ,n127);
    nand g5086(n6365 ,n5996 ,n6281);
    xnor g5087(n5639 ,n5296 ,n4368);
    xnor g5088(n1343 ,n1[116] ,n4[12]);
    nand g5089(n3491 ,n1963 ,n2795);
    nor g5090(n6405 ,n5440 ,n6353);
    xnor g5091(n1944 ,n1[103] ,n2[39]);
    nor g5092(n2403 ,n1[36] ,n719);
    xor g5093(n6829 ,n6986 ,n7018);
    nand g5094(n4790 ,n4532 ,n4401);
    nand g5095(n4099 ,n3678 ,n3564);
    nand g5096(n7048 ,n6689 ,n7125);
    nor g5097(n5357 ,n3537 ,n5138);
    nor g5098(n5526 ,n4290 ,n5353);
    nor g5099(n6590 ,n0[103] ,n0[71]);
    or g5100(n3871 ,n2133 ,n3497);
    xnor g5101(n6926 ,n229 ,n301);
    nand g5102(n125 ,n71 ,n124);
    nor g5103(n2123 ,n1961 ,n1885);
    xnor g5104(n1649 ,n0[35] ,n0[19]);
    or g5105(n3625 ,n1954 ,n2861);
    nor g5106(n6717 ,n6826 ,n6606);
    nor g5107(n3937 ,n2272 ,n3732);
    nand g5108(n2587 ,n0[3] ,n707);
    nor g5109(n1203 ,n786 ,n716);
    nor g5110(n2400 ,n1[46] ,n1958);
    or g5111(n2772 ,n1535 ,n2624);
    nor g5112(n6591 ,n0[113] ,n0[81]);
    nor g5113(n5661 ,n3728 ,n5563);
    not g5114(n3940 ,n3939);
    nor g5115(n5106 ,n706 ,n4991);
    nor g5116(n4389 ,n4345 ,n3997);
    nand g5117(n5013 ,n2172 ,n4779);
    xnor g5118(n1847 ,n0[3] ,n811);
    xor g5119(n3824 ,n2664 ,n1[72]);
    nor g5120(n856 ,n1[54] ,n2[54]);
    nor g5121(n5158 ,n2090 ,n4884);
    nand g5122(n6645 ,n1[80] ,n6579);
    nor g5123(n3554 ,n1954 ,n2957);
    or g5124(n4068 ,n3671 ,n3501);
    not g5125(n4234 ,n4233);
    nand g5126(n2577 ,n0[28] ,n707);
    nand g5127(n6698 ,n1[65] ,n6580);
    nor g5128(n477 ,n0[97] ,n6954);
    nand g5129(n9[125] ,n5306 ,n5882);
    nand g5130(n4280 ,n792 ,n4108);
    xnor g5131(n1442 ,n1[124] ,n2[60]);
    nand g5132(n7018 ,n6674 ,n7155);
    nand g5133(n628 ,n0[85] ,n622);
    not g5134(n765 ,n0[57]);
    nor g5135(n909 ,n734 ,n0[73]);
    xnor g5136(n5783 ,n5374 ,n5463);
    nand g5137(n6741 ,n0[43] ,n6737);
    or g5138(n490 ,n0[106] ,n6963);
    nand g5139(n6801 ,n1[97] ,n7088);
    or g5140(n9[38] ,n4501 ,n5828);
    or g5141(n4489 ,n3239 ,n4287);
    nand g5142(n5896 ,n717 ,n5837);
    nand g5143(n6993 ,n6633 ,n6815);
    nand g5144(n3703 ,n779 ,n3168);
    nand g5145(n3239 ,n7165 ,n2566);
    nand g5146(n67 ,n7081 ,n0[25]);
    xnor g5147(n2955 ,n1621 ,n1524);
    xnor g5148(n1443 ,n1[2] ,n2[2]);
    nor g5149(n5238 ,n3546 ,n5177);
    xnor g5150(n6904 ,n559 ,n595);
    nor g5151(n5040 ,n727 ,n4926);
    nor g5152(n5735 ,n711 ,n5583);
    xnor g5153(n1912 ,n1[51] ,n2[51]);
    not g5154(n2864 ,n2863);
    not g5155(n6733 ,n7090);
    nor g5156(n2168 ,n1959 ,n1430);
    nor g5157(n2278 ,n1956 ,n1607);
    nand g5158(n3147 ,n1[117] ,n2399);
    xnor g5159(n1348 ,n1[37] ,n4[29]);
    or g5160(n5702 ,n5026 ,n5559);
    or g5161(n180 ,n0[34] ,n1[34]);
    nand g5162(n6527 ,n6480 ,n6499);
    nand g5163(n1109 ,n7055 ,n796);
    not g5164(n982 ,n983);
    xnor g5165(n5469 ,n4805 ,n5060);
    nor g5166(n4228 ,n793 ,n3836);
    nand g5167(n1113 ,n6936 ,n796);
    nand g5168(n6326 ,n1955 ,n6308);
    nor g5169(n6363 ,n6300 ,n6297);
    nand g5170(n213 ,n0[39] ,n1[39]);
    nor g5171(n5632 ,n3411 ,n5410);
    nor g5172(n1817 ,n807 ,n1220);
    xnor g5173(n1618 ,n0[121] ,n1[121]);
    nor g5174(n2224 ,n1959 ,n1423);
    nand g5175(n1215 ,n1[115] ,n2[51]);
    nand g5176(n629 ,n0[74] ,n622);
    nand g5177(n2578 ,n1235 ,n1911);
    nand g5178(n1231 ,n0[35] ,n0[34]);
    nand g5179(n4097 ,n2966 ,n3809);
    nor g5180(n3271 ,n1222 ,n2817);
    xnor g5181(n4890 ,n4568 ,n4582);
    or g5182(n3031 ,n2302 ,n2301);
    nor g5183(n4117 ,n2783 ,n3705);
    nand g5184(n6770 ,n1[114] ,n7088);
    nand g5185(n4467 ,n2230 ,n4216);
    nor g5186(n2266 ,n1963 ,n1526);
    nand g5187(n9[89] ,n5497 ,n6363);
    nor g5188(n5641 ,n794 ,n5449);
    nor g5189(n5663 ,n5416 ,n5525);
    nand g5190(n4748 ,n708 ,n4589);
    nor g5191(n2131 ,n1960 ,n1929);
    nand g5192(n10[18] ,n4766 ,n5338);
    nand g5193(n6676 ,n1[91] ,n6580);
    nand g5194(n9[122] ,n4525 ,n6183);
    nand g5195(n6665 ,n1[87] ,n6579);
    not g5196(n2925 ,n2924);
    nor g5197(n3872 ,n3311 ,n3310);
    nor g5198(n3924 ,n787 ,n3792);
    nand g5199(n10[12] ,n4771 ,n5348);
    xnor g5200(n2837 ,n1254 ,n1276);
    nand g5201(n3104 ,n7167 ,n2569);
    xnor g5202(n1613 ,n0[99] ,n1[99]);
    nand g5203(n5606 ,n5107 ,n5487);
    xnor g5204(n5855 ,n5001 ,n5569);
    nor g5205(n1841 ,n753 ,n1220);
    nand g5206(n577 ,n522 ,n576);
    nand g5207(n6792 ,n1[100] ,n7088);
    nor g5208(n5127 ,n3507 ,n4947);
    xnor g5209(n1945 ,n1[105] ,n2[41]);
    xnor g5210(n3941 ,n2677 ,n2813);
    nand g5211(n4313 ,n3024 ,n4050);
    nand g5212(n5221 ,n4961 ,n5079);
    not g5213(n1220 ,n1221);
    xnor g5214(n227 ,n1[54] ,n0[54]);
    nor g5215(n5808 ,n5557 ,n5620);
    nand g5216(n3520 ,n2982 ,n2980);
    nand g5217(n1986 ,n1079 ,n1063);
    not g5218(n6420 ,n6419);
    nand g5219(n1070 ,n0[109] ,n789);
    nand g5220(n9[99] ,n4034 ,n6569);
    not g5221(n1959 ,n720);
    nor g5222(n3544 ,n1222 ,n2853);
    nand g5223(n9[60] ,n5733 ,n6029);
    nand g5224(n604 ,n494 ,n603);
    nor g5225(n2402 ,n0[56] ,n719);
    nand g5226(n305 ,n219 ,n304);
    nor g5227(n3581 ,n740 ,n2981);
    nand g5228(n6163 ,n6081 ,n6096);
    xnor g5229(n6836 ,n542 ,n561);
    nand g5230(n4954 ,n794 ,n4680);
    xnor g5231(n1714 ,n6894 ,n6895);
    nor g5232(n3121 ,n1884 ,n2044);
    or g5233(n2775 ,n2641 ,n2388);
    xnor g5234(n1452 ,n1[77] ,n2[13]);
    nor g5235(n3265 ,n1781 ,n3253);
    nand g5236(n6796 ,n1[116] ,n7088);
    nor g5237(n886 ,n731 ,n0[105]);
    nor g5238(n5024 ,n712 ,n4875);
    xnor g5239(n1424 ,n1[20] ,n2[20]);
    nand g5240(n501 ,n0[108] ,n6965);
    xnor g5241(n250 ,n1[46] ,n0[46]);
    nand g5242(n6193 ,n6 ,n6119);
    nand g5243(n975 ,n0[19] ,n714);
    nand g5244(n283 ,n202 ,n282);
    nand g5245(n152 ,n24 ,n151);
    nor g5246(n2044 ,n1998 ,n2014);
    nand g5247(n5615 ,n5421 ,n5420);
    nor g5248(n5246 ,n3368 ,n5021);
    nand g5249(n1195 ,n6899 ,n795);
    nand g5250(n6040 ,n1955 ,n5974);
    nand g5251(n3146 ,n2591 ,n2446);
    nor g5252(n6015 ,n3377 ,n5872);
    nor g5253(n5150 ,n727 ,n4923);
    xnor g5254(n1536 ,n0[51] ,n4[11]);
    nor g5255(n4090 ,n6803 ,n3727);
    not g5256(n711 ,n717);
    xor g5257(n4922 ,n4444 ,n2804);
    nand g5258(n2497 ,n0[59] ,n718);
    nand g5259(n1970 ,n1071 ,n1089);
    nor g5260(n2734 ,n0[1] ,n2568);
    xnor g5261(n2898 ,n1358 ,n1614);
    nand g5262(n3989 ,n0[21] ,n3490);
    xnor g5263(n1335 ,n0[121] ,n4[9]);
    or g5264(n5054 ,n713 ,n4874);
    or g5265(n169 ,n0[59] ,n1[59]);
    or g5266(n6126 ,n706 ,n6109);
    nor g5267(n3421 ,n2325 ,n2808);
    xnor g5268(n4879 ,n4583 ,n4575);
    nand g5269(n3988 ,n3598 ,n2245);
    nand g5270(n5755 ,n4695 ,n5644);
    xnor g5271(n2700 ,n1971 ,n1978);
    nand g5272(n412 ,n336 ,n411);
    or g5273(n319 ,n7036 ,n7004);
    nand g5274(n675 ,n1[28] ,n621);
    or g5275(n6478 ,n6410 ,n6416);
    xnor g5276(n1717 ,n0[45] ,n1[61]);
    xnor g5277(n5066 ,n4424 ,n4807);
    nand g5278(n7127 ,n6681 ,n6725);
    nand g5279(n6358 ,n6277 ,n6271);
    xnor g5280(n2657 ,n1[127] ,n1311);
    nand g5281(n464 ,n333 ,n463);
    nand g5282(n3241 ,n6807 ,n2602);
    nor g5283(n2487 ,n1957 ,n1460);
    nor g5284(n5317 ,n4740 ,n5179);
    nor g5285(n5351 ,n3424 ,n5073);
    not g5286(n806 ,n0[83]);
    nor g5287(n2310 ,n1957 ,n1624);
    nand g5288(n6996 ,n6654 ,n6812);
    or g5289(n5257 ,n4206 ,n5167);
    nor g5290(n4181 ,n3226 ,n3930);
    nand g5291(n7043 ,n6701 ,n7130);
    nor g5292(n6162 ,n3471 ,n6043);
    nand g5293(n4279 ,n0[85] ,n3918);
    xnor g5294(n2686 ,n0[111] ,n1627);
    nand g5295(n6691 ,n0[127] ,n0[95]);
    or g5296(n5427 ,n5107 ,n5266);
    nor g5297(n2330 ,n1[118] ,n1957);
    or g5298(n3926 ,n708 ,n3520);
    nand g5299(n5535 ,n4831 ,n5358);
    nand g5300(n6977 ,n6746 ,n6777);
    nand g5301(n589 ,n509 ,n588);
    nand g5302(n4531 ,n2326 ,n4225);
    nor g5303(n2099 ,n1958 ,n1604);
    nand g5304(n2395 ,n1964 ,n1574);
    nand g5305(n6637 ,n0[102] ,n0[70]);
    not g5306(n5457 ,n5456);
    or g5307(n4626 ,n3537 ,n4548);
    not g5308(n754 ,n0[97]);
    nor g5309(n2315 ,n1962 ,n1420);
    nand g5310(n6751 ,n0[48] ,n6737);
    not g5311(n6214 ,n6213);
    xnor g5312(n2811 ,n0[108] ,n1313);
    xnor g5313(n1557 ,n1[35] ,n1[3]);
    nor g5314(n5330 ,n3534 ,n5039);
    nand g5315(n3714 ,n830 ,n3195);
    nand g5316(n5549 ,n4818 ,n5366);
    nand g5317(n303 ,n206 ,n302);
    nand g5318(n3611 ,n1[40] ,n3043);
    not g5319(n2876 ,n2875);
    nand g5320(n1825 ,n807 ,n968);
    nor g5321(n6713 ,n6826 ,n6608);
    nand g5322(n3726 ,n1887 ,n3178);
    nor g5323(n2229 ,n1957 ,n1599);
    nor g5324(n2341 ,n1[47] ,n719);
    xnor g5325(n5582 ,n4660 ,n5262);
    or g5326(n2053 ,n951 ,n2028);
    nand g5327(n10[26] ,n4620 ,n5323);
    or g5328(n9[55] ,n4511 ,n5611);
    nand g5329(n3568 ,n1953 ,n2956);
    nand g5330(n10[4] ,n4616 ,n5316);
    or g5331(n166 ,n0[36] ,n1[36]);
    xnor g5332(n1342 ,n0[84] ,n7112);
    nand g5333(n1993 ,n1238 ,n1094);
    nand g5334(n3225 ,n1120 ,n2198);
    nand g5335(n5000 ,n1102 ,n4676);
    nand g5336(n5227 ,n5101 ,n5058);
    nor g5337(n2323 ,n724 ,n1746);
    nor g5338(n6293 ,n6234 ,n6200);
    nor g5339(n4754 ,n3501 ,n4417);
    nand g5340(n1996 ,n1076 ,n1212);
    nor g5341(n2453 ,n856 ,n1960);
    nor g5342(n5308 ,n5182 ,n5108);
    not g5343(n811 ,n0[2]);
    or g5344(n488 ,n0[99] ,n6956);
    nor g5345(n4527 ,n791 ,n4361);
    nand g5346(n6658 ,n0[117] ,n0[85]);
    nor g5347(n3013 ,n877 ,n2489);
    nand g5348(n9[77] ,n6026 ,n5968);
    nand g5349(n3423 ,n1953 ,n2930);
    xnor g5350(n237 ,n1[33] ,n0[33]);
    nand g5351(n587 ,n506 ,n586);
    nand g5352(n6624 ,n0[89] ,n6579);
    nor g5353(n2070 ,n1959 ,n1945);
    not g5354(n5940 ,n5939);
    nand g5355(n997 ,n0[68] ,n715);
    or g5356(n5477 ,n4704 ,n5328);
    xnor g5357(n1389 ,n1[80] ,n2[16]);
    xnor g5358(n407 ,n7005 ,n7037);
    nand g5359(n5168 ,n4237 ,n4857);
    nand g5360(n9[46] ,n3882 ,n5811);
    xnor g5361(n1685 ,n0[43] ,n0[27]);
    or g5362(n4215 ,n794 ,n3818);
    xnor g5363(n1263 ,n0[87] ,n7115);
    nor g5364(n2974 ,n2620 ,n2370);
    xnor g5365(n6931 ,n78 ,n151);
    nor g5366(n4978 ,n3529 ,n4611);
    nand g5367(n362 ,n7022 ,n6990);
    xnor g5368(n400 ,n6998 ,n7030);
    nor g5369(n5932 ,n4653 ,n5772);
    xnor g5370(n1258 ,n1[47] ,n4[7]);
    nor g5371(n4811 ,n4377 ,n4409);
    nand g5372(n5834 ,n4280 ,n5719);
    nor g5373(n2203 ,n1961 ,n1937);
    or g5374(n4737 ,n3526 ,n4550);
    xnor g5375(n1593 ,n0[96] ,n1[96]);
    nor g5376(n901 ,n1[4] ,n2[4]);
    xnor g5377(n6929 ,n382 ,n455);
    nor g5378(n2740 ,n1[33] ,n2593);
    nand g5379(n4507 ,n3619 ,n4276);
    nor g5380(n3474 ,n2303 ,n3031);
    nor g5381(n6165 ,n6099 ,n6084);
    nor g5382(n3441 ,n1954 ,n2955);
    nand g5383(n646 ,n0[66] ,n622);
    nand g5384(n3159 ,n2003 ,n2326);
    xor g5385(n6416 ,n6305 ,n6188);
    nand g5386(n2541 ,n1199 ,n1839);
    nand g5387(n6273 ,n6224 ,n6196);
    xnor g5388(n1617 ,n0[107] ,n1[107]);
    nor g5389(n2343 ,n0[85] ,n1956);
    xnor g5390(n5435 ,n4578 ,n5061);
    not g5391(n783 ,n7091);
    or g5392(n4138 ,n1960 ,n3849);
    nand g5393(n6317 ,n6301 ,n6303);
    xnor g5394(n1382 ,n6890 ,n6888);
    nand g5395(n3694 ,n1015 ,n3197);
    nor g5396(n5660 ,n4061 ,n5441);
    xnor g5397(n1621 ,n0[74] ,n1[74]);
    nor g5398(n2093 ,n1107 ,n1740);
    nand g5399(n5395 ,n5212 ,n5218);
    xnor g5400(n6864 ,n549 ,n575);
    nand g5401(n6577 ,n5125 ,n6575);
    nand g5402(n3757 ,n6806 ,n3064);
    nor g5403(n5810 ,n5558 ,n5619);
    xnor g5404(n6219 ,n5769 ,n6109);
    nand g5405(n9[66] ,n5023 ,n6132);
    xnor g5406(n1849 ,n0[19] ,n0[18]);
    nand g5407(n919 ,n0[81] ,n741);
    nand g5408(n7007 ,n6657 ,n7166);
    not g5409(n721 ,n1964);
    nor g5410(n2235 ,n1918 ,n1838);
    not g5411(n2929 ,n2928);
    nand g5412(n419 ,n364 ,n418);
    nand g5413(n4312 ,n3021 ,n3906);
    xnor g5414(n1561 ,n1[39] ,n1[7]);
    nand g5415(n4111 ,n2459 ,n3479);
    xor g5416(n705 ,n2658 ,n6414);
    nor g5417(n3719 ,n1954 ,n2953);
    xnor g5418(n4897 ,n2809 ,n4455);
    xnor g5419(n5747 ,n5458 ,n2652);
    nor g5420(n2423 ,n721 ,n1507);
    nand g5421(n1123 ,n6893 ,n796);
    nor g5422(n6308 ,n5115 ,n6194);
    xnor g5423(n1522 ,n0[81] ,n4[25]);
    nand g5424(n5387 ,n4819 ,n5161);
    nand g5425(n3214 ,n1135 ,n2113);
    nand g5426(n6093 ,n3325 ,n5954);
    nand g5427(n6284 ,n6004 ,n6208);
    xnor g5428(n4899 ,n2854 ,n4468);
    nor g5429(n1777 ,n0[69] ,n967);
    nor g5430(n5424 ,n1954 ,n690);
    nand g5431(n55 ,n7061 ,n0[5]);
    nor g5432(n3438 ,n1222 ,n2816);
    xnor g5433(n5391 ,n5154 ,n1542);
    nand g5434(n1038 ,n0[73] ,n810);
    nand g5435(n615 ,n500 ,n614);
    or g5436(n3326 ,n1954 ,n2877);
    or g5437(n4743 ,n3515 ,n4537);
    nand g5438(n596 ,n469 ,n595);
    nor g5439(n6188 ,n5398 ,n6144);
    nor g5440(n4413 ,n3498 ,n4334);
    nand g5441(n3991 ,n0[101] ,n3490);
    nand g5442(n5003 ,n2512 ,n4674);
    nor g5443(n3844 ,n3582 ,n2727);
    xnor g5444(n249 ,n1[45] ,n0[45]);
    nand g5445(n6959 ,n6763 ,n6795);
    nand g5446(n350 ,n7040 ,n7008);
    nand g5447(n422 ,n337 ,n421);
    nand g5448(n3583 ,n0[111] ,n2794);
    xnor g5449(n1270 ,n0[42] ,n1[58]);
    nor g5450(n6556 ,n5826 ,n6522);
    nand g5451(n7010 ,n6643 ,n7163);
    or g5452(n9[100] ,n5664 ,n6102);
    nor g5453(n4857 ,n3409 ,n4711);
    xnor g5454(n1478 ,n1[46] ,n2[46]);
    nor g5455(n3442 ,n6 ,n3248);
    nand g5456(n1065 ,n0[127] ,n710);
    nor g5457(n1884 ,n823 ,n929);
    nor g5458(n2071 ,n719 ,n1525);
    nor g5459(n3109 ,n1877 ,n2221);
    nor g5460(n3502 ,n1222 ,n2835);
    or g5461(n3889 ,n2180 ,n3421);
    xnor g5462(n5291 ,n4210 ,n4991);
    nand g5463(n5823 ,n2742 ,n5661);
    nand g5464(n118 ,n33 ,n117);
    nand g5465(n216 ,n0[51] ,n1[51]);
    nor g5466(n6174 ,n5116 ,n6069);
    xnor g5467(n2685 ,n1[117] ,n1535);
    or g5468(n478 ,n0[111] ,n6968);
    xnor g5469(n5279 ,n4988 ,n4662);
    nor g5470(n4045 ,n2546 ,n3360);
    not g5471(n2868 ,n2867);
    nor g5472(n2252 ,n1959 ,n1387);
    nor g5473(n5599 ,n712 ,n5435);
    nor g5474(n2392 ,n721 ,n1540);
    xnor g5475(n1410 ,n1[93] ,n2[29]);
    nand g5476(n6553 ,n5092 ,n6534);
    nand g5477(n6444 ,n6359 ,n6304);
    nand g5478(n4484 ,n4289 ,n4035);
    or g5479(n2079 ,n1962 ,n1931);
    or g5480(n6269 ,n712 ,n6243);
    nand g5481(n7006 ,n6644 ,n7167);
    nand g5482(n4237 ,n1966 ,n3947);
    nand g5483(n4226 ,n3858 ,n3926);
    xnor g5484(n6847 ,n88 ,n109);
    xnor g5485(n5782 ,n5270 ,n5461);
    not g5486(n5993 ,n5992);
    xor g5487(n688 ,n3947 ,n2847);
    nor g5488(n6440 ,n5163 ,n6357);
    nand g5489(n4078 ,n714 ,n3694);
    nand g5490(n207 ,n0[37] ,n1[37]);
    nor g5491(n3024 ,n2282 ,n2281);
    nand g5492(n162 ,n25 ,n161);
    nand g5493(n9[23] ,n5741 ,n6009);
    nor g5494(n2091 ,n1962 ,n1469);
    nand g5495(n7063 ,n655 ,n623);
    not g5496(n804 ,n0[0]);
    xnor g5497(n1357 ,n0[68] ,n0[52]);
    nand g5498(n4644 ,n3521 ,n4540);
    or g5499(n491 ,n0[103] ,n6960);
    nand g5500(n2586 ,n0[16] ,n1964);
    or g5501(n2102 ,n1962 ,n1470);
    nand g5502(n6649 ,n0[114] ,n0[82]);
    xnor g5503(n1589 ,n0[78] ,n1[78]);
    xnor g5504(n1672 ,n0[94] ,n4[22]);
    xnor g5505(n6856 ,n547 ,n571);
    nor g5506(n931 ,n746 ,n0[112]);
    xor g5507(n3822 ,n2681 ,n1[69]);
    nand g5508(n1201 ,n6836 ,n795);
    not g5509(n797 ,n6826);
    nand g5510(n3539 ,n6 ,n2793);
    nand g5511(n4064 ,n3664 ,n3503);
    xnor g5512(n1873 ,n0[17] ,n0[16]);
    nor g5513(n5329 ,n4147 ,n5029);
    nor g5514(n4552 ,n1166 ,n4246);
    nand g5515(n312 ,n181 ,n311);
    nor g5516(n5739 ,n1954 ,n5577);
    nand g5517(n5710 ,n3606 ,n5425);
    nand g5518(n4116 ,n3185 ,n3804);
    nand g5519(n6668 ,n0[95] ,n6580);
    nor g5520(n1739 ,n1049 ,n902);
    nand g5521(n6127 ,n717 ,n6106);
    nand g5522(n4938 ,n3394 ,n4723);
    nand g5523(n4986 ,n1190 ,n4787);
    xnor g5524(n4464 ,n3948 ,n2823);
    xnor g5525(n6937 ,n384 ,n459);
    nand g5526(n5094 ,n4244 ,n4958);
    xnor g5527(n533 ,n6977 ,n0[120]);
    or g5528(n2182 ,n1962 ,n1480);
    nand g5529(n3070 ,n1571 ,n2622);
    nand g5530(n597 ,n520 ,n596);
    nor g5531(n3476 ,n1954 ,n2946);
    nand g5532(n680 ,n1[18] ,n621);
    xnor g5533(n5078 ,n4668 ,n4425);
    xnor g5534(n5991 ,n5268 ,n5834);
    nor g5535(n3648 ,n1880 ,n3050);
    nor g5536(n6039 ,n1954 ,n5960);
    nand g5537(n2640 ,n773 ,n1964);
    nor g5538(n5074 ,n2737 ,n4968);
    not g5539(n6248 ,n6247);
    nand g5540(n1829 ,n0[72] ,n895);
    xnor g5541(n1935 ,n1[61] ,n2[61]);
    nand g5542(n3888 ,n708 ,n3511);
    nand g5543(n2172 ,n1016 ,n2015);
    nand g5544(n3376 ,n1953 ,n2913);
    nand g5545(n526 ,n0[106] ,n6963);
    nor g5546(n3964 ,n2406 ,n3716);
    nor g5547(n4169 ,n3723 ,n3933);
    xnor g5548(n4446 ,n2813 ,n3959);
    xnor g5549(n2805 ,n0[109] ,n1318);
    nand g5550(n460 ,n321 ,n459);
    nand g5551(n7157 ,n6581 ,n7122);
    xnor g5552(n1696 ,n6939 ,n6936);
    nand g5553(n1096 ,n0[61] ,n788);
    xnor g5554(n6940 ,n537 ,n613);
    nor g5555(n3088 ,n1221 ,n2359);
    xnor g5556(n1387 ,n1[36] ,n2[36]);
    not g5557(n5778 ,n5777);
    nor g5558(n5181 ,n6824 ,n4902);
    nand g5559(n1039 ,n6825 ,n6824);
    nand g5560(n5327 ,n790 ,n5173);
    nor g5561(n2242 ,n721 ,n1519);
    nand g5562(n9[29] ,n5400 ,n5909);
    nand g5563(n9[115] ,n4421 ,n6540);
    nand g5564(n6278 ,n6235 ,n6218);
    nand g5565(n5831 ,n4321 ,n5643);
    nand g5566(n3322 ,n1953 ,n2877);
    nand g5567(n5421 ,n4948 ,n5280);
    nor g5568(n6192 ,n792 ,n6131);
    nor g5569(n3068 ,n1813 ,n2423);
    xnor g5570(n6949 ,n387 ,n465);
    nor g5571(n2758 ,n1495 ,n2636);
    nand g5572(n5145 ,n6827 ,n4915);
    nor g5573(n5649 ,n6 ,n5528);
    nor g5574(n903 ,n800 ,n0[120]);
    xnor g5575(n1703 ,n6843 ,n6841);
    nand g5576(n1141 ,n6892 ,n796);
    or g5577(n4074 ,n710 ,n3797);
    nand g5578(n5939 ,n4393 ,n5773);
    not g5579(n829 ,n0[110]);
    nor g5580(n2120 ,n6 ,n1975);
    xnor g5581(n1367 ,n7094 ,n7052);
    nor g5582(n3795 ,n2488 ,n3188);
    xnor g5583(n1465 ,n1[92] ,n2[28]);
    nor g5584(n3361 ,n1[93] ,n2959);
    or g5585(n23 ,n7069 ,n0[13]);
    nor g5586(n3096 ,n975 ,n2643);
    nand g5587(n2546 ,n1159 ,n1807);
    nand g5588(n3202 ,n1112 ,n2119);
    nand g5589(n7086 ,n679 ,n636);
    nand g5590(n2568 ,n1[33] ,n707);
    nor g5591(n5030 ,n2325 ,n5005);
    nand g5592(n569 ,n511 ,n568);
    xnor g5593(n2696 ,n1[113] ,n1533);
    nor g5594(n3566 ,n1954 ,n2956);
    nand g5595(n6067 ,n4848 ,n5978);
    nand g5596(n2576 ,n714 ,n2023);
    nor g5597(n4189 ,n3750 ,n3988);
    nand g5598(n3156 ,n2006 ,n2326);
    xnor g5599(n88 ,n0[4] ,n7060);
    nor g5600(n2302 ,n1959 ,n1390);
    nor g5601(n6061 ,n5700 ,n5963);
    nor g5602(n5407 ,n711 ,n5267);
    nor g5603(n5409 ,n706 ,n5215);
    nand g5604(n6503 ,n6382 ,n6415);
    xnor g5605(n5464 ,n4578 ,n5060);
    nand g5606(n7146 ,n6622 ,n6706);
    nand g5607(n6805 ,n6581 ,n7109);
    nand g5608(n6963 ,n6740 ,n6785);
    nand g5609(n3970 ,n3583 ,n3113);
    nor g5610(n888 ,n728 ,n0[80]);
    or g5611(n4141 ,n1959 ,n3816);
    nor g5612(n5234 ,n3488 ,n5166);
    nand g5613(n1860 ,n0[23] ,n1221);
    nor g5614(n2285 ,n6 ,n1763);
    not g5615(n729 ,n0[8]);
    or g5616(n2048 ,n1962 ,n1938);
    nand g5617(n599 ,n521 ,n598);
    nor g5618(n4162 ,n6 ,n4103);
    nand g5619(n6981 ,n6767 ,n6791);
    nand g5620(n2349 ,n774 ,n718);
    nor g5621(n2319 ,n1957 ,n1593);
    nor g5622(n5690 ,n5559 ,n5434);
    nor g5623(n2244 ,n1961 ,n1422);
    xnor g5624(n1520 ,n0[13] ,n1[13]);
    not g5625(n3945 ,n3944);
    nor g5626(n5359 ,n3526 ,n5140);
    nand g5627(n6746 ,n0[56] ,n6737);
    nand g5628(n1136 ,n6939 ,n795);
    xnor g5629(n1311 ,n1[63] ,n1[31]);
    nor g5630(n3525 ,n2177 ,n2976);
    nand g5631(n6465 ,n6401 ,n6423);
    nor g5632(n5044 ,n791 ,n4929);
    nand g5633(n6767 ,n0[60] ,n6737);
    nand g5634(n6968 ,n6749 ,n6779);
    nor g5635(n2460 ,n956 ,n1805);
    nor g5636(n2065 ,n721 ,n1489);
    nand g5637(n144 ,n30 ,n143);
    nor g5638(n3592 ,n765 ,n3044);
    or g5639(n9[103] ,n5668 ,n6239);
    nand g5640(n3990 ,n0[4] ,n3491);
    nor g5641(n1048 ,n0[57] ,n0[56]);
    nor g5642(n3515 ,n6825 ,n2807);
    xnor g5643(n1467 ,n1[41] ,n2[41]);
    nand g5644(n4303 ,n2771 ,n3860);
    xnor g5645(n6840 ,n543 ,n563);
    xor g5646(n6033 ,n5931 ,n2702);
    xnor g5647(n2911 ,n1678 ,n1510);
    nand g5648(n2396 ,n1964 ,n1499);
    xnor g5649(n3832 ,n1[81] ,n2696);
    nand g5650(n3541 ,n6 ,n2718);
    xnor g5651(n6415 ,n6307 ,n6143);
    nor g5652(n3803 ,n2143 ,n3069);
    nand g5653(n4536 ,n1119 ,n4127);
    or g5654(n2068 ,n1962 ,n1944);
    nand g5655(n4542 ,n1167 ,n4138);
    nor g5656(n3605 ,n764 ,n2797);
    nand g5657(n5838 ,n4954 ,n5643);
    xnor g5658(n1347 ,n0[13] ,n4[29]);
    nand g5659(n1144 ,n6859 ,n797);
    nand g5660(n4777 ,n1955 ,n4571);
    xnor g5661(n92 ,n0[8] ,n7064);
    nand g5662(n4322 ,n3647 ,n3856);
    not g5663(n774 ,n1[57]);
    xnor g5664(n1550 ,n1[34] ,n1[2]);
    nand g5665(n971 ,n0[88] ,n723);
    xor g5666(n7112 ,n0[52] ,n0[20]);
    or g5667(n5820 ,n4315 ,n5628);
    xnor g5668(n1471 ,n1[74] ,n2[10]);
    or g5669(n335 ,n7027 ,n6995);
    not g5670(n1529 ,n1528);
    xnor g5671(n1926 ,n1[30] ,n2[30]);
    or g5672(n3807 ,n6825 ,n2819);
    nand g5673(n4796 ,n3593 ,n4392);
    nand g5674(n3728 ,n7128 ,n3107);
    xnor g5675(n1692 ,n6914 ,n6915);
    nand g5676(n1016 ,n806 ,n728);
    nand g5677(n5796 ,n5625 ,n5617);
    nand g5678(n5813 ,n3596 ,n5621);
    nand g5679(n1062 ,n0[36] ,n710);
    nor g5680(n5602 ,n4686 ,n5454);
    nand g5681(n6969 ,n6751 ,n6781);
    nand g5682(n1164 ,n6923 ,n796);
    xnor g5683(n1668 ,n0[108] ,n4[4]);
    or g5684(n4738 ,n3527 ,n4556);
    nor g5685(n2275 ,n1957 ,n1635);
    nand g5686(n5759 ,n5423 ,n5603);
    xor g5687(n4904 ,n4457 ,n2851);
    nand g5688(n4568 ,n2526 ,n4215);
    nand g5689(n126 ,n36 ,n125);
    nor g5690(n5491 ,n3465 ,n5241);
    nor g5691(n914 ,n0[71] ,n788);
    nand g5692(n6660 ,n1[85] ,n6579);
    xnor g5693(n6922 ,n228 ,n299);
    nand g5694(n6700 ,n0[81] ,n6579);
    nand g5695(n2755 ,n1577 ,n2633);
    xnor g5696(n1640 ,n0[22] ,n1[22]);
    nand g5697(n3150 ,n1[116] ,n2360);
    nand g5698(n9[105] ,n4975 ,n6395);
    not g5699(n2870 ,n2869);
    or g5700(n2156 ,n1959 ,n1471);
    nand g5701(n9[7] ,n5654 ,n5824);
    xnor g5702(n3814 ,n2651 ,n2711);
    nand g5703(n9[64] ,n5307 ,n6525);
    nand g5704(n458 ,n345 ,n457);
    nor g5705(n6144 ,n793 ,n6044);
    nor g5706(n6070 ,n792 ,n5970);
    nand g5707(n6680 ,n0[122] ,n0[90]);
    nor g5708(n3617 ,n774 ,n2994);
    nor g5709(n3893 ,n2197 ,n3742);
    nand g5710(n3216 ,n1180 ,n2152);
    nor g5711(n2225 ,n1959 ,n1415);
    nor g5712(n4009 ,n3217 ,n3613);
    xnor g5713(n2718 ,n1724 ,n1570);
    nor g5714(n4441 ,n3881 ,n4144);
    nand g5715(n4309 ,n7134 ,n3920);
    nand g5716(n3163 ,n714 ,n2503);
    xnor g5717(n4842 ,n0[14] ,n4571);
    or g5718(n2747 ,n2147 ,n2059);
    xnor g5719(n2716 ,n1722 ,n1564);
    nand g5720(n4981 ,n3312 ,n4720);
    nor g5721(n3256 ,n0[72] ,n2405);
    nand g5722(n4980 ,n3320 ,n4721);
    nand g5723(n3995 ,n0[103] ,n3490);
    nor g5724(n5506 ,n5304 ,n5293);
    nand g5725(n7136 ,n6652 ,n6716);
    nand g5726(n6010 ,n3301 ,n5857);
    nand g5727(n3232 ,n1209 ,n2101);
    nand g5728(n159 ,n44 ,n158);
    nand g5729(n1151 ,n6853 ,n795);
    nand g5730(n5884 ,n5096 ,n5754);
    nand g5731(n2965 ,n2522 ,n2307);
    nand g5732(n6651 ,n0[90] ,n6580);
    nor g5733(n2015 ,n741 ,n984);
    nand g5734(n4072 ,n3306 ,n3682);
    or g5735(n473 ,n0[123] ,n6980);
    or g5736(n5633 ,n3453 ,n5476);
    nor g5737(n5673 ,n2325 ,n5529);
    nand g5738(n280 ,n175 ,n279);
    nand g5739(n57 ,n7058 ,n0[2]);
    not g5740(n777 ,n0[87]);
    xnor g5741(n6841 ,n391 ,n411);
    xnor g5742(n6917 ,n379 ,n449);
    nand g5743(n5968 ,n1953 ,n5849);
    not g5744(n6218 ,n6217);
    xnor g5745(n1378 ,n6897 ,n6896);
    nand g5746(n3674 ,n0[12] ,n3082);
    nand g5747(n3799 ,n2535 ,n3057);
    nand g5748(n3226 ,n1184 ,n2201);
    nand g5749(n6632 ,n1[70] ,n6579);
    xnor g5750(n4473 ,n2798 ,n3938);
    or g5751(n2140 ,n1045 ,n1892);
    nor g5752(n882 ,n0[117] ,n6);
    nand g5753(n4643 ,n794 ,n4461);
    or g5754(n4750 ,n3512 ,n4543);
    xnor g5755(n1461 ,n0[85] ,n0[69]);
    nor g5756(n1017 ,n751 ,n0[42]);
    not g5757(n1025 ,n1024);
    xnor g5758(n3951 ,n2832 ,n2850);
    not g5759(n828 ,n1[60]);
    not g5760(n5108 ,n5020);
    nand g5761(n3977 ,n0[111] ,n3490);
    not g5762(n790 ,n708);
    or g5763(n5543 ,n3462 ,n5384);
    nand g5764(n7049 ,n6692 ,n7124);
    not g5765(n5172 ,n5171);
    nand g5766(n6290 ,n3309 ,n6177);
    nand g5767(n2022 ,n1000 ,n1047);
    nor g5768(n1168 ,n785 ,n716);
    nor g5769(n4295 ,n3620 ,n3994);
    nand g5770(n664 ,n1[22] ,n621);
    nand g5771(n3161 ,n1969 ,n2326);
    nor g5772(n5987 ,n713 ,n5934);
    not g5773(n6209 ,n6208);
    nand g5774(n6500 ,n5982 ,n6433);
    or g5775(n17 ,n7083 ,n0[27]);
    nor g5776(n1246 ,n823 ,n725);
    xnor g5777(n1678 ,n0[39] ,n1[55]);
    nand g5778(n463 ,n348 ,n462);
    nor g5779(n2247 ,n1962 ,n1428);
    xnor g5780(n1490 ,n0[8] ,n1[8]);
    nand g5781(n917 ,n0[74] ,n724);
    nor g5782(n5494 ,n6 ,n5377);
    nor g5783(n2002 ,n864 ,n926);
    nor g5784(n4263 ,n1962 ,n3825);
    nand g5785(n4270 ,n2075 ,n3966);
    nand g5786(n6161 ,n3349 ,n6049);
    nand g5787(n4584 ,n4063 ,n4275);
    nand g5788(n4985 ,n1177 ,n4765);
    nand g5789(n3260 ,n2011 ,n2265);
    nor g5790(n5417 ,n711 ,n5228);
    nor g5791(n3953 ,n3563 ,n3432);
    or g5792(n176 ,n0[57] ,n1[57]);
    not g5793(n753 ,n0[126]);
    not g5794(n4581 ,n4582);
    xnor g5795(n4671 ,n4245 ,n1983);
    xnor g5796(n5262 ,n5001 ,n5008);
    not g5797(n5266 ,n5265);
    nor g5798(n2773 ,n888 ,n2595);
    nand g5799(n2006 ,n1059 ,n883);
    nand g5800(n5918 ,n4521 ,n5808);
    xnor g5801(n1705 ,n0[69] ,n1[85]);
    nand g5802(n1116 ,n6935 ,n796);
    nor g5803(n4490 ,n4165 ,n4352);
    nand g5804(n4323 ,n2597 ,n3859);
    nand g5805(n5121 ,n798 ,n4915);
    or g5806(n3372 ,n1954 ,n2911);
    nor g5807(n5005 ,n4260 ,n4648);
    nand g5808(n6457 ,n3548 ,n6347);
    nand g5809(n4504 ,n1039 ,n4119);
    or g5810(n1015 ,n750 ,n0[10]);
    xnor g5811(n1606 ,n0[70] ,n1[70]);
    nor g5812(n4194 ,n6 ,n4106);
    or g5813(n3111 ,n748 ,n2215);
    nor g5814(n5488 ,n5382 ,n5308);
    or g5815(n3338 ,n1954 ,n2894);
    nor g5816(n2422 ,n791 ,n1587);
    or g5817(n9[95] ,n5257 ,n6017);
    nand g5818(n513 ,n0[98] ,n6955);
    nand g5819(n6455 ,n3351 ,n6362);
    nand g5820(n1240 ,n3[2] ,n3[1]);
    xnor g5821(n2883 ,n1298 ,n1361);
    nand g5822(n5926 ,n4480 ,n5800);
    nor g5823(n5764 ,n5101 ,n5633);
    nand g5824(n3651 ,n0[18] ,n3093);
    nand g5825(n64 ,n7075 ,n0[19]);
    nand g5826(n3755 ,n7144 ,n3063);
    nor g5827(n4746 ,n3806 ,n4567);
    xor g5828(n7102 ,n0[42] ,n0[10]);
    nor g5829(n2162 ,n1963 ,n1563);
    xnor g5830(n1688 ,n6934 ,n6935);
    nor g5831(n4033 ,n3768 ,n2754);
    xnor g5832(n2956 ,n1705 ,n1547);
    nor g5833(n4561 ,n1178 ,n4249);
    nor g5834(n996 ,n0[59] ,n0[56]);
    nand g5835(n3753 ,n7146 ,n3054);
    nand g5836(n4073 ,n3357 ,n3685);
    nand g5837(n3230 ,n7164 ,n2562);
    nand g5838(n498 ,n0[117] ,n6974);
    nand g5839(n6533 ,n6483 ,n6500);
    nor g5840(n2792 ,n1499 ,n2604);
    xnor g5841(n4926 ,n2844 ,n4464);
    or g5842(n3430 ,n788 ,n3260);
    or g5843(n5499 ,n4688 ,n5354);
    nand g5844(n3164 ,n1971 ,n2326);
    nor g5845(n3054 ,n1801 ,n2273);
    nor g5846(n1178 ,n846 ,n716);
    nand g5847(n682 ,n1[0] ,n621);
    nand g5848(n3037 ,n1005 ,n2476);
    nand g5849(n2528 ,n984 ,n1905);
    nor g5850(n6456 ,n6371 ,n6282);
    nor g5851(n3916 ,n2317 ,n3759);
    xnor g5852(n2704 ,n0[114] ,n1519);
    nand g5853(n7024 ,n6632 ,n7149);
    nand g5854(n6382 ,n3569 ,n6269);
    nor g5855(n5283 ,n4624 ,n5071);
    nand g5856(n2021 ,n714 ,n1035);
    nand g5857(n9[78] ,n4340 ,n5799);
    nand g5858(n2632 ,n799 ,n1964);
    nand g5859(n1835 ,n752 ,n1048);
    nand g5860(n147 ,n46 ,n146);
    nand g5861(n6697 ,n0[67] ,n6580);
    or g5862(n3355 ,n1954 ,n2902);
    xnor g5863(n1537 ,n0[28] ,n1[28]);
    nor g5864(n6305 ,n4931 ,n6192);
    xnor g5865(n1386 ,n1[33] ,n2[33]);
    nor g5866(n2256 ,n1957 ,n1633);
    xnor g5867(n1936 ,n1[90] ,n2[26]);
    xnor g5868(n2655 ,n1[126] ,n1355);
    nand g5869(n5923 ,n3967 ,n5746);
    nand g5870(n4771 ,n2560 ,n4436);
    nand g5871(n4331 ,n0[61] ,n3898);
    nand g5872(n1115 ,n6952 ,n796);
    nand g5873(n5216 ,n5036 ,n5035);
    nor g5874(n6253 ,n6023 ,n6213);
    nor g5875(n3211 ,n1189 ,n2096);
    xor g5876(n694 ,n5260 ,n1547);
    or g5877(n332 ,n7020 ,n6988);
    nand g5878(n616 ,n485 ,n615);
    nand g5879(n1064 ,n0[28] ,n791);
    xnor g5880(n1359 ,n0[47] ,n0[31]);
    xnor g5881(n2855 ,n1335 ,n1525);
    nand g5882(n4291 ,n4000 ,n3927);
    nand g5883(n160 ,n29 ,n159);
    nor g5884(n2143 ,n886 ,n1766);
    nand g5885(n9[57] ,n5705 ,n6552);
    nand g5886(n7066 ,n660 ,n629);
    or g5887(n4415 ,n4351 ,n4089);
    nand g5888(n5931 ,n4423 ,n5775);
    not g5889(n4998 ,n4997);
    xnor g5890(n2930 ,n1672 ,n1586);
    xnor g5891(n1716 ,n0[41] ,n1[57]);
    not g5892(n758 ,n0[33]);
    nand g5893(n520 ,n0[115] ,n6972);
    xnor g5894(n6895 ,n100 ,n133);
    nor g5895(n4856 ,n3403 ,n4709);
    xnor g5896(n1588 ,n0[100] ,n1[100]);
    nand g5897(n3020 ,n1569 ,n2639);
    nand g5898(n6970 ,n6764 ,n6783);
    xnor g5899(n3810 ,n0[77] ,n2648);
    nand g5900(n10[8] ,n4768 ,n5345);
    nand g5901(n4535 ,n2326 ,n4218);
    nor g5902(n2317 ,n1962 ,n1419);
    xnor g5903(n6854 ,n242 ,n265);
    nand g5904(n613 ,n505 ,n612);
    xnor g5905(n4468 ,n2836 ,n3960);
    nor g5906(n3885 ,n2067 ,n3740);
    nand g5907(n3637 ,n1[53] ,n2983);
    or g5908(n28 ,n7058 ,n0[2]);
    or g5909(n4610 ,n2561 ,n4465);
    not g5910(n713 ,n717);
    xor g5911(n7095 ,n0[35] ,n0[3]);
    nand g5912(n5269 ,n4190 ,n5063);
    not g5913(n1036 ,n1035);
    nand g5914(n4582 ,n1098 ,n4229);
    nand g5915(n10[9] ,n4789 ,n5514);
    nand g5916(n1186 ,n6864 ,n796);
    or g5917(n4152 ,n2738 ,n4064);
    nand g5918(n6080 ,n5634 ,n5988);
    nand g5919(n3704 ,n2072 ,n3170);
    or g5920(n5652 ,n5188 ,n5432);
    nor g5921(n1742 ,n0[120] ,n1009);
    nand g5922(n3298 ,n1952 ,n2873);
    nor g5923(n4540 ,n1203 ,n4136);
    xnor g5924(n1530 ,n1[20] ,n782);
    nand g5925(n4784 ,n1138 ,n4504);
    nand g5926(n9[111] ,n5860 ,n6169);
    nor g5927(n5626 ,n1954 ,n5447);
    or g5928(n9[53] ,n4513 ,n5767);
    nand g5929(n288 ,n189 ,n287);
    nand g5930(n259 ,n209 ,n258);
    nand g5931(n652 ,n0[83] ,n622);
    xnor g5932(n536 ,n6980 ,n0[123]);
    nor g5933(n5047 ,n715 ,n4929);
    nor g5934(n3527 ,n6825 ,n2837);
    nor g5935(n3424 ,n1954 ,n2929);
    nand g5936(n583 ,n501 ,n582);
    nand g5937(n1000 ,n0[34] ,n758);
    xor g5938(n697 ,n1584 ,n5464);
    nor g5939(n6106 ,n3905 ,n5981);
    nor g5940(n2207 ,n721 ,n1537);
    nand g5941(n1897 ,n0[62] ,n1221);
    nor g5942(n938 ,n746 ,n0[113]);
    nor g5943(n6721 ,n6826 ,n6607);
    nand g5944(n5240 ,n5083 ,n5064);
    nor g5945(n1222 ,n726 ,n845);
    nand g5946(n500 ,n0[124] ,n6981);
    xnor g5947(n1632 ,n0[93] ,n1[93]);
    nand g5948(n6491 ,n6459 ,n6455);
    nor g5949(n5021 ,n711 ,n4876);
    xnor g5950(n3841 ,n2700 ,n1975);
    not g5951(n622 ,n6826);
    nand g5952(n2616 ,n735 ,n1964);
    xnor g5953(n1612 ,n0[124] ,n1[124]);
    or g5954(n6371 ,n3321 ,n6260);
    nand g5955(n1834 ,n0[27] ,n1221);
    nand g5956(n984 ,n0[80] ,n714);
    nand g5957(n137 ,n48 ,n136);
    xnor g5958(n2830 ,n0[102] ,n1278);
    nand g5959(n1907 ,n0[65] ,n990);
    not g5960(n1555 ,n1554);
    nand g5961(n1887 ,n0[127] ,n1221);
    nand g5962(n6750 ,n0[57] ,n6737);
    or g5963(n6180 ,n711 ,n6141);
    nand g5964(n446 ,n320 ,n445);
    nor g5965(n3329 ,n1954 ,n2891);
    nand g5966(n1882 ,n0[20] ,n966);
    not g5967(n5844 ,n5845);
    xnor g5968(n1426 ,n1[21] ,n2[21]);
    nand g5969(n9[117] ,n5765 ,n6022);
    xor g5970(n704 ,n6413 ,n2671);
    nor g5971(n4672 ,n793 ,n4408);
    or g5972(n5335 ,n4066 ,n5110);
    nor g5973(n3851 ,n2189 ,n3559);
    xnor g5974(n6933 ,n383 ,n457);
    nand g5975(n5743 ,n1953 ,n695);
    nor g5976(n3074 ,n1843 ,n2477);
    xnor g5977(n2942 ,n1590 ,n1505);
    nand g5978(n5161 ,n798 ,n4918);
    nor g5979(n5871 ,n711 ,n5836);
    or g5980(n9[9] ,n4798 ,n6441);
    xnor g5981(n6912 ,n530 ,n599);
    not g5982(n716 ,n797);
    not g5983(n964 ,n965);
    not g5984(n1034 ,n1033);
    nand g5985(n6288 ,n6232 ,n6212);
    nor g5986(n4429 ,n2263 ,n4228);
    nand g5987(n5374 ,n3574 ,n5063);
    xnor g5988(n6858 ,n243 ,n267);
    nand g5989(n7035 ,n6648 ,n7138);
    nand g5990(n3710 ,n841 ,n3184);
    nor g5991(n2273 ,n721 ,n1525);
    xnor g5992(n535 ,n6979 ,n0[122]);
    nand g5993(n6354 ,n5987 ,n6282);
    not g5994(n1513 ,n1512);
    xnor g5995(n1580 ,n0[57] ,n4[17]);
    nor g5996(n4173 ,n2545 ,n3935);
    or g5997(n9[40] ,n4482 ,n6560);
    nand g5998(n632 ,n0[86] ,n622);
    nor g5999(n4988 ,n2515 ,n4678);
    nor g6000(n6110 ,n5494 ,n5981);
    nor g6001(n6711 ,n6826 ,n6587);
    or g6002(n3363 ,n983 ,n3256);
    xnor g6003(n240 ,n1[36] ,n0[36]);
    xnor g6004(n2826 ,n0[104] ,n1376);
    nand g6005(n6759 ,n0[36] ,n6737);
    not g6006(n2947 ,n2946);
    nand g6007(n5377 ,n4069 ,n5027);
    nand g6008(n6810 ,n6581 ,n7104);
    nand g6009(n2389 ,n707 ,n1498);
    not g6010(n1003 ,n1002);
    nor g6011(n5402 ,n5105 ,n5264);
    xnor g6012(n1631 ,n0[95] ,n1[95]);
    not g6013(n748 ,n0[27]);
    nand g6014(n3194 ,n1970 ,n2326);
    nand g6015(n5681 ,n3455 ,n5476);
    or g6016(n4224 ,n792 ,n3838);
    nor g6017(n2329 ,n1783 ,n2022);
    xnor g6018(n1558 ,n0[21] ,n1[21]);
    nand g6019(n1979 ,n879 ,n1088);
    nand g6020(n53 ,n7071 ,n0[15]);
    nand g6021(n3186 ,n728 ,n2528);
    or g6022(n2088 ,n1961 ,n1446);
    nand g6023(n3538 ,n6 ,n2716);
    nand g6024(n203 ,n0[33] ,n1[33]);
    or g6025(n331 ,n7023 ,n6991);
    nor g6026(n5230 ,n3337 ,n5089);
    nand g6027(n4950 ,n2769 ,n4815);
    nor g6028(n1864 ,n822 ,n995);
    or g6029(n27 ,n7061 ,n0[5]);
    nand g6030(n3463 ,n1953 ,n2939);
    nand g6031(n6359 ,n5780 ,n6283);
    xnor g6032(n6250 ,n6113 ,n1679);
    nand g6033(n5881 ,n1952 ,n5817);
    xnor g6034(n6206 ,n5833 ,n6105);
    nor g6035(n6544 ,n713 ,n6513);
    nand g6036(n3752 ,n7147 ,n3061);
    nor g6037(n2240 ,n719 ,n1618);
    not g6038(n1484 ,n1485);
    nand g6039(n1905 ,n0[82] ,n939);
    nand g6040(n3616 ,n1[56] ,n2992);
    xnor g6041(n7054 ,n236 ,n315);
    or g6042(n25 ,n7086 ,n0[30]);
    nor g6043(n4599 ,n4205 ,n4384);
    nand g6044(n309 ,n201 ,n308);
    nor g6045(n5512 ,n5315 ,n5336);
    or g6046(n6092 ,n5687 ,n5988);
    xnor g6047(n1396 ,n1[39] ,n2[39]);
    nand g6048(n5466 ,n3568 ,n5286);
    nor g6049(n5102 ,n713 ,n5000);
    xnor g6050(n1422 ,n1[9] ,n2[9]);
    nor g6051(n5600 ,n1954 ,n691);
    not g6052(n6194 ,n6193);
    nand g6053(n612 ,n473 ,n611);
    xnor g6054(n2817 ,n1319 ,n1670);
    nand g6055(n1156 ,n6921 ,n795);
    not g6056(n733 ,n0[90]);
    nor g6057(n1729 ,n0[0] ,n972);
    xnor g6058(n2804 ,n1375 ,n1658);
    nand g6059(n1876 ,n0[50] ,n1221);
    not g6060(n816 ,n0[5]);
    nand g6061(n6980 ,n6760 ,n6793);
    nand g6062(n6983 ,n6752 ,n6780);
    nand g6063(n296 ,n182 ,n295);
    nand g6064(n6736 ,n3[3] ,n6733);
    xnor g6065(n1275 ,n1[40] ,n4[0]);
    nor g6066(n2258 ,n1962 ,n1927);
    nor g6067(n4310 ,n2552 ,n3896);
    nor g6068(n2062 ,n907 ,n1960);
    or g6069(n2187 ,n1960 ,n1939);
    nand g6070(n9[90] ,n5648 ,n6163);
    nand g6071(n3175 ,n1979 ,n2326);
    nor g6072(n3485 ,n1954 ,n2951);
    xnor g6073(n101 ,n0[17] ,n7073);
    nor g6074(n4130 ,n710 ,n4113);
    nand g6075(n6053 ,n6001 ,n5777);
    xnor g6076(n4422 ,n3813 ,n1984);
    nand g6077(n4862 ,n3340 ,n4636);
    nand g6078(n3126 ,n1[35] ,n2616);
    nand g6079(n4550 ,n1124 ,n4265);
    xnor g6080(n6838 ,n238 ,n257);
    nor g6081(n3440 ,n1792 ,n2725);
    or g6082(n38 ,n7079 ,n0[23]);
    nand g6083(n3255 ,n922 ,n2053);
    nand g6084(n197 ,n0[44] ,n1[44]);
    nor g6085(n6542 ,n706 ,n6510);
    nand g6086(n562 ,n484 ,n561);
    nand g6087(n4515 ,n3670 ,n4202);
    nand g6088(n4245 ,n6 ,n3841);
    xnor g6089(n2844 ,n1280 ,n1338);
    nor g6090(n4627 ,n3746 ,n4380);
    not g6091(n4909 ,n4908);
    not g6092(n1577 ,n1576);
    nand g6093(n6096 ,n6021 ,n5781);
    xnor g6094(n4916 ,n2815 ,n4440);
    nor g6095(n3501 ,n1222 ,n2828);
    nor g6096(n3536 ,n6825 ,n2799);
    nor g6097(n5618 ,n711 ,n5430);
    xnor g6098(n1671 ,n6886 ,n6887);
    nand g6099(n2545 ,n1155 ,n1811);
    nand g6100(n3981 ,n0[30] ,n3490);
    nand g6101(n4500 ,n2326 ,n4360);
    or g6102(n5787 ,n5597 ,n5555);
    nand g6103(n9[112] ,n5827 ,n6504);
    nor g6104(n1858 ,n820 ,n1220);
    nand g6105(n5532 ,n4832 ,n5357);
    or g6106(n484 ,n0[98] ,n6955);
    nand g6107(n4327 ,n2593 ,n3937);
    nand g6108(n425 ,n370 ,n424);
    xnor g6109(n5994 ,n5836 ,n5841);
    nand g6110(n6447 ,n3307 ,n6325);
    nand g6111(n128 ,n23 ,n127);
    xnor g6112(n2682 ,n1668 ,n1612);
    xnor g6113(n394 ,n6992 ,n7024);
    nand g6114(n6765 ,n0[39] ,n6737);
    xnor g6115(n2953 ,n1652 ,n1516);
    xnor g6116(n1712 ,n6862 ,n6863);
    nand g6117(n6787 ,n1[98] ,n7088);
    nor g6118(n2409 ,n724 ,n1861);
    nor g6119(n5438 ,n3294 ,n5223);
    nand g6120(n4766 ,n2560 ,n4444);
    nor g6121(n5959 ,n711 ,n5937);
    nand g6122(n3792 ,n3191 ,n3187);
    xnor g6123(n6898 ,n253 ,n287);
    nor g6124(n5134 ,n727 ,n4896);
    nor g6125(n4387 ,n3205 ,n4272);
    xnor g6126(n75 ,n0[22] ,n7078);
    nor g6127(n4749 ,n6 ,n4447);
    xnor g6128(n1721 ,n6942 ,n6943);
    nor g6129(n173 ,n0[33] ,n1[33]);
    nand g6130(n6530 ,n6498 ,n6487);
    nand g6131(n3600 ,n0[39] ,n2794);
    nand g6132(n6971 ,n6755 ,n6770);
    or g6133(n5814 ,n4333 ,n5610);
    xnor g6134(n6191 ,n5831 ,n6112);
    xnor g6135(n4903 ,n4578 ,n4574);
    nand g6136(n9[83] ,n5242 ,n6545);
    nor g6137(n2768 ,n2092 ,n2091);
    nor g6138(n6407 ,n6240 ,n6320);
    xnor g6139(n2939 ,n1589 ,n1541);
    or g6140(n876 ,n724 ,n0[0]);
    nand g6141(n3144 ,n2607 ,n2461);
    nor g6142(n4665 ,n880 ,n4470);
    or g6143(n2057 ,n719 ,n1519);
    nor g6144(n2390 ,n0[42] ,n719);
    xnor g6145(n396 ,n6994 ,n7026);
    xnor g6146(n6074 ,n5938 ,n1345);
    nor g6147(n4021 ,n3206 ,n3396);
    or g6148(n2160 ,n1962 ,n1434);
    nand g6149(n4349 ,n2531 ,n3974);
    nand g6150(n4244 ,n1966 ,n3946);
    nand g6151(n7152 ,n6581 ,n7053);
    nand g6152(n141 ,n64 ,n140);
    nor g6153(n3608 ,n831 ,n2797);
    nor g6154(n3286 ,n1954 ,n2886);
    nor g6155(n900 ,n806 ,n0[82]);
    nor g6156(n2452 ,n817 ,n721);
    xnor g6157(n6120 ,n5942 ,n5948);
    nand g6158(n3770 ,n7127 ,n3001);
    nand g6159(n4637 ,n717 ,n4427);
    nand g6160(n5372 ,n3675 ,n5043);
    xnor g6161(n234 ,n1[61] ,n0[61]);
    nand g6162(n572 ,n491 ,n571);
    xnor g6163(n5852 ,n5567 ,n4677);
    nor g6164(n5414 ,n1954 ,n5219);
    nand g6165(n2480 ,n714 ,n1910);
    nand g6166(n6639 ,n0[66] ,n6579);
    nor g6167(n3961 ,n3425 ,n3454);
    not g6168(n808 ,n0[43]);
    nor g6169(n4316 ,n844 ,n3878);
    or g6170(n19 ,n7080 ,n0[24]);
    nand g6171(n4759 ,n3843 ,n4437);
    xnor g6172(n2647 ,n1989 ,n2000);
    nand g6173(n1968 ,n1096 ,n1061);
    nand g6174(n4047 ,n3629 ,n2063);
    nand g6175(n1180 ,n6863 ,n796);
    nor g6176(n4195 ,n6 ,n3957);
    xnor g6177(n1574 ,n1[41] ,n1[9]);
    xnor g6178(n99 ,n0[15] ,n7071);
    nor g6179(n1793 ,n728 ,n11);
    nor g6180(n6245 ,n5448 ,n6142);
    or g6181(n1857 ,n0[49] ,n979);
    xnor g6182(n6422 ,n6280 ,n6246);
    nor g6183(n5912 ,n5675 ,n5736);
    nand g6184(n6739 ,n0[54] ,n6737);
    xnor g6185(n5946 ,n5831 ,n1380);
    nand g6186(n2726 ,n937 ,n2428);
    xnor g6187(n1377 ,n0[89] ,n7117);
    or g6188(n2525 ,n6 ,n1972);
    nand g6189(n3748 ,n7153 ,n3072);
    nand g6190(n5765 ,n1953 ,n5593);
    nor g6191(n1026 ,n810 ,n0[74]);
    nor g6192(n5332 ,n3528 ,n5132);
    nand g6193(n6318 ,n6278 ,n6275);
    xnor g6194(n1582 ,n0[119] ,n0[103]);
    xnor g6195(n1291 ,n0[22] ,n0[6]);
    nor g6196(n4158 ,n3778 ,n4056);
    nor g6197(n6715 ,n6826 ,n6593);
    not g6198(n2592 ,n2591);
    nand g6199(n5483 ,n4706 ,n5301);
    nand g6200(n6546 ,n1952 ,n6514);
    xnor g6201(n1395 ,n1[40] ,n2[40]);
    nand g6202(n2606 ,n934 ,n1879);
    nor g6203(n5904 ,n706 ,n5831);
    nor g6204(n3416 ,n1222 ,n2844);
    or g6205(n5689 ,n5098 ,n5465);
    xnor g6206(n5277 ,n4670 ,n4992);
    nand g6207(n4795 ,n3983 ,n4437);
    nor g6208(n4989 ,n2502 ,n4675);
    nand g6209(n6758 ,n0[51] ,n6737);
    xnor g6210(n1726 ,n0[90] ,n4[18]);
    xnor g6211(n5475 ,n4210 ,n5156);
    nor g6212(n4384 ,n722 ,n4358);
    or g6213(n6086 ,n6015 ,n5991);
    nand g6214(n349 ,n7030 ,n6998);
    nor g6215(n1759 ,n0[17] ,n975);
    or g6216(n4722 ,n711 ,n4571);
    nand g6217(n298 ,n178 ,n297);
    nand g6218(n3679 ,n3147 ,n2170);
    nand g6219(n6182 ,n5544 ,n6122);
    xnor g6220(n2881 ,n1365 ,n1587);
    or g6221(n9[36] ,n4484 ,n5922);
    xnor g6222(n2691 ,n0[95] ,n1279);
    or g6223(n4615 ,n2561 ,n4466);
    nor g6224(n5049 ,n4713 ,n4880);
    xnor g6225(n98 ,n0[14] ,n7070);
    xnor g6226(n6843 ,n87 ,n107);
    nand g6227(n879 ,n0[23] ,n715);
    xnor g6228(n6985 ,n388 ,n467);
    nor g6229(n4029 ,n3696 ,n3274);
    nor g6230(n5302 ,n5084 ,n5053);
    nor g6231(n1813 ,n745 ,n11);
    not g6232(n5984 ,n5983);
    nand g6233(n3992 ,n0[38] ,n3490);
    nand g6234(n3182 ,n1978 ,n2326);
    nor g6235(n6129 ,n712 ,n6107);
    not g6236(n4689 ,n4688);
    or g6237(n2313 ,n1962 ,n1926);
    nand g6238(n9[34] ,n5136 ,n6154);
    or g6239(n4623 ,n3798 ,n4547);
    nor g6240(n5666 ,n4792 ,n5483);
    nand g6241(n7150 ,n6612 ,n6702);
    not g6242(n1960 ,n720);
    nand g6243(n906 ,n0[42] ,n724);
    nand g6244(n2029 ,n723 ,n1032);
    nor g6245(n2797 ,n1221 ,n2326);
    nand g6246(n4127 ,n2560 ,n3946);
    nand g6247(n4831 ,n1966 ,n4457);
    xnor g6248(n6509 ,n6385 ,n1556);
    nand g6249(n1906 ,n0[1] ,n972);
    nand g6250(n528 ,n0[96] ,n6953);
    nand g6251(n4405 ,n794 ,n4221);
    xnor g6252(n6885 ,n402 ,n433);
    xor g6253(n7116 ,n0[56] ,n0[24]);
    nand g6254(n6822 ,n6581 ,n7092);
    nor g6255(n4246 ,n1959 ,n3827);
    not g6256(n4878 ,n4877);
    nor g6257(n1775 ,n0[88] ,n1008);
    nand g6258(n6768 ,n0[40] ,n6737);
    xnor g6259(n6906 ,n255 ,n291);
    nor g6260(n1014 ,n0[89] ,n0[88]);
    nand g6261(n4651 ,n4008 ,n4529);
    xnor g6262(n1250 ,n6885 ,n6884);
    not g6263(n1962 ,n720);
    nand g6264(n4493 ,n792 ,n4359);
    xnor g6265(n4435 ,n2827 ,n3955);
    nand g6266(n260 ,n184 ,n259);
    xnor g6267(n1372 ,n6854 ,n6852);
    nor g6268(n5869 ,n713 ,n5730);
    nor g6269(n6018 ,n3441 ,n5893);
    xnor g6270(n2962 ,n1709 ,n1626);
    or g6271(n3026 ,n2290 ,n2289);
    nand g6272(n6743 ,n0[44] ,n6737);
    nand g6273(n4717 ,n3514 ,n4552);
    nor g6274(n6353 ,n5982 ,n6282);
    nor g6275(n4284 ,n762 ,n3884);
    nor g6276(n5259 ,n4304 ,n5025);
    nand g6277(n9[26] ,n6052 ,n6458);
    xnor g6278(n1602 ,n0[37] ,n0[21]);
    nand g6279(n2515 ,n1891 ,n1848);
    xor g6280(n693 ,n4213 ,n5158);
    nand g6281(n5530 ,n5326 ,n5252);
    xnor g6282(n241 ,n1[37] ,n0[37]);
    nand g6283(n509 ,n0[111] ,n6968);
    xnor g6284(n2829 ,n0[112] ,n1316);
    nand g6285(n6148 ,n3285 ,n6050);
    nand g6286(n4512 ,n3993 ,n4171);
    nor g6287(n4660 ,n2234 ,n4469);
    xnor g6288(n1521 ,n0[19] ,n1[19]);
    nor g6289(n4101 ,n2721 ,n3660);
    xnor g6290(n1919 ,n1[28] ,n2[28]);
    nor g6291(n4382 ,n3733 ,n4251);
    nand g6292(n571 ,n516 ,n570);
    xnor g6293(n2840 ,n1253 ,n1680);
    nand g6294(n1805 ,n794 ,n935);
    xor g6295(n7106 ,n0[46] ,n0[14]);
    or g6296(n4174 ,n2178 ,n3887);
    nand g6297(n1157 ,n6835 ,n795);
    nand g6298(n677 ,n1[17] ,n621);
    nand g6299(n4356 ,n7151 ,n3904);
    xnor g6300(n1943 ,n1[82] ,n2[18]);
    nand g6301(n3083 ,n1220 ,n2365);
    nand g6302(n2967 ,n1220 ,n2380);
    nand g6303(n6401 ,n3358 ,n6328);
    xnor g6304(n2798 ,n1384 ,n1362);
    nand g6305(n602 ,n482 ,n601);
    xnor g6306(n5751 ,n4666 ,n5464);
    nand g6307(n6685 ,n0[125] ,n0[93]);
    xnor g6308(n1358 ,n0[73] ,n4[1]);
    xnor g6309(n1523 ,n0[10] ,n1[10]);
    xnor g6310(n4893 ,n2840 ,n4449);
    nor g6311(n5440 ,n2325 ,n5275);
    nor g6312(n2264 ,n1958 ,n1615);
    xnor g6313(n1300 ,n0[100] ,n7096);
    nor g6314(n6397 ,n5549 ,n6317);
    nand g6315(n4354 ,n3666 ,n4029);
    xnor g6316(n1648 ,n0[38] ,n1[54]);
    nand g6317(n9[114] ,n4505 ,n6184);
    nand g6318(n3384 ,n2200 ,n2779);
    nor g6319(n6388 ,n712 ,n6314);
    or g6320(n4601 ,n711 ,n4582);
    nand g6321(n3743 ,n7158 ,n3165);
    xnor g6322(n5589 ,n5198 ,n1248);
    nor g6323(n4941 ,n4207 ,n4745);
    xnor g6324(n5199 ,n1715 ,n4879);
    nor g6325(n3465 ,n1954 ,n2939);
    xnor g6326(n1937 ,n1[11] ,n2[11]);
    nand g6327(n7019 ,n6698 ,n7154);
    not g6328(n6201 ,n6200);
    nand g6329(n112 ,n27 ,n111);
    xnor g6330(n1315 ,n6878 ,n6876);
    nand g6331(n59 ,n7074 ,n0[18]);
    nand g6332(n657 ,n1[26] ,n621);
    nor g6333(n3575 ,n2013 ,n3115);
    xnor g6334(n6113 ,n5846 ,n5945);
    xnor g6335(n5734 ,n5454 ,n2680);
    nor g6336(n2333 ,n0[61] ,n1958);
    xnor g6337(n2703 ,n1702 ,n1549);
    or g6338(n2152 ,n1962 ,n1438);
    nand g6339(n934 ,n0[58] ,n724);
    nand g6340(n3452 ,n1952 ,n2936);
    nand g6341(n3254 ,n906 ,n2199);
    nand g6342(n5763 ,n1953 ,n5708);
    nand g6343(n5403 ,n692 ,n5225);
    or g6344(n4147 ,n3769 ,n4054);
    xnor g6345(n1600 ,n0[108] ,n1[108]);
    nor g6346(n1964 ,n7090 ,n1232);
    nand g6347(n158 ,n18 ,n157);
    nor g6348(n2633 ,n0[11] ,n1963);
    not g6349(n2944 ,n2943);
    nand g6350(n206 ,n0[56] ,n1[56]);
    xnor g6351(n2662 ,n1[107] ,n1576);
    nor g6352(n1800 ,n731 ,n1220);
    nand g6353(n5911 ,n5526 ,n5759);
    nor g6354(n3052 ,n1798 ,n2185);
    nor g6355(n860 ,n1[64] ,n2[0]);
    nand g6356(n3875 ,n3245 ,n3585);
    xor g6357(n4898 ,n4212 ,n4586);
    nand g6358(n1061 ,n0[93] ,n710);
    nand g6359(n3621 ,n1[44] ,n2795);
    nand g6360(n6998 ,n6666 ,n6810);
    nor g6361(n4652 ,n6 ,n4453);
    nand g6362(n2597 ,n0[0] ,n707);
    xnor g6363(n5571 ,n1559 ,n5277);
    nand g6364(n5805 ,n4314 ,n5622);
    nand g6365(n6957 ,n6759 ,n6792);
    or g6366(n37 ,n7073 ,n0[17]);
    nor g6367(n3370 ,n1954 ,n2863);
    nor g6368(n5157 ,n2284 ,n4884);
    nand g6369(n1152 ,n6865 ,n795);
    nor g6370(n2249 ,n1963 ,n1509);
    nor g6371(n6246 ,n5670 ,n6144);
    nand g6372(n7046 ,n6683 ,n7127);
    nor g6373(n2476 ,n1000 ,n1768);
    nand g6374(n5325 ,n788 ,n5074);
    nand g6375(n5555 ,n4820 ,n5233);
    nor g6376(n1792 ,n0[17] ,n869);
    nor g6377(n4469 ,n793 ,n4211);
    xnor g6378(n1645 ,n0[97] ,n4[9]);
    nor g6379(n6555 ,n711 ,n6511);
    nor g6380(n6031 ,n3605 ,n5867);
    nand g6381(n3997 ,n3663 ,n3731);
    xnor g6382(n1542 ,n0[12] ,n1[12]);
    xnor g6383(n5726 ,n4805 ,n5455);
    nand g6384(n1196 ,n6940 ,n796);
    nand g6385(n6160 ,n3339 ,n6040);
    nand g6386(n5971 ,n4149 ,n5888);
    nand g6387(n5470 ,n4702 ,n5330);
    xnor g6388(n91 ,n0[7] ,n7063);
    nand g6389(n117 ,n61 ,n116);
    not g6390(n731 ,n0[106]);
    nand g6391(n594 ,n471 ,n593);
    nand g6392(n7080 ,n671 ,n641);
    nand g6393(n9[45] ,n5451 ,n6063);
    or g6394(n700 ,n6002 ,n5782);
    nor g6395(n5450 ,n2325 ,n5376);
    nor g6396(n4447 ,n4254 ,n4204);
    nand g6397(n5251 ,n4967 ,n5069);
    nand g6398(n2555 ,n1230 ,n1909);
    nor g6399(n899 ,n1[5] ,n2[5]);
    nor g6400(n6350 ,n706 ,n6311);
    xnor g6401(n84 ,n7087 ,n0[31]);
    nand g6402(n109 ,n69 ,n108);
    not g6403(n5936 ,n5935);
    nand g6404(n5744 ,n1953 ,n5581);
    nor g6405(n5046 ,n3449 ,n4891);
    nand g6406(n1129 ,n6908 ,n796);
    not g6407(n3809 ,n3790);
    xnor g6408(n546 ,n6959 ,n0[102]);
    nor g6409(n1871 ,n0[17] ,n976);
    nand g6410(n993 ,n0[27] ,n723);
    nor g6411(n5082 ,n2745 ,n4962);
    or g6412(n3297 ,n2407 ,n3253);
    nand g6413(n5685 ,n3464 ,n5397);
    nand g6414(n5699 ,n4861 ,n5469);
    nor g6415(n2916 ,n1865 ,n2609);
    xor g6416(n691 ,n2656 ,n5061);
    or g6417(n344 ,n7024 ,n6992);
    nand g6418(n4799 ,n4500 ,n4492);
    nand g6419(n6532 ,n5538 ,n6491);
    nand g6420(n5006 ,n4802 ,n4752);
    xnor g6421(n5208 ,n4840 ,n1578);
    nand g6422(n7060 ,n659 ,n650);
    or g6423(n3389 ,n1954 ,n2919);
    nor g6424(n4962 ,n988 ,n4781);
    nor g6425(n5367 ,n3798 ,n5149);
    nor g6426(n6439 ,n6379 ,n6145);
    xnor g6427(n3837 ,n1[79] ,n2672);
    or g6428(n470 ,n0[100] ,n6957);
    nor g6429(n2236 ,n719 ,n1611);
    nor g6430(n5964 ,n1954 ,n5851);
    nand g6431(n3142 ,n2580 ,n2419);
    xnor g6432(n1583 ,n0[123] ,n1[123]);
    nand g6433(n3134 ,n1[62] ,n2385);
    nor g6434(n2590 ,n0[48] ,n1788);
    nand g6435(n4569 ,n2527 ,n4216);
    xnor g6436(n2957 ,n1330 ,n1595);
    nand g6437(n6138 ,n6075 ,n6065);
    nor g6438(n4632 ,n3529 ,n4545);
    not g6439(n727 ,n6827);
    nand g6440(n6008 ,n5598 ,n5928);
    or g6441(n323 ,n7042 ,n7010);
    xnor g6442(n1433 ,n1[1] ,n2[1]);
    nor g6443(n3537 ,n6825 ,n2853);
    nand g6444(n3399 ,n1953 ,n2921);
    or g6445(n5846 ,n3442 ,n5718);
    nand g6446(n6794 ,n1[101] ,n7088);
    xnor g6447(n2857 ,n1336 ,n1629);
    xnor g6448(n1704 ,n0[75] ,n4[3]);
    nand g6449(n5693 ,n4618 ,n5396);
    nand g6450(n5353 ,n4331 ,n5172);
    xnor g6451(n4908 ,n2835 ,n4433);
    nand g6452(n2795 ,n788 ,n2326);
    nor g6453(n6143 ,n4854 ,n6069);
    nand g6454(n4588 ,n3198 ,n4347);
    nor g6455(n2054 ,n1958 ,n1509);
    nand g6456(n1980 ,n1092 ,n950);
    not g6457(n4576 ,n4577);
    nor g6458(n5841 ,n4412 ,n5718);
    or g6459(n165 ,n0[51] ,n1[51]);
    nand g6460(n1193 ,n6872 ,n795);
    or g6461(n4060 ,n3657 ,n3510);
    nand g6462(n5537 ,n4830 ,n5359);
    nand g6463(n136 ,n37 ,n135);
    nor g6464(n3922 ,n2437 ,n3766);
    nor g6465(n6016 ,n3405 ,n5878);
    nand g6466(n3131 ,n2427 ,n2474);
    nor g6467(n987 ,n738 ,n0[114]);
    nand g6468(n3540 ,n6 ,n2720);
    nand g6469(n4104 ,n3557 ,n3459);
    nor g6470(n5085 ,n6824 ,n4896);
    not g6471(n4362 ,n4361);
    nand g6472(n3843 ,n1965 ,n3461);
    nand g6473(n4788 ,n3034 ,n4516);
    nor g6474(n3295 ,n1954 ,n2867);
    xnor g6475(n1472 ,n1[125] ,n2[61]);
    nor g6476(n3615 ,n770 ,n2974);
    xor g6477(n689 ,n3948 ,n2799);
    nand g6478(n201 ,n0[59] ,n1[59]);
    nand g6479(n1898 ,n0[59] ,n1221);
    xnor g6480(n1414 ,n1[78] ,n2[14]);
    nor g6481(n6229 ,n3782 ,n6125);
    nand g6482(n4355 ,n2156 ,n4084);
    xnor g6483(n1938 ,n1[87] ,n2[23]);
    or g6484(n6823 ,n3[1] ,n6735);
    nand g6485(n5712 ,n5169 ,n5437);
    not g6486(n1234 ,n1233);
    not g6487(n1952 ,n1954);
    nor g6488(n4614 ,n727 ,n4476);
    nand g6489(n6615 ,n0[68] ,n6579);
    not g6490(n5997 ,n5996);
    nand g6491(n965 ,n794 ,n708);
    xnor g6492(n1427 ,n1[109] ,n2[45]);
    nor g6493(n6372 ,n3341 ,n6251);
    nand g6494(n4098 ,n2417 ,n3570);
    or g6495(n4186 ,n1960 ,n3832);
    xnor g6496(n100 ,n0[16] ,n7072);
    nand g6497(n6292 ,n3555 ,n6180);
    nand g6498(n194 ,n0[53] ,n1[53]);
    nand g6499(n3434 ,n709 ,n2916);
    nand g6500(n5381 ,n4829 ,n5119);
    nor g6501(n4932 ,n4357 ,n4742);
    or g6502(n4692 ,n1965 ,n4455);
    nand g6503(n5502 ,n4686 ,n5313);
    nand g6504(n4570 ,n1085 ,n4215);
    nor g6505(n2061 ,n1957 ,n1492);
    xnor g6506(n1279 ,n0[127] ,n7123);
    or g6507(n4657 ,n3513 ,n4541);
    xnor g6508(n1492 ,n0[0] ,n1[0]);
    not g6509(n4806 ,n4807);
    nand g6510(n3718 ,n2184 ,n3199);
    nor g6511(n5348 ,n4717 ,n5189);
    xnor g6512(n1273 ,n1[68] ,n4[12]);
    nand g6513(n5643 ,n6 ,n5445);
    nand g6514(n5091 ,n4237 ,n4960);
    not g6515(n2575 ,n2574);
    xnor g6516(n1641 ,n0[23] ,n1[23]);
    not g6517(n5079 ,n5078);
    xnor g6518(n6919 ,n75 ,n145);
    nor g6519(n5915 ,n5801 ,n5388);
    nand g6520(n6272 ,n6221 ,n6222);
    nor g6521(n5815 ,n4399 ,n5711);
    xor g6522(n3831 ,n2666 ,n1[68]);
    nand g6523(n6295 ,n6152 ,n6206);
    xnor g6524(n1519 ,n0[2] ,n1[2]);
    xor g6525(n7098 ,n0[38] ,n0[6]);
    or g6526(n4230 ,n792 ,n3839);
    nand g6527(n4239 ,n1966 ,n3938);
    or g6528(n4619 ,n2561 ,n4449);
    not g6529(n4875 ,n4876);
    nor g6530(n6559 ,n5168 ,n6517);
    xnor g6531(n1319 ,n6949 ,n6948);
    nor g6532(n2052 ,n1962 ,n1455);
    nand g6533(n3639 ,n1[55] ,n2988);
    nor g6534(n6529 ,n6384 ,n6505);
    nand g6535(n3248 ,n917 ,n2050);
    or g6536(n9[101] ,n5665 ,n6156);
    nor g6537(n2037 ,n1963 ,n1482);
    nand g6538(n1863 ,n0[49] ,n1221);
    nor g6539(n2196 ,n1956 ,n1613);
    nand g6540(n9[22] ,n5740 ,n5804);
    xnor g6541(n3956 ,n2823 ,n2805);
    not g6542(n5081 ,n5080);
    not g6543(n5645 ,n5637);
    nor g6544(n4358 ,n4015 ,n3892);
    nand g6545(n6535 ,n6484 ,n6502);
    xor g6546(n5287 ,n4211 ,n5002);
    nand g6547(n6764 ,n0[49] ,n6737);
    xnor g6548(n5956 ,n5206 ,n5724);
    xnor g6549(n1559 ,n0[61] ,n4[21]);
    nor g6550(n3353 ,n1[49] ,n3144);
    nor g6551(n6702 ,n6826 ,n6605);
    nor g6552(n4492 ,n2543 ,n4172);
    nor g6553(n5186 ,n6824 ,n4911);
    nor g6554(n5603 ,n706 ,n5422);
    xnor g6555(n6175 ,n5934 ,n6034);
    xnor g6556(n1409 ,n1[58] ,n2[58]);
    nand g6557(n1207 ,n1[5] ,n2[5]);
    nand g6558(n6496 ,n6452 ,n6346);
    xnor g6559(n2862 ,n1633 ,n1575);
    xnor g6560(n6837 ,n390 ,n409);
    nor g6561(n6728 ,n6826 ,n6604);
    nand g6562(n4378 ,n791 ,n4235);
    nor g6563(n3512 ,n6825 ,n2825);
    nand g6564(n3628 ,n2443 ,n2786);
    nor g6565(n2004 ,n867 ,n923);
    nor g6566(n4375 ,n722 ,n4368);
    xnor g6567(n6343 ,n6244 ,n6173);
    xnor g6568(n1608 ,n0[126] ,n0[110]);
    xnor g6569(n1636 ,n0[122] ,n1[122]);
    nand g6570(n2503 ,n1235 ,n1998);
    nor g6571(n4180 ,n3225 ,n3929);
    nand g6572(n4364 ,n2016 ,n3845);
    xnor g6573(n2851 ,n1370 ,n1341);
    nand g6574(n4496 ,n3016 ,n4339);
    nor g6575(n1874 ,n760 ,n11);
    or g6576(n2184 ,n719 ,n1632);
    xnor g6577(n1656 ,n0[40] ,n0[24]);
    nand g6578(n5617 ,n4940 ,n5472);
    nand g6579(n5610 ,n4197 ,n5544);
    nand g6580(n3601 ,n0[103] ,n2794);
    nor g6581(n6710 ,n6826 ,n6586);
    nor g6582(n6398 ,n712 ,n701);
    not g6583(n824 ,n0[12]);
    nor g6584(n1086 ,n840 ,n790);
    nor g6585(n3984 ,n708 ,n3794);
    xnor g6586(n4902 ,n2837 ,n4466);
    nand g6587(n2540 ,n1157 ,n1853);
    nor g6588(n2790 ,n2328 ,n2608);
    nor g6589(n4085 ,n6802 ,n3726);
    nor g6590(n2759 ,n1515 ,n2630);
    not g6591(n776 ,n1[55]);
    nand g6592(n3768 ,n7130 ,n3059);
    xnor g6593(n2861 ,n1349 ,n1491);
    nand g6594(n6964 ,n6741 ,n6772);
    xnor g6595(n5265 ,n4876 ,n5002);
    nand g6596(n5793 ,n5534 ,n5629);
    nand g6597(n4543 ,n1118 ,n4139);
    nand g6598(n6235 ,n3397 ,n6123);
    nand g6599(n1211 ,n7089 ,n7091);
    nand g6600(n7089 ,n3[0] ,n6730);
    nor g6601(n2808 ,n1864 ,n2585);
    nand g6602(n5676 ,n4191 ,n5536);
    nand g6603(n3614 ,n1[46] ,n2973);
    nand g6604(n6224 ,n3414 ,n6139);
    nand g6605(n1244 ,n0[67] ,n723);
    nand g6606(n510 ,n0[120] ,n6977);
    nor g6607(n1740 ,n0[58] ,n996);
    nor g6608(n4003 ,n836 ,n3272);
    xnor g6609(n2954 ,n1704 ,n1591);
    nand g6610(n6752 ,n0[62] ,n6737);
    nor g6611(n6378 ,n5385 ,n6263);
    xnor g6612(n95 ,n0[11] ,n7067);
    nor g6613(n1643 ,n1049 ,n1051);
    or g6614(n2421 ,n1960 ,n1424);
    not g6615(n2637 ,n2636);
    or g6616(n339 ,n7025 ,n6993);
    nand g6617(n4235 ,n3280 ,n3857);
    xnor g6618(n1321 ,n0[123] ,n7119);
    nor g6619(n6362 ,n6252 ,n6281);
    nand g6620(n6757 ,n0[63] ,n6737);
    nor g6621(n3508 ,n6825 ,n2817);
    not g6622(n2600 ,n2599);
    nand g6623(n46 ,n7078 ,n0[22]);
    or g6624(n4121 ,n2561 ,n3943);
    not g6625(n728 ,n0[81]);
    nor g6626(n3471 ,n1954 ,n2944);
    nand g6627(n6755 ,n0[50] ,n6737);
    nand g6628(n6271 ,n6140 ,n6220);
    nor g6629(n4254 ,n708 ,n4111);
    nand g6630(n6635 ,n0[109] ,n0[77]);
    not g6631(n784 ,n6909);
    xnor g6632(n2720 ,n1723 ,n1502);
    nor g6633(n3494 ,n2327 ,n3131);
    nor g6634(n2209 ,n1961 ,n1934);
    nor g6635(n6042 ,n711 ,n5969);
    or g6636(n5797 ,n4342 ,n5679);
    or g6637(n2087 ,n1961 ,n1447);
    not g6638(n2325 ,n2326);
    xnor g6639(n1569 ,n839 ,n1[0]);
    nor g6640(n4631 ,n3505 ,n4544);
    nand g6641(n1233 ,n0[32] ,n714);
    nand g6642(n943 ,n0[23] ,n708);
    nand g6643(n4544 ,n1139 ,n4129);
    nand g6644(n210 ,n0[36] ,n1[36]);
    nand g6645(n129 ,n47 ,n128);
    not g6646(n981 ,n980);
    xnor g6647(n2874 ,n1353 ,n1596);
    nand g6648(n2767 ,n1504 ,n2628);
    or g6649(n9[42] ,n4790 ,n6182);
    not g6650(n1041 ,n1040);
    nand g6651(n933 ,n0[10] ,n724);
    nand g6652(n2512 ,n793 ,n1974);
    xnor g6653(n6512 ,n6305 ,n6415);
    nor g6654(n5616 ,n5414 ,n5409);
    nor g6655(n6431 ,n3398 ,n702);
    xnor g6656(n1669 ,n0[47] ,n1[63]);
    nor g6657(n2318 ,n721 ,n1491);
    nand g6658(n5222 ,n4889 ,n5032);
    not g6659(n5076 ,n5075);
    xnor g6660(n2863 ,n1598 ,n1517);
    nor g6661(n6538 ,n5474 ,n6507);
    xnor g6662(n5854 ,n694 ,n1585);
    nand g6663(n5167 ,n4243 ,n4984);
    nand g6664(n2308 ,n792 ,n1991);
    not g6665(n2605 ,n2604);
    nor g6666(n3405 ,n1954 ,n2940);
    nand g6667(n4272 ,n2068 ,n3972);
    nand g6668(n430 ,n340 ,n429);
    nand g6669(n6105 ,n4493 ,n5978);
    xnor g6670(n6886 ,n250 ,n281);
    or g6671(n2791 ,n1514 ,n2642);
    nor g6672(n2986 ,n2590 ,n2585);
    nand g6673(n4238 ,n1966 ,n3945);
    nand g6674(n5050 ,n3269 ,n4898);
    nor g6675(n3481 ,n1954 ,n2948);
    nor g6676(n1023 ,n741 ,n0[81]);
    nand g6677(n1890 ,n0[124] ,n1221);
    nand g6678(n6136 ,n6062 ,n6064);
    xnor g6679(n6903 ,n102 ,n137);
    nor g6680(n4634 ,n3499 ,n4546);
    nor g6681(n3028 ,n0[96] ,n2323);
    or g6682(n9[94] ,n5256 ,n5716);
    xnor g6683(n1281 ,n0[117] ,n4[5]);
    or g6684(n3565 ,n1954 ,n2958);
    xnor g6685(n3817 ,n1[85] ,n2685);
    xnor g6686(n2902 ,n1686 ,n1630);
    nor g6687(n957 ,n0[114] ,n0[112]);
    nand g6688(n1902 ,n0[90] ,n1018);
    xnor g6689(n2674 ,n0[126] ,n1249);
    nor g6690(n4612 ,n727 ,n4477);
    nor g6691(n1176 ,n784 ,n716);
    nand g6692(n7057 ,n674 ,n648);
    nor g6693(n4163 ,n722 ,n3954);
    nand g6694(n4813 ,n1966 ,n4435);
    xnor g6695(n2879 ,n1303 ,n1649);
    nand g6696(n4508 ,n3702 ,n4176);
    or g6697(n5126 ,n2325 ,n5007);
    nor g6698(n4851 ,n722 ,n4682);
    xnor g6699(n2854 ,n1306 ,n1692);
    nand g6700(n5973 ,n4643 ,n5888);
    xnor g6701(n1630 ,n0[105] ,n1[105]);
    nor g6702(n2373 ,n1[44] ,n719);
    or g6703(n3913 ,n2766 ,n3774);
    nand g6704(n6999 ,n6672 ,n6809);
    nand g6705(n642 ,n0[64] ,n622);
    nand g6706(n9[107] ,n6543 ,n6576);
    nand g6707(n5036 ,n4860 ,n4888);
    nor g6708(n5908 ,n4354 ,n5819);
    nor g6709(n3547 ,n1954 ,n2962);
    xnor g6710(n2890 ,n1301 ,n1653);
    xnor g6711(n6945 ,n386 ,n463);
    nor g6712(n980 ,n725 ,n0[59]);
    xnor g6713(n1457 ,n0[126] ,n1[126]);
    or g6714(n5217 ,n4062 ,n5130);
    nand g6715(n105 ,n51 ,n104);
    xnor g6716(n1473 ,n1[3] ,n2[3]);
    xnor g6717(n1603 ,n0[104] ,n1[104]);
    or g6718(n345 ,n7044 ,n7012);
    nor g6719(n2727 ,n1030 ,n2609);
    nand g6720(n1095 ,n0[81] ,n0[80]);
    nor g6721(n874 ,n725 ,n0[8]);
    nand g6722(n5214 ,n4938 ,n5081);
    nand g6723(n2553 ,n1133 ,n1897);
    or g6724(n2973 ,n2629 ,n2348);
    nor g6725(n3284 ,n1222 ,n2809);
    nand g6726(n504 ,n0[113] ,n6970);
    xnor g6727(n2681 ,n1[101] ,n1544);
    nand g6728(n922 ,n0[66] ,n724);
    nor g6729(n4459 ,n4262 ,n4120);
    nor g6730(n1738 ,n1052 ,n942);
    nor g6731(n2128 ,n905 ,n1962);
    nor g6732(n2268 ,n1961 ,n1410);
    nand g6733(n5508 ,n3347 ,n5224);
    nand g6734(n5545 ,n4813 ,n5362);
    nor g6735(n857 ,n791 ,n0[101]);
    nor g6736(n1875 ,n769 ,n11);
    not g6737(n1504 ,n1503);
    xnor g6738(n389 ,n6987 ,n7019);
    nand g6739(n9[54] ,n5034 ,n5627);
    nor g6740(n6360 ,n5776 ,n6283);
    not g6741(n6212 ,n6211);
    xnor g6742(n1934 ,n1[91] ,n2[27]);
    nand g6743(n2009 ,n0[88] ,n1008);
    or g6744(n3387 ,n3002 ,n2268);
    xnor g6745(n4478 ,n3943 ,n2810);
    nand g6746(n3666 ,n0[13] ,n3094);
    xnor g6747(n6417 ,n6280 ,n6309);
    xnor g6748(n1700 ,n0[98] ,n4[10]);
    xnor g6749(n1507 ,n0[24] ,n1[24]);
    or g6750(n2776 ,n1579 ,n2635);
    nand g6751(n7076 ,n672 ,n625);
    nand g6752(n5517 ,n5250 ,n5281);
    nor g6753(n6055 ,n5896 ,n5977);
    nor g6754(n4412 ,n6 ,n4219);
    nand g6755(n347 ,n7047 ,n7015);
    or g6756(n9[41] ,n4799 ,n6412);
    nand g6757(n1057 ,n0[125] ,n789);
    nand g6758(n4553 ,n1160 ,n4128);
    nand g6759(n2458 ,n0[83] ,n2015);
    xnor g6760(n6924 ,n533 ,n605);
    xnor g6761(n6196 ,n6108 ,n5833);
    nand g6762(n5008 ,n2507 ,n4674);
    nor g6763(n6300 ,n6229 ,n6203);
    or g6764(n6137 ,n711 ,n6105);
    not g6765(n732 ,n0[15]);
    nor g6766(n3107 ,n1874 ,n2034);
    not g6767(n714 ,n724);
    nand g6768(n2447 ,n0[58] ,n718);
    xnor g6769(n5445 ,n4593 ,n5017);
    nor g6770(n2561 ,n845 ,n1966);
    nand g6771(n4106 ,n1904 ,n3549);
    nand g6772(n928 ,n0[13] ,n709);
    nand g6773(n3385 ,n2465 ,n2778);
    nand g6774(n6960 ,n6765 ,n6798);
    nor g6775(n2399 ,n0[117] ,n1958);
    xnor g6776(n1661 ,n6910 ,n6911);
    nand g6777(n6560 ,n4730 ,n6520);
    not g6778(n2935 ,n2934);
    not g6779(n5840 ,n5841);
    nand g6780(n10[0] ,n4941 ,n4708);
    nand g6781(n9[98] ,n5112 ,n6135);
    nand g6782(n3644 ,n0[54] ,n2796);
    nand g6783(n6164 ,n5889 ,n6074);
    nand g6784(n6647 ,n0[73] ,n6580);
    nand g6785(n5111 ,n710 ,n5011);
    nand g6786(n5950 ,n1953 ,n5855);
    nor g6787(n2134 ,n6 ,n1756);
    nor g6788(n5272 ,n794 ,n5055);
    nand g6789(n998 ,n0[65] ,n820);
    nand g6790(n6766 ,n0[53] ,n6737);
    nand g6791(n6681 ,n0[124] ,n0[92]);
    xnor g6792(n2692 ,n1[115] ,n1496);
    nor g6793(n1768 ,n0[32] ,n1047);
    nor g6794(n6571 ,n5673 ,n6557);
    nor g6795(n1824 ,n739 ,n11);
    nand g6796(n6807 ,n6581 ,n7107);
    nand g6797(n5880 ,n5762 ,n5755);
    nand g6798(n2570 ,n0[31] ,n707);
    xnor g6799(n2702 ,n0[120] ,n1490);
    nand g6800(n2508 ,n0[59] ,n2017);
    nand g6801(n212 ,n0[38] ,n1[38]);
    nand g6802(n2752 ,n1513 ,n2618);
    nand g6803(n4510 ,n3703 ,n4175);
    nor g6804(n4529 ,n4292 ,n4316);
    or g6805(n472 ,n0[116] ,n6973);
    nand g6806(n6989 ,n6697 ,n6819);
    nor g6807(n6430 ,n3381 ,n6323);
    not g6808(n738 ,n0[112]);
    nand g6809(n5879 ,n5566 ,n5757);
    xnor g6810(n1673 ,n0[34] ,n1[50]);
    or g6811(n181 ,n0[61] ,n1[61]);
    nand g6812(n6979 ,n6769 ,n6782);
    not g6813(n848 ,n6877);
    or g6814(n33 ,n7064 ,n0[8]);
    nor g6815(n4470 ,n793 ,n4213);
    xnor g6816(n1420 ,n1[17] ,n2[17]);
    nor g6817(n5038 ,n712 ,n4999);
    nor g6818(n5608 ,n5097 ,n5466);
    nor g6819(n5090 ,n6824 ,n4897);
    xnor g6820(n4463 ,n3946 ,n2826);
    nand g6821(n1209 ,n1[117] ,n2[53]);
    nand g6822(n588 ,n478 ,n587);
    xnor g6823(n6892 ,n556 ,n589);
    nand g6824(n988 ,n723 ,n760);
    not g6825(n801 ,n0[18]);
    xnor g6826(n86 ,n0[2] ,n7058);
    or g6827(n5153 ,n4060 ,n4979);
    nand g6828(n276 ,n164 ,n275);
    nor g6829(n2441 ,n0[5] ,n1545);
    or g6830(n14 ,n7060 ,n0[4]);
    xnor g6831(n5593 ,n5266 ,n2653);
    nand g6832(n3178 ,n1988 ,n2326);
    nand g6833(n6672 ,n0[77] ,n6580);
    nand g6834(n2478 ,n0[12] ,n1964);
    nor g6835(n2777 ,n2054 ,n2105);
    nand g6836(n681 ,n1[25] ,n621);
    nand g6837(n1150 ,n6883 ,n796);
    xnor g6838(n2838 ,n0[116] ,n1342);
    or g6839(n2307 ,n715 ,n1429);
    xnor g6840(n1644 ,n1[23] ,n4[23]);
    nor g6841(n6254 ,n6006 ,n6214);
    nand g6842(n6965 ,n6743 ,n6774);
    nand g6843(n6285 ,n6226 ,n6211);
    nand g6844(n66 ,n7065 ,n0[9]);
    nand g6845(n353 ,n7045 ,n7013);
    nand g6846(n1030 ,n0[90] ,n809);
    nor g6847(n1802 ,n800 ,n1220);
    nand g6848(n6325 ,n717 ,n6309);
    nand g6849(n307 ,n220 ,n306);
    nor g6850(n5120 ,n3267 ,n4898);
    xnor g6851(n1330 ,n0[99] ,n4[11]);
    nor g6852(n4958 ,n3530 ,n4774);
    xnor g6853(n1271 ,n6865 ,n6864);
    nand g6854(n1081 ,n0[28] ,n787);
    nor g6855(n3487 ,n6 ,n2808);
    nor g6856(n5627 ,n5520 ,n5532);
    nor g6857(n5803 ,n1954 ,n5591);
    nand g6858(n6610 ,n0[100] ,n0[68]);
    nand g6859(n1243 ,n0[50] ,n723);
    nand g6860(n5761 ,n1953 ,n5586);
    nor g6861(n4945 ,n2325 ,n4808);
    xnor g6862(n2923 ,n1340 ,n1631);
    or g6863(n2085 ,n1034 ,n1729);
    nor g6864(n4249 ,n1960 ,n3837);
    xnor g6865(n1698 ,n0[66] ,n1[82]);
    or g6866(n2992 ,n2623 ,n2402);
    or g6867(n3564 ,n791 ,n3260);
    nand g6868(n1840 ,n0[5] ,n1221);
    xnor g6869(n78 ,n0[25] ,n7081);
    nor g6870(n6393 ,n3336 ,n6322);
    or g6871(n2056 ,n1961 ,n1454);
    xnor g6872(n6121 ,n5391 ,n5941);
    nand g6873(n4564 ,n1170 ,n4125);
    nor g6874(n873 ,n0[67] ,n0[66]);
    not g6875(n789 ,n791);
    nor g6876(n5345 ,n4737 ,n5184);
    nor g6877(n5827 ,n4330 ,n5684);
    xnor g6878(n255 ,n1[51] ,n0[51]);
    or g6879(n5344 ,n5117 ,n5160);
    nor g6880(n5319 ,n4738 ,n5181);
    xnor g6881(n1604 ,n0[97] ,n1[97]);
    not g6882(n791 ,n8);
    nand g6883(n5363 ,n3514 ,n5144);
    xnor g6884(n1544 ,n1[37] ,n1[5]);
    nor g6885(n2304 ,n1956 ,n1916);
    nor g6886(n2381 ,n0[36] ,n1958);
    nand g6887(n429 ,n375 ,n428);
    nor g6888(n3458 ,n2291 ,n3026);
    nand g6889(n1098 ,n0[79] ,n792);
    nand g6890(n6469 ,n6292 ,n6418);
    nand g6891(n7158 ,n6581 ,n7121);
    nand g6892(n1812 ,n0[42] ,n1221);
    nor g6893(n3065 ,n1826 ,n2310);
    not g6894(n837 ,n1[86]);
    nor g6895(n3038 ,n1221 ,n2345);
    xnor g6896(n1493 ,n1[47] ,n1[15]);
    or g6897(n4187 ,n1961 ,n3829);
    nand g6898(n4318 ,n792 ,n4102);
    nand g6899(n1154 ,n6852 ,n796);
    nor g6900(n4294 ,n732 ,n4018);
    or g6901(n3019 ,n2270 ,n2269);
    nor g6902(n872 ,n725 ,n0[18]);
    nand g6903(n5146 ,n6827 ,n4916);
    xnor g6904(n1448 ,n1[111] ,n2[47]);
    xor g6905(n3830 ,n2665 ,n1[71]);
    or g6906(n4143 ,n3361 ,n4081);
    nand g6907(n1989 ,n1057 ,n1060);
    nand g6908(n6614 ,n0[92] ,n6579);
    nor g6909(n5026 ,n4684 ,n4878);
    nor g6910(n2254 ,n1962 ,n1935);
    not g6911(n3247 ,n3246);
    or g6912(n3444 ,n789 ,n3258);
    nand g6913(n5978 ,n6 ,n5852);
    not g6914(n2583 ,n2582);
    nand g6915(n6808 ,n6581 ,n7106);
    not g6916(n2326 ,n722);
    nand g6917(n4286 ,n3999 ,n3853);
    nand g6918(n7009 ,n6682 ,n7164);
    xor g6919(n7113 ,n0[53] ,n0[21]);
    nand g6920(n4639 ,n2749 ,n4387);
    nor g6921(n3657 ,n742 ,n3085);
    nor g6922(n3480 ,n1954 ,n2889);
    nand g6923(n671 ,n1[24] ,n621);
    nor g6924(n4380 ,n722 ,n4363);
    xnor g6925(n5847 ,n5575 ,n3494);
    nor g6926(n2269 ,n1958 ,n1620);
    or g6927(n9[102] ,n5913 ,n5803);
    xnor g6928(n6875 ,n95 ,n123);
    nand g6929(n2574 ,n0[11] ,n1964);
    xnor g6930(n3939 ,n2674 ,n2833);
    not g6931(n3262 ,n3232);
    nand g6932(n1165 ,n6903 ,n795);
    nor g6933(n3531 ,n6825 ,n2841);
    nor g6934(n5298 ,n706 ,n5114);
    not g6935(n802 ,n0[80]);
    xnor g6936(n232 ,n1[59] ,n0[59]);
    nand g6937(n6824 ,n6732 ,n6733);
    nor g6938(n5242 ,n4852 ,n5124);
    nor g6939(n3045 ,n1793 ,n2314);
    nor g6940(n4711 ,n6824 ,n688);
    nand g6941(n3775 ,n7125 ,n2756);
    nor g6942(n870 ,n708 ,n0[15]);
    nand g6943(n6961 ,n6768 ,n6799);
    nor g6944(n4729 ,n2325 ,n4462);
    nor g6945(n6084 ,n6014 ,n5984);
    nand g6946(n2443 ,n1[62] ,n1483);
    nand g6947(n3292 ,n1952 ,n2918);
    xnor g6948(n3839 ,n2646 ,n2645);
    nor g6949(n3456 ,n1222 ,n2848);
    nand g6950(n2636 ,n817 ,n707);
    xnor g6951(n6845 ,n392 ,n413);
    nor g6952(n5504 ,n5246 ,n5294);
    or g6953(n2351 ,n721 ,n1569);
    nor g6954(n6322 ,n713 ,n6308);
    xnor g6955(n5724 ,n4456 ,n5531);
    xnor g6956(n5574 ,n5380 ,n5375);
    nand g6957(n3209 ,n1141 ,n2130);
    nand g6958(n3187 ,n2009 ,n2433);
    not g6959(n4925 ,n4924);
    xnor g6960(n235 ,n1[62] ,n0[62]);
    not g6961(n698 ,n699);
    nor g6962(n6332 ,n711 ,n6306);
    nor g6963(n5113 ,n4491 ,n4943);
    nand g6964(n1839 ,n0[34] ,n1221);
    xnor g6965(n2806 ,n0[118] ,n1267);
    nand g6966(n3586 ,n2456 ,n3105);
    xnor g6967(n230 ,n1[57] ,n0[57]);
    nor g6968(n6564 ,n5393 ,n6555);
    xnor g6969(n2669 ,n1985 ,n2001);
    xnor g6970(n6314 ,n6066 ,n6191);
    nor g6971(n5014 ,n2822 ,n4780);
    or g6972(n2077 ,n719 ,n1520);
    xnor g6973(n5390 ,n5016 ,n4459);
    xnor g6974(n5077 ,n4667 ,n4454);
    nor g6975(n4339 ,n2479 ,n4087);
    nand g6976(n1125 ,n6888 ,n796);
    nand g6977(n1140 ,n6831 ,n796);
    nand g6978(n5528 ,n5325 ,n5253);
    nand g6979(n3551 ,n1953 ,n2958);
    nor g6980(n6225 ,n1954 ,n6146);
    nand g6981(n610 ,n497 ,n609);
    nand g6982(n5562 ,n4692 ,n5229);
    nor g6983(n904 ,n0[98] ,n714);
    nor g6984(n2745 ,n1750 ,n2500);
    or g6985(n468 ,n0[107] ,n6964);
    nor g6986(n5766 ,n1954 ,n5592);
    nor g6987(n6019 ,n3484 ,n5897);
    nand g6988(n1120 ,n6927 ,n795);
    nand g6989(n1868 ,n0[30] ,n964);
    xnor g6990(n1581 ,n0[87] ,n4[31]);
    nand g6991(n3745 ,n7160 ,n3109);
    nand g6992(n54 ,n7080 ,n0[24]);
    nand g6993(n4265 ,n720 ,n3824);
    xnor g6994(n3958 ,n2820 ,n2803);
    nand g6995(n467 ,n366 ,n466);
    nand g6996(n591 ,n512 ,n590);
    nand g6997(n3750 ,n6809 ,n3114);
    nor g6998(n2188 ,n1956 ,n1591);
    or g6999(n2198 ,n1959 ,n1436);
    nand g7000(n9[68] ,n5794 ,n5899);
    nand g7001(n4773 ,n2560 ,n4442);
    nand g7002(n1160 ,n6949 ,n795);
    nand g7003(n2439 ,n0[43] ,n2019);
    nand g7004(n4201 ,n708 ,n3965);
    nor g7005(n5963 ,n1954 ,n5850);
    nor g7006(n999 ,n0[123] ,n0[120]);
    not g7007(n4712 ,n4711);
    nand g7008(n63 ,n7064 ,n0[8]);
    not g7009(n5897 ,n5896);
    nand g7010(n116 ,n35 ,n115);
    not g7011(n4475 ,n4474);
    nand g7012(n114 ,n40 ,n113);
    xnor g7013(n6909 ,n377 ,n445);
    nor g7014(n3582 ,n809 ,n2739);
    nand g7015(n3693 ,n2313 ,n3159);
    xnor g7016(n5061 ,n4805 ,n4429);
    nand g7017(n3120 ,n1[60] ,n2640);
    nand g7018(n1059 ,n0[47] ,n790);
    xnor g7019(n1393 ,n1[15] ,n2[15]);
    nor g7020(n2124 ,n980 ,n1752);
    nor g7021(n2073 ,n1958 ,n1523);
    nand g7022(n5903 ,n3298 ,n5748);
    xnor g7023(n5590 ,n5196 ,n5195);
    nor g7024(n4288 ,n4005 ,n3681);
    xnor g7025(n1284 ,n0[127] ,n0[15]);
    nand g7026(n6701 ,n1[89] ,n6580);
    not g7027(n4699 ,n4698);
    or g7028(n5696 ,n5382 ,n5408);
    nor g7029(n3560 ,n709 ,n3255);
    nand g7030(n511 ,n0[101] ,n6958);
    nor g7031(n1843 ,n746 ,n11);
    or g7032(n2316 ,n1959 ,n1449);
    nor g7033(n3850 ,n3592 ,n2724);
    nor g7034(n6458 ,n6241 ,n6361);
    xnor g7035(n4590 ,n4223 ,n4225);
    not g7036(n2567 ,n2566);
    nand g7037(n4736 ,n717 ,n4568);
    nor g7038(n6443 ,n5381 ,n6318);
    nand g7039(n4555 ,n1172 ,n4298);
    or g7040(n4140 ,n1960 ,n3848);
    nor g7041(n2234 ,n6 ,n1744);
    or g7042(n10[29] ,n4865 ,n4700);
    nand g7043(n3766 ,n7168 ,n3102);
    not g7044(n4993 ,n4994);
    nor g7045(n867 ,n709 ,n0[38]);
    nand g7046(n6818 ,n6581 ,n7096);
    nand g7047(n1159 ,n6832 ,n797);
    nor g7048(n2618 ,n0[10] ,n1963);
    nand g7049(n3789 ,n7150 ,n3015);
    nand g7050(n9[84] ,n5689 ,n6020);
    nand g7051(n3213 ,n1197 ,n2106);
    nand g7052(n5375 ,n4259 ,n5111);
    xnor g7053(n1462 ,n0[30] ,n0[6]);
    xnor g7054(n4450 ,n3943 ,n2832);
    or g7055(n408 ,n376 ,n325);
    nand g7056(n4864 ,n4142 ,n4631);
    nand g7057(n1190 ,n6881 ,n795);
    xnor g7058(n1515 ,n1[46] ,n1[14]);
    xor g7059(n4892 ,n4212 ,n4575);
    nor g7060(n4417 ,n722 ,n4214);
    xnor g7061(n1514 ,n1[38] ,n1[6]);
    nor g7062(n4022 ,n3227 ,n3395);
    nand g7063(n4129 ,n2560 ,n3942);
    nand g7064(n2446 ,n0[34] ,n718);
    nor g7065(n4951 ,n3796 ,n4816);
    nor g7066(n2410 ,n0[73] ,n1771);
    nor g7067(n2092 ,n1956 ,n1491);
    nor g7068(n885 ,n803 ,n0[106]);
    nor g7069(n2429 ,n1[62] ,n1483);
    nor g7070(n1872 ,n0[25] ,n994);
    not g7071(n2614 ,n2613);
    or g7072(n2736 ,n2626 ,n2408);
    nor g7073(n4778 ,n0[99] ,n4394);
    xnor g7074(n2948 ,n1694 ,n1522);
    nand g7075(n7081 ,n681 ,n647);
    xnor g7076(n1392 ,n1[50] ,n2[50]);
    nor g7077(n2284 ,n6 ,n2006);
    nor g7078(n3920 ,n2463 ,n3687);
    nand g7079(n6221 ,n6151 ,n6073);
    nor g7080(n5307 ,n4970 ,n5192);
    nand g7081(n6954 ,n6754 ,n6801);
    or g7082(n1736 ,n978 ,n987);
    nand g7083(n3158 ,n2601 ,n2472);
    nand g7084(n5063 ,n6 ,n4846);
    xnor g7085(n4839 ,n4429 ,n4570);
    nand g7086(n924 ,n0[126] ,n708);
    nand g7087(n5563 ,n4690 ,n5230);
    xnor g7088(n4369 ,n3957 ,n3953);
    xnor g7089(n6936 ,n536 ,n611);
    not g7090(n4229 ,n4228);
    or g7091(n3514 ,n6825 ,n2848);
    nor g7092(n2136 ,n1961 ,n1474);
    nand g7093(n505 ,n0[123] ,n6980);
    xnor g7094(n1480 ,n1[83] ,n2[19]);
    nor g7095(n1999 ,n870 ,n927);
    xnor g7096(n1653 ,n0[41] ,n0[25]);
    nor g7097(n6391 ,n5093 ,n6383);
    nor g7098(n5316 ,n4741 ,n5178);
    nor g7099(n5999 ,n3329 ,n5901);
    nand g7100(n427 ,n374 ,n426);
    nor g7101(n5750 ,n5495 ,n5608);
    or g7102(n4742 ,n3535 ,n4565);
    nand g7103(n5009 ,n3864 ,n4753);
    nand g7104(n6775 ,n1[109] ,n7088);
    nor g7105(n5613 ,n1954 ,n5431);
    nor g7106(n4044 ,n3761 ,n3033);
    xnor g7107(n3815 ,n1[78] ,n2678);
    nand g7108(n3195 ,n2570 ,n2496);
    nor g7109(n3124 ,n1915 ,n2186);
    or g7110(n2222 ,n1959 ,n1458);
    xnor g7111(n1894 ,n1[29] ,n2[29]);
    nor g7112(n3059 ,n1810 ,n2434);
    not g7113(n5295 ,n5226);
    nor g7114(n1748 ,n0[97] ,n1226);
    nand g7115(n3930 ,n2995 ,n3595);
    nand g7116(n5828 ,n3992 ,n5614);
    nor g7117(n3342 ,n1954 ,n2945);
    xnor g7118(n1318 ,n0[77] ,n7105);
    nand g7119(n3404 ,n2056 ,n2744);
    nor g7120(n2280 ,n719 ,n1621);
    nor g7121(n5784 ,n794 ,n5596);
    nor g7122(n2311 ,n1957 ,n1636);
    xnor g7123(n4896 ,n2825 ,n4451);
    nor g7124(n6116 ,n712 ,n6067);
    nor g7125(n3867 ,n2539 ,n3721);
    nor g7126(n2634 ,n0[8] ,n721);
    xnor g7127(n96 ,n0[12] ,n7068);
    nand g7128(n6568 ,n5126 ,n6551);
    nor g7129(n5961 ,n711 ,n5936);
    nor g7130(n3579 ,n1222 ,n2854);
    nor g7131(n3978 ,n710 ,n3800);
    xnor g7132(n1651 ,n0[92] ,n4[20]);
    nand g7133(n4554 ,n1134 ,n4307);
    nand g7134(n3975 ,n0[7] ,n3491);
    nor g7135(n2194 ,n1958 ,n1603);
    or g7136(n2132 ,n1962 ,n1472);
    nand g7137(n5598 ,n4699 ,n5455);
    nor g7138(n893 ,n1[115] ,n2[51]);
    nand g7139(n649 ,n0[82] ,n622);
    xnor g7140(n2927 ,n1606 ,n1532);
    or g7141(n4868 ,n3970 ,n4639);
    nor g7142(n4602 ,n706 ,n4576);
    nand g7143(n70 ,n7066 ,n0[10]);
    not g7144(n5933 ,n5932);
    nand g7145(n4094 ,n7140 ,n3474);
    nor g7146(n2404 ,n1[117] ,n719);
    xnor g7147(n6853 ,n394 ,n417);
    xnor g7148(n6848 ,n545 ,n567);
    nor g7149(n4747 ,n4309 ,n4506);
    nor g7150(n3877 ,n787 ,n3791);
    not g7151(n2908 ,n2907);
    xnor g7152(n1683 ,n0[96] ,n4[8]);
    xnor g7153(n6195 ,n6108 ,n5973);
    nand g7154(n4760 ,n2560 ,n4443);
    nand g7155(n5682 ,n4024 ,n5510);
    nor g7156(n5444 ,n6 ,n5375);
    or g7157(n4528 ,n791 ,n4364);
    nand g7158(n5733 ,n717 ,n5580);
    nor g7159(n5232 ,n3456 ,n5189);
    nand g7160(n4052 ,n789 ,n3522);
    nand g7161(n5824 ,n5653 ,n5713);
    xnor g7162(n2917 ,n1650 ,n1618);
    nand g7163(n6819 ,n6581 ,n7095);
    xnor g7164(n1539 ,n1[40] ,n1[8]);
    nor g7165(n3516 ,n1222 ,n2798);
    nor g7166(n5669 ,n4328 ,n5450);
    nor g7167(n4185 ,n1960 ,n3821);
    nor g7168(n3061 ,n1818 ,n2271);
    nor g7169(n946 ,n0[116] ,n6);
    nand g7170(n3638 ,n1[54] ,n2985);
    nand g7171(n4077 ,n3645 ,n3639);
    nor g7172(n5398 ,n6 ,n5380);
    or g7173(n2023 ,n0[32] ,n1067);
    nand g7174(n4827 ,n1966 ,n4434);
    xnor g7175(n5569 ,n5200 ,n2697);
    nand g7176(n4825 ,n1966 ,n4446);
    nand g7177(n4253 ,n710 ,n4111);
    xnor g7178(n1900 ,n1[81] ,n2[17]);
    nand g7179(n3135 ,n1579 ,n2562);
    nor g7180(n4409 ,n715 ,n4361);
    nand g7181(n1118 ,n6929 ,n797);
    xnor g7182(n1374 ,n0[82] ,n7110);
    nor g7183(n3649 ,n799 ,n3086);
    nand g7184(n3570 ,n723 ,n2993);
    nor g7185(n5974 ,n4850 ,n5887);
    nand g7186(n5474 ,n4687 ,n5332);
    nor g7187(n5965 ,n5623 ,n5918);
    nor g7188(n2097 ,n893 ,n1961);
    xor g7189(n6830 ,n1[32] ,n0[32]);
    xnor g7190(n1509 ,n0[3] ,n1[3]);
    nand g7191(n3574 ,n794 ,n3246);
    xnor g7192(n1354 ,n0[23] ,n0[7]);
    nor g7193(n2623 ,n0[24] ,n1963);
    xnor g7194(n6934 ,n231 ,n305);
    xnor g7195(n2650 ,n1281 ,n1527);
    nand g7196(n6366 ,n3673 ,n6268);
    nor g7197(n3845 ,n3581 ,n2728);
    nand g7198(n1184 ,n6931 ,n795);
    nand g7199(n3417 ,n1953 ,n2927);
    nand g7200(n5559 ,n4832 ,n5237);
    nor g7201(n3688 ,n3153 ,n2454);
    nand g7202(n3747 ,n7154 ,n3071);
    nand g7203(n2058 ,n792 ,n1984);
    not g7204(n5770 ,n5769);
    nor g7205(n6592 ,n0[106] ,n0[74]);
    xnor g7206(n1506 ,n1[54] ,n1[22]);
    or g7207(n5695 ,n2325 ,n5530);
    nand g7208(n6330 ,n717 ,n6307);
    nor g7209(n5650 ,n6 ,n5530);
    nand g7210(n5218 ,n4955 ,n5076);
    nand g7211(n3624 ,n2432 ,n3128);
    nand g7212(n4345 ,n3587 ,n3989);
    nand g7213(n4079 ,n2478 ,n3597);
    nand g7214(n1967 ,n1082 ,n1087);
    nand g7215(n3971 ,n3584 ,n2121);
    nand g7216(n2524 ,n1099 ,n1745);
    xnor g7217(n1332 ,n6919 ,n6916);
    nand g7218(n7033 ,n6642 ,n7140);
    xnor g7219(n1510 ,n0[55] ,n4[15]);
    nand g7220(n5607 ,n5099 ,n5485);
    nor g7221(n3289 ,n1954 ,n2865);
    nand g7222(n4350 ,n3599 ,n4013);
    nor g7223(n6228 ,n3290 ,n6116);
    nor g7224(n1722 ,n1054 ,n1013);
    nand g7225(n6185 ,n5552 ,n6165);
    nor g7226(n952 ,n759 ,n0[113]);
    nor g7227(n6520 ,n5537 ,n6489);
    nor g7228(n6601 ,n0[124] ,n0[92]);
    nor g7229(n4184 ,n3498 ,n3894);
    xnor g7230(n2656 ,n1331 ,n1293);
    or g7231(n4741 ,n3534 ,n4554);
    nand g7232(n6659 ,n0[75] ,n6579);
    xnor g7233(n1400 ,n1[52] ,n2[52]);
    nor g7234(n2175 ,n1961 ,n1912);
    nand g7235(n6611 ,n0[94] ,n6580);
    nand g7236(n3733 ,n7129 ,n3051);
    nor g7237(n5902 ,n713 ,n5832);
    or g7238(n2990 ,n1[56] ,n2594);
    xnor g7239(n392 ,n6990 ,n7022);
    xnor g7240(n6928 ,n534 ,n607);
    nor g7241(n871 ,n710 ,n0[62]);
    xnor g7242(n1791 ,n0[74] ,n734);
    nor g7243(n6135 ,n6060 ,n6056);
    not g7244(n794 ,n6);
    nor g7245(n5996 ,n711 ,n5931);
    xnor g7246(n2818 ,n1250 ,n1671);
    xnor g7247(n404 ,n7002 ,n7034);
    xnor g7248(n2958 ,n1706 ,n1501);
    xor g7249(n7096 ,n0[36] ,n0[4]);
    nand g7250(n2519 ,n794 ,n1980);
    nand g7251(n2259 ,n792 ,n2004);
    nor g7252(n2615 ,n0[25] ,n721);
    nand g7253(n1212 ,n0[125] ,n709);
    nor g7254(n1972 ,n1074 ,n1083);
    nand g7255(n6005 ,n5554 ,n5874);
    nor g7256(n3577 ,n2325 ,n3247);
    not g7257(n4917 ,n4916);
    nand g7258(n6408 ,n6369 ,n6145);
    not g7259(n842 ,n0[62]);
    nor g7260(n2055 ,n1962 ,n1921);
    nand g7261(n4296 ,n2570 ,n4085);
    or g7262(n5505 ,n2209 ,n5383);
    xnor g7263(n225 ,n1[52] ,n0[52]);
    nand g7264(n6771 ,n1[125] ,n7088);
    or g7265(n6435 ,n6381 ,n6283);
    nand g7266(n271 ,n215 ,n270);
    nand g7267(n2571 ,n0[30] ,n1964);
    nand g7268(n438 ,n324 ,n437);
    nor g7269(n3932 ,n722 ,n3493);
    xnor g7270(n6563 ,n6509 ,n1287);
    not g7271(n5010 ,n5009);
    nor g7272(n2621 ,n0[22] ,n1963);
    or g7273(n179 ,n0[37] ,n1[37]);
    nor g7274(n4150 ,n1961 ,n3820);
    nand g7275(n5084 ,n4243 ,n4936);
    nand g7276(n523 ,n0[121] ,n6978);
    nor g7277(n1107 ,n752 ,n0[56]);
    xnor g7278(n2847 ,n1285 ,n1703);
    or g7279(n5684 ,n3911 ,n5548);
    xnor g7280(n1718 ,n6831 ,n6828);
    nand g7281(n155 ,n68 ,n154);
    nand g7282(n525 ,n0[99] ,n6956);
    nor g7283(n3419 ,n1954 ,n2927);
    xnor g7284(n1288 ,n0[73] ,n7101);
    nor g7285(n6570 ,n4945 ,n6558);
    nor g7286(n2250 ,n1957 ,n1601);
    nor g7287(n4293 ,n817 ,n4017);
    xnor g7288(n2893 ,n1255 ,n1351);
    or g7289(n4702 ,n1965 ,n4463);
    nor g7290(n6588 ,n0[102] ,n0[70]);
    nand g7291(n5369 ,n3805 ,n5151);
    xnor g7292(n1619 ,n0[75] ,n1[75]);
    or g7293(n6065 ,n5632 ,n5975);
    xnor g7294(n1439 ,n0[84] ,n1[84]);
    nor g7295(n2060 ,n1777 ,n1779);
    xnor g7296(n1313 ,n0[76] ,n7104);
    nand g7297(n6518 ,n6479 ,n6493);
    nand g7298(n2017 ,n723 ,n1048);
    nand g7299(n9[12] ,n6094 ,n6178);
    or g7300(n6485 ,n6437 ,n6345);
    or g7301(n2072 ,n1961 ,n1894);
    or g7302(n30 ,n7077 ,n0[21]);
    nand g7303(n465 ,n347 ,n464);
    nand g7304(n3177 ,n2562 ,n2493);
    or g7305(n483 ,n0[101] ,n6958);
    nor g7306(n4530 ,n722 ,n4220);
    nand g7307(n6641 ,n1[68] ,n6579);
    or g7308(n2988 ,n2635 ,n2364);
    or g7309(n493 ,n0[113] ,n6970);
    nor g7310(n1776 ,n0[73] ,n1026);
    or g7311(n5310 ,n3416 ,n5179);
    not g7312(n5162 ,n5161);
    nor g7313(n3165 ,n1878 ,n2565);
    not g7314(n5073 ,n5072);
    nand g7315(n9[10] ,n6179 ,n6291);
    xnor g7316(n5942 ,n5845 ,n1523);
    nor g7317(n3529 ,n6825 ,n2839);
endmodule
