module top (n0, n1, n7, n8, n9, n2, n3, n4, n5, n14, n15, n6, n16, n17, n10, n11, n12, n13);
    input n0, n1, n2, n3, n4, n5, n6;
    input [6:0] n7;
    input [7:0] n8;
    output [7:0] n9, n10, n11, n12, n13;
    output n14, n15, n16, n17;
    wire n0, n1, n2, n3, n4, n5, n6;
    wire [6:0] n7;
    wire [7:0] n8;
    wire [7:0] n9, n10, n11, n12, n13;
    wire n14, n15, n16, n17;
    wire [2:0] n18;
    wire [4:0] n19;
    wire [4:0] n20;
    wire [3:0] n21;
    wire [15:0] n22;
    wire [7:0] n23;
    wire [7:0] n24;
    wire [7:0] n25;
    wire [7:0] n26;
    wire [7:0] n27;
    wire [7:0] n28;
    wire [7:0] n29;
    wire [7:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [7:0] n36;
    wire [7:0] n37;
    wire [7:0] n38;
    wire [3:0] n39;
    wire [3:0] n40;
    wire [7:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [7:0] n44;
    wire [7:0] n45;
    wire [7:0] n46;
    wire [7:0] n47;
    wire [7:0] n48;
    wire [7:0] n49;
    wire [7:0] n50;
    wire [7:0] n51;
    wire [7:0] n52;
    wire [7:0] n53;
    wire [7:0] n54;
    wire [7:0] n55;
    wire [7:0] n56;
    wire [7:0] n57;
    wire [3:0] n58;
    wire [3:0] n59;
    wire [7:0] n60;
    wire n61, n62, n63, n64, n65, n66, n67, n68;
    wire n69, n70, n71, n72, n73, n74, n75, n76;
    wire n77, n78, n79, n80, n81, n82, n83, n84;
    wire n85, n86, n87, n88, n89, n90, n91, n92;
    wire n93, n94, n95, n96, n97, n98, n99, n100;
    wire n101, n102, n103, n104, n105, n106, n107, n108;
    wire n109, n110, n111, n112, n113, n114, n115, n116;
    wire n117, n118, n119, n120, n121, n122, n123, n124;
    wire n125, n126, n127, n128, n129, n130, n131, n132;
    wire n133, n134, n135, n136, n137, n138, n139, n140;
    wire n141, n142, n143, n144, n145, n146, n147, n148;
    wire n149, n150, n151, n152, n153, n154, n155, n156;
    wire n157, n158, n159, n160, n161, n162, n163, n164;
    wire n165, n166, n167, n168, n169, n170, n171, n172;
    wire n173, n174, n175, n176, n177, n178, n179, n180;
    wire n181, n182, n183, n184, n185, n186, n187, n188;
    wire n189, n190, n191, n192, n193, n194, n195, n196;
    wire n197, n198, n199, n200, n201, n202, n203, n204;
    wire n205, n206, n207, n208, n209, n210, n211, n212;
    wire n213, n214, n215, n216, n217, n218, n219, n220;
    wire n221, n222, n223, n224, n225, n226, n227, n228;
    wire n229, n230, n231, n232, n233, n234, n235, n236;
    wire n237, n238, n239, n240, n241, n242, n243, n244;
    wire n245, n246, n247, n248, n249, n250, n251, n252;
    wire n253, n254, n255, n256, n257, n258, n259, n260;
    wire n261, n262, n263, n264, n265, n266, n267, n268;
    wire n269, n270, n271, n272, n273, n274, n275, n276;
    wire n277, n278, n279, n280, n281, n282, n283, n284;
    wire n285, n286, n287, n288, n289, n290, n291, n292;
    wire n293, n294, n295, n296, n297, n298, n299, n300;
    wire n301, n302, n303, n304, n305, n306, n307, n308;
    wire n309, n310, n311, n312, n313, n314, n315, n316;
    wire n317, n318, n319, n320, n321, n322, n323, n324;
    wire n325, n326, n327, n328, n329, n330, n331, n332;
    wire n333, n334, n335, n336, n337, n338, n339, n340;
    wire n341, n342, n343, n344, n345, n346, n347, n348;
    wire n349, n350, n351, n352, n353, n354, n355, n356;
    wire n357, n358, n359, n360, n361, n362, n363, n364;
    wire n365, n366, n367, n368, n369, n370, n371, n372;
    wire n373, n374, n375, n376, n377, n378, n379, n380;
    wire n381, n382, n383, n384, n385, n386, n387, n388;
    wire n389, n390, n391, n392, n393, n394, n395, n396;
    wire n397, n398, n399, n400, n401, n402, n403, n404;
    wire n405, n406, n407, n408, n409, n410, n411, n412;
    wire n413, n414, n415, n416, n417, n418, n419, n420;
    wire n421, n422, n423, n424, n425, n426, n427, n428;
    wire n429, n430, n431, n432, n433, n434, n435, n436;
    wire n437, n438, n439, n440, n441, n442, n443, n444;
    wire n445, n446, n447, n448, n449, n450, n451, n452;
    wire n453, n454, n455, n456, n457, n458, n459, n460;
    wire n461, n462, n463, n464, n465, n466, n467, n468;
    wire n469, n470, n471, n472, n473, n474, n475, n476;
    wire n477, n478, n479, n480, n481, n482, n483, n484;
    wire n485, n486, n487, n488, n489, n490, n491, n492;
    wire n493, n494, n495, n496, n497, n498, n499, n500;
    wire n501, n502, n503, n504, n505, n506, n507, n508;
    wire n509, n510, n511, n512, n513, n514, n515, n516;
    wire n517, n518, n519, n520, n521, n522, n523, n524;
    wire n525, n526, n527, n528, n529, n530, n531, n532;
    wire n533, n534, n535, n536, n537, n538, n539, n540;
    wire n541, n542, n543, n544, n545, n546, n547, n548;
    wire n549, n550, n551, n552, n553, n554, n555, n556;
    wire n557, n558, n559, n560, n561, n562, n563, n564;
    wire n565, n566, n567, n568, n569, n570, n571, n572;
    wire n573, n574, n575, n576, n577, n578, n579, n580;
    wire n581, n582, n583, n584, n585, n586, n587, n588;
    wire n589, n590, n591, n592, n593, n594, n595, n596;
    wire n597, n598, n599, n600, n601, n602, n603, n604;
    wire n605, n606, n607, n608, n609, n610, n611, n612;
    wire n613, n614, n615, n616, n617, n618, n619, n620;
    wire n621, n622, n623, n624, n625, n626, n627, n628;
    wire n629, n630, n631, n632, n633, n634, n635, n636;
    wire n637, n638, n639, n640, n641, n642, n643, n644;
    wire n645, n646, n647, n648, n649, n650, n651, n652;
    wire n653, n654, n655, n656, n657, n658, n659, n660;
    wire n661, n662, n663, n664, n665, n666, n667, n668;
    wire n669, n670, n671, n672, n673, n674, n675, n676;
    wire n677, n678, n679, n680, n681, n682, n683, n684;
    wire n685, n686, n687, n688, n689, n690, n691, n692;
    wire n693, n694, n695, n696, n697, n698, n699, n700;
    wire n701, n702, n703, n704, n705, n706, n707, n708;
    wire n709, n710, n711, n712, n713, n714, n715, n716;
    wire n717, n718, n719, n720, n721, n722, n723, n724;
    wire n725, n726, n727, n728, n729, n730, n731, n732;
    wire n733, n734, n735, n736, n737, n738, n739, n740;
    wire n741, n742, n743, n744, n745, n746, n747, n748;
    wire n749, n750, n751, n752, n753, n754, n755, n756;
    wire n757, n758, n759, n760, n761, n762, n763, n764;
    wire n765, n766, n767, n768, n769, n770, n771, n772;
    wire n773, n774, n775, n776, n777, n778, n779, n780;
    wire n781, n782, n783, n784, n785, n786, n787, n788;
    wire n789, n790, n791, n792, n793, n794, n795, n796;
    wire n797, n798, n799, n800, n801, n802, n803, n804;
    wire n805, n806, n807, n808, n809, n810, n811, n812;
    wire n813, n814, n815, n816, n817, n818, n819, n820;
    wire n821, n822, n823, n824, n825, n826, n827, n828;
    wire n829, n830, n831, n832, n833, n834, n835, n836;
    wire n837, n838, n839, n840, n841, n842, n843, n844;
    wire n845, n846, n847, n848, n849, n850, n851, n852;
    wire n853, n854, n855, n856, n857, n858, n859, n860;
    wire n861, n862, n863, n864, n865, n866, n867, n868;
    wire n869, n870, n871, n872, n873, n874, n875, n876;
    wire n877, n878, n879, n880, n881, n882, n883, n884;
    wire n885, n886, n887, n888, n889, n890, n891, n892;
    wire n893, n894, n895, n896, n897, n898, n899, n900;
    wire n901, n902, n903, n904, n905, n906, n907, n908;
    wire n909, n910, n911, n912, n913, n914, n915, n916;
    wire n917, n918, n919, n920, n921, n922, n923, n924;
    wire n925, n926, n927, n928, n929, n930, n931, n932;
    wire n933, n934, n935, n936, n937, n938, n939, n940;
    wire n941, n942, n943, n944, n945, n946, n947, n948;
    wire n949, n950, n951, n952, n953, n954, n955, n956;
    wire n957, n958, n959, n960, n961, n962, n963, n964;
    wire n965, n966, n967, n968, n969, n970, n971, n972;
    wire n973, n974, n975, n976, n977, n978, n979, n980;
    wire n981, n982, n983, n984, n985, n986, n987, n988;
    wire n989, n990, n991, n992, n993, n994, n995, n996;
    wire n997, n998, n999, n1000, n1001, n1002, n1003, n1004;
    wire n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012;
    wire n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
    wire n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
    wire n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
    wire n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044;
    wire n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
    wire n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060;
    wire n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068;
    wire n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076;
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084;
    wire n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092;
    wire n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100;
    wire n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108;
    wire n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116;
    wire n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124;
    wire n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132;
    wire n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140;
    wire n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148;
    wire n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156;
    wire n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164;
    wire n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172;
    wire n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180;
    wire n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188;
    wire n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196;
    wire n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204;
    wire n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
    wire n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220;
    wire n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228;
    wire n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236;
    wire n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244;
    wire n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252;
    wire n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260;
    wire n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268;
    wire n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276;
    wire n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284;
    wire n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292;
    wire n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300;
    wire n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308;
    wire n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;
    wire n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;
    wire n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332;
    wire n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340;
    wire n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348;
    wire n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356;
    wire n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364;
    wire n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372;
    wire n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380;
    wire n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388;
    wire n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;
    wire n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404;
    wire n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412;
    wire n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;
    wire n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428;
    wire n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436;
    wire n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444;
    wire n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452;
    wire n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;
    wire n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468;
    wire n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476;
    wire n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
    wire n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492;
    wire n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500;
    wire n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508;
    wire n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516;
    wire n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524;
    wire n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532;
    wire n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540;
    wire n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548;
    wire n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556;
    wire n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564;
    wire n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572;
    wire n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580;
    wire n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588;
    wire n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596;
    wire n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604;
    wire n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612;
    wire n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620;
    wire n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628;
    wire n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636;
    wire n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644;
    wire n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652;
    wire n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660;
    wire n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668;
    wire n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676;
    wire n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684;
    wire n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692;
    wire n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700;
    wire n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708;
    wire n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716;
    wire n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724;
    wire n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732;
    wire n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740;
    wire n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748;
    wire n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756;
    wire n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764;
    wire n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772;
    wire n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780;
    wire n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788;
    wire n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796;
    wire n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804;
    wire n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812;
    wire n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820;
    wire n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828;
    wire n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836;
    wire n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844;
    wire n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852;
    wire n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860;
    wire n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868;
    wire n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876;
    wire n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884;
    wire n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892;
    wire n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900;
    wire n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908;
    wire n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916;
    wire n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924;
    wire n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932;
    wire n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940;
    wire n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948;
    wire n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956;
    wire n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964;
    wire n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972;
    wire n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980;
    wire n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988;
    wire n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996;
    wire n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004;
    wire n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012;
    wire n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020;
    wire n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028;
    wire n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036;
    wire n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044;
    wire n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052;
    wire n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060;
    wire n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068;
    wire n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076;
    wire n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084;
    wire n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092;
    wire n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100;
    wire n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108;
    wire n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116;
    wire n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124;
    wire n2125, n2126, n2127, n2128, n2129, n2130;
    nor g0(n1913 ,n1438 ,n1704);
    not g1(n97 ,n22[4]);
    nand g2(n1049 ,n2115 ,n868);
    not g3(n197 ,n196);
    nand g4(n582 ,n8[1] ,n456);
    nand g5(n1450 ,n41[4] ,n1307);
    nand g6(n292 ,n22[13] ,n245);
    nor g7(n1439 ,n41[0] ,n1315);
    nand g8(n1371 ,n657 ,n1230);
    not g9(n2080 ,n18[1]);
    nor g10(n231 ,n162 ,n59[1]);
    nand g11(n1642 ,n56[4] ,n1341);
    nand g12(n1193 ,n578 ,n855);
    nand g13(n1797 ,n31[6] ,n1555);
    nor g14(n106 ,n97 ,n105);
    nor g15(n771 ,n54[0] ,n600);
    nand g16(n1857 ,n1646 ,n1616);
    nor g17(n1704 ,n36[0] ,n1546);
    nand g18(n681 ,n26[5] ,n420);
    nor g19(n761 ,n155 ,n425);
    nand g20(n1221 ,n58[2] ,n1079);
    dff g21(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1051), .Q(n54[7]));
    nand g22(n317 ,n304 ,n313);
    nand g23(n1500 ,n41[7] ,n1316);
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1813), .Q(n26[4]));
    nand g25(n1220 ,n58[1] ,n1079);
    nand g26(n1849 ,n1638 ,n1676);
    nand g27(n1166 ,n57[5] ,n871);
    nand g28(n534 ,n8[7] ,n395);
    nand g29(n1962 ,n1424 ,n1738);
    not g30(n150 ,n42[4]);
    nand g31(n1604 ,n46[2] ,n1340);
    nand g32(n1517 ,n45[7] ,n1386);
    nand g33(n1367 ,n381 ,n1202);
    nand g34(n567 ,n8[4] ,n450);
    nand g35(n1350 ,n736 ,n1224);
    nand g36(n1148 ,n549 ,n786);
    not g37(n1386 ,n1385);
    nand g38(n790 ,n54[6] ,n601);
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n437), .Q(n22[5]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1169), .Q(n53[6]));
    nand g41(n741 ,n37[4] ,n415);
    nand g42(n1815 ,n1284 ,n1518);
    nand g43(n2009 ,n1481 ,n1773);
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1102), .Q(n49[4]));
    nand g45(n1593 ,n45[0] ,n1386);
    nand g46(n1839 ,n1684 ,n1629);
    nand g47(n2024 ,n1435 ,n1760);
    nor g48(n309 ,n140 ,n272);
    nand g49(n1468 ,n41[5] ,n1310);
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1600), .Q(n19[1]));
    nand g51(n835 ,n47[5] ,n617);
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1815), .Q(n26[2]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1212), .Q(n21[2]));
    nor g54(n305 ,n148 ,n276);
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1970), .Q(n24[7]));
    nand g56(n1066 ,n60[3] ,n865);
    nand g57(n1108 ,n532 ,n828);
    nand g58(n1134 ,n558 ,n850);
    nand g59(n822 ,n49[5] ,n603);
    nand g60(n901 ,n56[4] ,n595);
    nand g61(n1768 ,n37[2] ,n1543);
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1991), .Q(n31[6]));
    nand g63(n339 ,n39[0] ,n311);
    or g64(n1396 ,n921 ,n1370);
    not g65(n99 ,n22[12]);
    nand g66(n662 ,n24[6] ,n418);
    not g67(n1266 ,n1199);
    nor g68(n1895 ,n1425 ,n1699);
    nand g69(n1613 ,n55[4] ,n1382);
    nor g70(n1438 ,n41[0] ,n1323);
    nand g71(n2120 ,n2073 ,n2074);
    nand g72(n1829 ,n1670 ,n1621);
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n210), .Q(n10[7]));
    nand g74(n1837 ,n1667 ,n1686);
    nand g75(n287 ,n22[5] ,n245);
    nand g76(n2011 ,n1466 ,n1740);
    nand g77(n1431 ,n41[1] ,n1311);
    or g78(n177 ,n154 ,n3);
    nand g79(n1061 ,n568 ,n797);
    nand g80(n1056 ,n522 ,n800);
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n20[4]));
    nand g82(n1207 ,n590 ,n1178);
    nand g83(n269 ,n141 ,n255);
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1109), .Q(n48[3]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1208), .Q(n57[1]));
    nand g86(n1165 ,n20[1] ,n873);
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1238), .Q(n57[0]));
    nor g88(n395 ,n261 ,n385);
    nand g89(n424 ,n1 ,n364);
    nand g90(n1562 ,n49[3] ,n1334);
    nor g91(n2109 ,n121 ,n123);
    nand g92(n848 ,n45[5] ,n607);
    nand g93(n203 ,n22[2] ,n22[3]);
    xnor g94(n2089 ,n58[2] ,n94);
    nor g95(n1227 ,n1007 ,n1006);
    not g96(n428 ,n389);
    nor g97(n167 ,n22[8] ,n22[9]);
    nand g98(n1376 ,n1025 ,n1235);
    nor g99(n107 ,n22[5] ,n106);
    nand g100(n1675 ,n46[4] ,n1340);
    nand g101(n1356 ,n1035 ,n1196);
    nor g102(n759 ,n161 ,n460);
    nand g103(n949 ,n721 ,n653);
    nand g104(n657 ,n30[3] ,n417);
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2016), .Q(n37[2]));
    nand g106(n1982 ,n1492 ,n1788);
    nand g107(n791 ,n54[5] ,n601);
    nand g108(n1632 ,n56[5] ,n1341);
    nand g109(n831 ,n48[1] ,n605);
    nand g110(n696 ,n37[2] ,n415);
    not g111(n1085 ,n1084);
    nand g112(n738 ,n25[2] ,n459);
    nand g113(n640 ,n34[3] ,n416);
    nand g114(n2062 ,n1940 ,n2056);
    not g115(n111 ,n110);
    nand g116(n796 ,n53[5] ,n615);
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n996), .Q(n45[0]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1168), .Q(n56[4]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1884), .Q(n34[1]));
    nor g120(n627 ,n327 ,n452);
    nand g121(n1603 ,n43[7] ,n1384);
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1269), .Q(n15));
    not g123(n1340 ,n1339);
    nand g124(n1764 ,n37[6] ,n1543);
    nand g125(n1092 ,n477 ,n814);
    not g126(n154 ,n18[2]);
    nand g127(n891 ,n51[2] ,n613);
    nand g128(n344 ,n2126 ,n302);
    not g129(n871 ,n870);
    nand g130(n1771 ,n1522 ,n1693);
    nand g131(n1574 ,n34[7] ,n1332);
    nor g132(n1302 ,n218 ,n1263);
    nand g133(n795 ,n53[6] ,n615);
    nor g134(n1712 ,n933 ,n1401);
    xnor g135(n2100 ,n22[4] ,n105);
    nand g136(n912 ,n651 ,n692);
    nand g137(n1616 ,n44[3] ,n1381);
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1193), .Q(n44[3]));
    nand g139(n280 ,n22[10] ,n245);
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1152), .Q(n42[5]));
    nand g141(n1760 ,n23[3] ,n1535);
    nand g142(n1198 ,n344 ,n1164);
    nand g143(n716 ,n33[7] ,n422);
    nand g144(n1584 ,n34[3] ,n1332);
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n20[3]));
    nand g146(n1960 ,n1423 ,n1739);
    nand g147(n1156 ,n471 ,n880);
    nand g148(n1114 ,n557 ,n835);
    not g149(n390 ,n391);
    nand g150(n913 ,n337 ,n742);
    nand g151(n1352 ,n60[5] ,n1252);
    nand g152(n1807 ,n1275 ,n1506);
    nand g153(n1650 ,n56[2] ,n1341);
    nand g154(n911 ,n55[1] ,n619);
    nand g155(n1140 ,n544 ,n911);
    nor g156(n473 ,n8[0] ,n394);
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n993), .Q(n47[0]));
    nor g158(n1289 ,n41[0] ,n1250);
    nand g159(n1360 ,n60[6] ,n1252);
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1268), .Q(n41[0]));
    buf g161(n13[4], n10[6]);
    nand g162(n433 ,n284 ,n371);
    or g163(n1407 ,n966 ,n1350);
    nand g164(n1037 ,n40[0] ,n872);
    nand g165(n1687 ,n51[6] ,n1342);
    not g166(n95 ,n94);
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1192), .Q(n55[2]));
    nand g168(n1129 ,n593 ,n849);
    nand g169(n1115 ,n536 ,n836);
    nand g170(n864 ,n1 ,n625);
    nand g171(n1039 ,n762 ,n882);
    nor g172(n296 ,n140 ,n266);
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2058), .Q(n60[3]));
    nand g174(n541 ,n8[3] ,n395);
    nand g175(n1462 ,n41[4] ,n1314);
    nor g176(n1912 ,n1855 ,n1854);
    buf g177(n13[2], n10[0]);
    nand g178(n248 ,n158 ,n231);
    nand g179(n1282 ,n41[4] ,n1244);
    nand g180(n1447 ,n41[1] ,n1303);
    nand g181(n824 ,n49[2] ,n603);
    nand g182(n527 ,n8[3] ,n409);
    nor g183(n1267 ,n41[0] ,n1247);
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1018), .Q(n56[0]));
    nand g185(n1413 ,n41[6] ,n1319);
    nand g186(n717 ,n36[7] ,n458);
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1134), .Q(n45[1]));
    nor g188(n605 ,n140 ,n407);
    nand g189(n1671 ,n54[2] ,n1383);
    nand g190(n1831 ,n1672 ,n1625);
    nand g191(n2013 ,n1479 ,n1772);
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1073), .Q(n51[7]));
    not g193(n327 ,n328);
    nand g194(n530 ,n8[7] ,n401);
    nand g195(n224 ,n11[1] ,n1);
    nand g196(n1210 ,n427 ,n1158);
    nand g197(n1195 ,n788 ,n1154);
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2025), .Q(n23[4]));
    nand g199(n1731 ,n28[2] ,n1549);
    nor g200(n240 ,n204 ,n209);
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2027), .Q(n23[6]));
    nor g202(n496 ,n8[0] ,n446);
    not g203(n91 ,n90);
    nand g204(n1868 ,n1656 ,n1561);
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1997), .Q(n58[3]));
    nand g206(n1793 ,n32[3] ,n1553);
    not g207(n1319 ,n1320);
    nand g208(n1859 ,n1565 ,n1649);
    nand g209(n477 ,n8[7] ,n399);
    nor g210(n426 ,n18[0] ,n348);
    nand g211(n1643 ,n48[3] ,n1335);
    nor g212(n1001 ,n490 ,n773);
    nor g213(n465 ,n8[0] ,n404);
    or g214(n209 ,n156 ,n21[3]);
    not g215(n1549 ,n1548);
    nand g216(n518 ,n8[7] ,n456);
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1961), .Q(n27[3]));
    nand g218(n88 ,n59[2] ,n87);
    nand g219(n2007 ,n1500 ,n1775);
    nand g220(n580 ,n8[1] ,n447);
    nand g221(n1571 ,n42[1] ,n1387);
    nand g222(n246 ,n155 ,n182);
    nand g223(n1977 ,n1488 ,n1785);
    nand g224(n1284 ,n41[2] ,n1244);
    nand g225(n1293 ,n41[7] ,n1246);
    nand g226(n202 ,n22[0] ,n149);
    nand g227(n299 ,n147 ,n268);
    buf g228(n11[4], 1'b0);
    not g229(n410 ,n411);
    or g230(n1000 ,n929 ,n920);
    not g231(n147 ,n21[1]);
    nand g232(n1128 ,n542 ,n909);
    nor g233(n328 ,n140 ,n314);
    nor g234(n1441 ,n41[0] ,n1301);
    not g235(n1535 ,n1534);
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1191), .Q(n49[2]));
    nand g237(n2037 ,n1622 ,n1900);
    nand g238(n2018 ,n1484 ,n1765);
    nor g239(n997 ,n976 ,n975);
    nand g240(n1525 ,n47[5] ,n1338);
    nand g241(n445 ,n289 ,n376);
    or g242(n1014 ,n932 ,n974);
    nand g243(n757 ,n26[2] ,n420);
    nor g244(n1224 ,n992 ,n1000);
    nand g245(n1792 ,n32[4] ,n1553);
    xnor g246(n2103 ,n22[7] ,n110);
    nor g247(n464 ,n8[0] ,n396);
    nand g248(n1212 ,n784 ,n1138);
    nand g249(n643 ,n24[0] ,n418);
    nand g250(n238 ,n167 ,n170);
    nand g251(n1975 ,n1430 ,n1753);
    nand g252(n802 ,n52[6] ,n597);
    nand g253(n1669 ,n52[0] ,n1333);
    nor g254(n462 ,n235 ,n424);
    nand g255(n336 ,n9[4] ,n311);
    dff g256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1052), .Q(n54[6]));
    nand g257(n1640 ,n1066 ,n1351);
    nand g258(n1548 ,n1 ,n1320);
    nand g259(n306 ,n9[0] ,n275);
    nand g260(n1566 ,n47[2] ,n1338);
    dff g261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1115), .Q(n47[4]));
    nor g262(n1926 ,n1410 ,n1708);
    nand g263(n1733 ,n27[7] ,n1551);
    or g264(n1005 ,n939 ,n937);
    nand g265(n1370 ,n751 ,n1229);
    not g266(n131 ,n130);
    nand g267(n1588 ,n34[1] ,n1332);
    nand g268(n934 ,n637 ,n670);
    nor g269(n1711 ,n922 ,n1396);
    nor g270(n2036 ,n1923 ,n1922);
    nand g271(n1809 ,n1276 ,n1507);
    nand g272(n1318 ,n187 ,n1258);
    nand g273(n1232 ,n41[1] ,n1077);
    nor g274(n1015 ,n140 ,n780);
    nand g275(n588 ,n8[5] ,n409);
    nand g276(n529 ,n8[1] ,n409);
    nand g277(n289 ,n22[7] ,n245);
    nor g278(n1019 ,n501 ,n779);
    nand g279(n1610 ,n30[7] ,n1330);
    nand g280(n1294 ,n41[6] ,n1251);
    dff g281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n40[2]));
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1894), .Q(n27[0]));
    nand g283(n875 ,n192 ,n466);
    nand g284(n1736 ,n27[4] ,n1551);
    nand g285(n1869 ,n1657 ,n1615);
    nand g286(n826 ,n48[6] ,n605);
    nand g287(n733 ,n29[4] ,n423);
    xnor g288(n2102 ,n22[6] ,n108);
    dff g289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1377), .Q(n41[5]));
    nand g290(n1526 ,n43[5] ,n1384);
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1978), .Q(n58[2]));
    or g292(n264 ,n238 ,n239);
    nand g293(n1559 ,n42[3] ,n1387);
    nor g294(n1258 ,n40[1] ,n1085);
    nor g295(n1938 ,n1608 ,n1851);
    not g296(n160 ,n58[1]);
    nand g297(n2004 ,n1494 ,n1777);
    nand g298(n378 ,n2098 ,n326);
    nand g299(n2034 ,n1916 ,n1915);
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1041), .Q(n59[2]));
    nand g301(n661 ,n26[6] ,n420);
    not g302(n1315 ,n1316);
    nand g303(n633 ,n26[1] ,n420);
    nand g304(n250 ,n157 ,n195);
    nor g305(n1338 ,n184 ,n1259);
    nand g306(n1181 ,n507 ,n898);
    nand g307(n752 ,n23[0] ,n419);
    nand g308(n366 ,n14 ,n334);
    nand g309(n1274 ,n41[4] ,n1248);
    nand g310(n1374 ,n1027 ,n1233);
    nand g311(n608 ,n1 ,n404);
    nand g312(n1479 ,n41[4] ,n1324);
    nand g313(n1167 ,n20[0] ,n873);
    nand g314(n598 ,n1 ,n410);
    nand g315(n1959 ,n1421 ,n1736);
    nand g316(n1368 ,n647 ,n1227);
    dff g317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1097), .Q(n50[2]));
    nand g318(n1565 ,n43[2] ,n1384);
    nand g319(n1753 ,n24[2] ,n1557);
    nand g320(n1954 ,n1417 ,n1731);
    nand g321(n290 ,n22[3] ,n245);
    nor g322(n1903 ,n1836 ,n1837);
    not g323(n1313 ,n1314);
    nand g324(n832 ,n47[7] ,n617);
    not g325(n257 ,n256);
    nand g326(n1832 ,n1690 ,n1601);
    nor g327(n615 ,n140 ,n456);
    dff g328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1149), .Q(n43[1]));
    nand g329(n1089 ,n579 ,n812);
    or g330(n1924 ,n1887 ,n1886);
    nor g331(n1915 ,n1860 ,n1859);
    not g332(n183 ,n184);
    nand g333(n1473 ,n41[6] ,n1316);
    nand g334(n737 ,n36[4] ,n458);
    nand g335(n495 ,n8[2] ,n391);
    nand g336(n512 ,n8[2] ,n399);
    nand g337(n522 ,n8[3] ,n401);
    nand g338(n1836 ,n1628 ,n1668);
    nor g339(n865 ,n193 ,n626);
    nand g340(n727 ,n29[6] ,n423);
    nand g341(n1625 ,n44[6] ,n1381);
    nand g342(n261 ,n59[1] ,n194);
    nand g343(n1035 ,n40[1] ,n872);
    nand g344(n675 ,n34[2] ,n416);
    nand g345(n1217 ,n1037 ,n1085);
    nand g346(n483 ,n8[6] ,n405);
    nor g347(n769 ,n46[0] ,n608);
    nand g348(n1052 ,n535 ,n790);
    nand g349(n1759 ,n23[4] ,n1535);
    nand g350(n1806 ,n1274 ,n1505);
    nand g351(n486 ,n8[2] ,n405);
    or g352(n1401 ,n931 ,n1369);
    nand g353(n282 ,n22[6] ,n245);
    dff g354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1143), .Q(n43[7]));
    nand g355(n117 ,n22[10] ,n116);
    nand g356(n1679 ,n50[5] ,n1337);
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1217), .Q(n40[0]));
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1807), .Q(n30[3]));
    or g359(n258 ,n214 ,n182);
    nand g360(n260 ,n59[2] ,n231);
    nand g361(n1503 ,n30[5] ,n1330);
    dff g362(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1988), .Q(n32[2]));
    dff g363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1116), .Q(n47[3]));
    dff g364(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1967), .Q(n25[4]));
    nand g365(n1144 ,n546 ,n859);
    nand g366(n1296 ,n41[4] ,n1251);
    nand g367(n1655 ,n52[2] ,n1333);
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1965), .Q(n25[3]));
    nand g369(n1595 ,n49[6] ,n1334);
    nand g370(n1063 ,n564 ,n799);
    buf g371(n12[3], 1'b0);
    nand g372(n895 ,n2082 ,n627);
    nor g373(n1703 ,n37[0] ,n1542);
    dff g374(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1882), .Q(n34[2]));
    nand g375(n438 ,n293 ,n356);
    dff g376(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1944), .Q(n29[5]));
    nor g377(n405 ,n250 ,n359);
    nand g378(n672 ,n24[5] ,n418);
    nor g379(n459 ,n188 ,n363);
    nand g380(n939 ,n709 ,n643);
    not g381(n609 ,n608);
    nand g382(n108 ,n22[5] ,n106);
    nand g383(n663 ,n27[0] ,n412);
    nand g384(n1627 ,n56[6] ,n1341);
    nand g385(n1023 ,n41[5] ,n867);
    nand g386(n1164 ,n20[2] ,n873);
    nand g387(n1133 ,n543 ,n897);
    or g388(n1013 ,n977 ,n979);
    nand g389(n762 ,n353 ,n388);
    dff g390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1596), .Q(n19[4]));
    nand g391(n1349 ,n1167 ,n1240);
    nand g392(n1950 ,n1413 ,n1726);
    nand g393(n1331 ,n1 ,n1247);
    nor g394(n1709 ,n31[0] ,n1554);
    dff g395(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1211), .Q(n57[4]));
    nand g396(n1662 ,n48[0] ,n1335);
    nand g397(n538 ,n8[2] ,n447);
    nand g398(n436 ,n283 ,n378);
    xnor g399(n2111 ,n22[15] ,n124);
    dff g400(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n441), .Q(n22[15]));
    dff g401(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1358), .Q(n19[0]));
    nand g402(n1272 ,n41[6] ,n1248);
    not g403(n127 ,n126);
    dff g404(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1356), .Q(n40[1]));
    not g405(n400 ,n401);
    nand g406(n1372 ,n1022 ,n1231);
    nand g407(n1639 ,n54[6] ,n1383);
    nand g408(n920 ,n739 ,n672);
    nand g409(n1878 ,n1279 ,n1580);
    nand g410(n2125 ,n62 ,n61);
    nand g411(n1434 ,n41[4] ,n1317);
    dff g412(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1820), .Q(n38[5]));
    dff g413(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n980), .Q(n52[0]));
    dff g414(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1373), .Q(n41[1]));
    not g415(n225 ,n224);
    nand g416(n468 ,n427 ,n387);
    nor g417(n765 ,n50[0] ,n620);
    dff g418(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1698), .Q(n26[0]));
    or g419(n985 ,n967 ,n956);
    nand g420(n1042 ,n351 ,n895);
    nand g421(n1882 ,n1288 ,n1577);
    nand g422(n1778 ,n35[5] ,n1541);
    nand g423(n363 ,n39[1] ,n331);
    not g424(n109 ,n108);
    nand g425(n726 ,n33[6] ,n422);
    nand g426(n1729 ,n28[4] ,n1549);
    dff g427(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1124), .Q(n46[2]));
    nand g428(n594 ,n1 ,n390);
    not g429(n221 ,n220);
    nand g430(n1160 ,n319 ,n884);
    nor g431(n873 ,n310 ,n625);
    nand g432(n1670 ,n57[7] ,n1380);
    nand g433(n1788 ,n33[1] ,n1545);
    nand g434(n979 ,n676 ,n756);
    nand g435(n948 ,n652 ,n659);
    nand g436(n1279 ,n41[4] ,n1246);
    nand g437(n1233 ,n41[2] ,n1077);
    nand g438(n1437 ,n41[1] ,n1317);
    nand g439(n838 ,n47[2] ,n617);
    dff g440(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1132), .Q(n45[3]));
    dff g441(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1999), .Q(n33[6]));
    nand g442(n2002 ,n1482 ,n1780);
    nand g443(n1053 ,n560 ,n792);
    dff g444(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1050), .Q(n51[5]));
    nand g445(n2074 ,n20[0] ,n2069);
    nand g446(n1513 ,n26[6] ,n1326);
    nand g447(n793 ,n54[3] ,n601);
    nor g448(n781 ,n386 ,n764);
    nor g449(n999 ,n936 ,n935);
    nand g450(n784 ,n21[2] ,n628);
    nor g451(n245 ,n213 ,n198);
    nand g452(n1032 ,n775 ,n785);
    nand g453(n507 ,n8[7] ,n391);
    nand g454(n1790 ,n32[6] ,n1553);
    dff g455(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1204), .Q(n57[7]));
    nand g456(n682 ,n24[3] ,n418);
    nand g457(n367 ,n2101 ,n326);
    nor g458(n603 ,n140 ,n409);
    dff g459(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2008), .Q(n36[1]));
    dff g460(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1375), .Q(n41[3]));
    nand g461(n1984 ,n1442 ,n1790);
    nand g462(n705 ,n29[1] ,n423);
    nor g463(n867 ,n222 ,n626);
    not g464(n1557 ,n1556);
    nand g465(n566 ,n8[5] ,n393);
    nand g466(n1515 ,n26[4] ,n1326);
    nand g467(n1605 ,n43[3] ,n1384);
    nand g468(n575 ,n8[4] ,n401);
    nand g469(n924 ,n748 ,n749);
    not g470(n451 ,n452);
    nor g471(n872 ,n140 ,n625);
    not g472(n610 ,n611);
    nor g473(n279 ,n257 ,n247);
    nand g474(n905 ,n56[1] ,n595);
    nand g475(n1783 ,n33[6] ,n1545);
    nand g476(n1814 ,n1283 ,n1516);
    nand g477(n876 ,n42[6] ,n599);
    nor g478(n516 ,n244 ,n424);
    nand g479(n1299 ,n41[2] ,n1251);
    nor g480(n1898 ,n1824 ,n1823);
    dff g481(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1098), .Q(n50[1]));
    xnor g482(n2119 ,n2124 ,n84);
    nand g483(n1999 ,n1485 ,n1783);
    or g484(n995 ,n928 ,n927);
    or g485(n259 ,n158 ,n227);
    dff g486(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1004), .Q(n53[0]));
    nand g487(n288 ,n22[12] ,n245);
    nand g488(n1149 ,n551 ,n978);
    nand g489(n1214 ,n58[0] ,n1079);
    dff g490(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1129), .Q(n45[4]));
    nand g491(n1135 ,n591 ,n851);
    nand g492(n1470 ,n41[3] ,n1310);
    nand g493(n440 ,n291 ,n384);
    nor g494(n1541 ,n140 ,n1316);
    nand g495(n1763 ,n37[7] ,n1543);
    nand g496(n1465 ,n41[1] ,n1314);
    nand g497(n1964 ,n1467 ,n1742);
    dff g498(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1136), .Q(n44[6]));
    nand g499(n204 ,n21[0] ,n21[1]);
    nor g500(n601 ,n140 ,n393);
    nand g501(n1430 ,n41[2] ,n1311);
    nand g502(n134 ,n279 ,n317);
    nand g503(n500 ,n8[1] ,n391);
    nand g504(n1287 ,n41[5] ,n1246);
    nand g505(n721 ,n38[7] ,n448);
    nor g506(n1018 ,n463 ,n777);
    not g507(n145 ,n39[2]);
    nand g508(n1630 ,n1172 ,n1360);
    nand g509(n526 ,n8[6] ,n401);
    nand g510(n1290 ,n41[1] ,n1246);
    nand g511(n641 ,n26[3] ,n420);
    nor g512(n767 ,n48[0] ,n604);
    nor g513(n1270 ,n41[0] ,n1245);
    nand g514(n548 ,n8[3] ,n454);
    nand g515(n815 ,n50[6] ,n621);
    nor g516(n870 ,n346 ,n627);
    nand g517(n1461 ,n41[5] ,n1314);
    nor g518(n77 ,n20[2] ,n20[0]);
    nand g519(n1631 ,n48[5] ,n1335);
    nand g520(n1752 ,n24[4] ,n1557);
    nand g521(n807 ,n52[2] ,n597);
    nand g522(n1876 ,n1583 ,n1582);
    nand g523(n2003 ,n1489 ,n1779);
    nand g524(n2047 ,n1688 ,n2030);
    nand g525(n1773 ,n36[2] ,n1547);
    nand g526(n132 ,n40[2] ,n131);
    nand g527(n1735 ,n27[5] ,n1551);
    nand g528(n931 ,n750 ,n636);
    nand g529(n760 ,n330 ,n425);
    not g530(n64 ,n63);
    dff g531(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1242), .Q(n18[1]));
    nand g532(n1621 ,n44[7] ,n1381);
    or g533(n2046 ,n1660 ,n2041);
    nand g534(n348 ,n14 ,n335);
    nand g535(n285 ,n22[11] ,n245);
    nand g536(n2040 ,n1569 ,n1917);
    dff g537(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1090), .Q(n51[2]));
    nand g538(n1635 ,n1126 ,n1352);
    dff g539(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1374), .Q(n41[2]));
    not g540(n606 ,n607);
    dff g541(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1694), .Q(n30[0]));
    nand g542(n2073 ,n19[0] ,n2081);
    dff g543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1133), .Q(n45[2]));
    nand g544(n747 ,n37[3] ,n415);
    nand g545(n656 ,n34[6] ,n416);
    dff g546(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1984), .Q(n32[6]));
    or g547(n2066 ,n1767 ,n2065);
    nand g548(n1123 ,n497 ,n844);
    nand g549(n1172 ,n60[5] ,n865);
    nor g550(n986 ,n481 ,n766);
    nand g551(n799 ,n53[2] ,n615);
    nor g552(n1336 ,n189 ,n1262);
    dff g553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1816), .Q(n26[1]));
    nor g554(n302 ,n140 ,n275);
    dff g555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2011), .Q(n36[5]));
    nand g556(n1867 ,n1573 ,n1626);
    nand g557(n1499 ,n41[7] ,n1324);
    nand g558(n851 ,n44[7] ,n623);
    not g559(n1317 ,n1318);
    nor g560(n1412 ,n41[0] ,n1313);
    nand g561(n1346 ,n1044 ,n1265);
    dff g562(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1071), .Q(n52[1]));
    nand g563(n1787 ,n33[2] ,n1545);
    nand g564(n1295 ,n41[5] ,n1251);
    nor g565(n1410 ,n41[0] ,n1304);
    nor g566(n1314 ,n190 ,n1263);
    nand g567(n565 ,n8[7] ,n409);
    nand g568(n1359 ,n60[7] ,n1252);
    nand g569(n858 ,n43[7] ,n611);
    nand g570(n2008 ,n1474 ,n1774);
    nand g571(n525 ,n8[5] ,n401);
    nor g572(n297 ,n20[4] ,n277);
    nor g573(n1316 ,n215 ,n1257);
    nand g574(n1483 ,n41[1] ,n1316);
    xnor g575(n2087 ,n39[3] ,n92);
    nand g576(n581 ,n8[2] ,n407);
    dff g577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1150), .Q(n42[7]));
    nand g578(n1871 ,n1658 ,n1523);
    nand g579(n308 ,n212 ,n269);
    nand g580(n1064 ,n582 ,n890);
    dff g581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1160), .Q(n39[3]));
    nor g582(n1271 ,n41[0] ,n1249);
    dff g583(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1057), .Q(n54[1]));
    dff g584(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1064), .Q(n53[1]));
    nand g585(n1427 ,n41[5] ,n1311);
    nand g586(n1065 ,n487 ,n801);
    dff g587(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n20[0]));
    nand g588(n1182 ,n499 ,n899);
    dff g589(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1968), .Q(n25[2]));
    nand g590(n1568 ,n49[2] ,n1334);
    dff g591(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1878), .Q(n34[4]));
    nand g592(n553 ,n8[2] ,n403);
    nor g593(n300 ,n2 ,n279);
    nor g594(n1539 ,n140 ,n1310);
    dff g595(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2013), .Q(n36[4]));
    nand g596(n1120 ,n483 ,n841);
    nand g597(n294 ,n22[9] ,n245);
    nand g598(n110 ,n22[6] ,n109);
    nor g599(n1268 ,n1020 ,n1241);
    nand g600(n2020 ,n1493 ,n1764);
    nand g601(n583 ,n8[1] ,n452);
    dff g602(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1959), .Q(n27[4]));
    nand g603(n1844 ,n1634 ,n1525);
    nand g604(n1883 ,n1665 ,n1666);
    nand g605(n1969 ,n1472 ,n1747);
    nor g606(n326 ,n303 ,n313);
    nand g607(n1205 ,n587 ,n1175);
    nand g608(n892 ,n48[7] ,n605);
    nand g609(n803 ,n52[5] ,n597);
    nor g610(n984 ,n467 ,n765);
    nand g611(n1445 ,n41[3] ,n1303);
    nand g612(n818 ,n50[2] ,n621);
    nor g613(n450 ,n248 ,n385);
    dff g614(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1598), .Q(n19[2]));
    nand g615(n511 ,n8[6] ,n397);
    nand g616(n1045 ,n2117 ,n863);
    not g617(n161 ,n20[4]);
    not g618(n1330 ,n1329);
    nand g619(n1178 ,n57[3] ,n871);
    dff g620(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1952), .Q(n28[4]));
    nand g621(n1353 ,n60[1] ,n1252);
    nor g622(n989 ,n925 ,n924);
    nand g623(n1436 ,n41[2] ,n1317);
    nor g624(n2097 ,n102 ,n100);
    nor g625(n430 ,n223 ,n366);
    nand g626(n1345 ,n340 ,n1264);
    nor g627(n466 ,n226 ,n424);
    dff g628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2007), .Q(n35[7]));
    nand g629(n1942 ,n1496 ,n1718);
    nand g630(n2113 ,n71 ,n70);
    nand g631(n286 ,n22[1] ,n245);
    xor g632(n2127 ,n20[3] ,n63);
    nand g633(n1561 ,n50[1] ,n1337);
    not g634(n137 ,n138);
    nand g635(n789 ,n54[7] ,n601);
    nor g636(n1341 ,n217 ,n1260);
    nand g637(n1422 ,n41[3] ,n1321);
    nand g638(n1170 ,n60[1] ,n865);
    nand g639(n1554 ,n1 ,n1308);
    dff g640(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1003), .Q(n42[0]));
    nand g641(n502 ,n8[2] ,n397);
    nor g642(n776 ,n51[0] ,n612);
    nand g643(n1949 ,n1454 ,n1725);
    nor g644(n2053 ,n1842 ,n2049);
    nand g645(n1026 ,n41[2] ,n867);
    nand g646(n1576 ,n45[1] ,n1386);
    nand g647(n653 ,n32[7] ,n421);
    nor g648(n364 ,n18[1] ,n330);
    nand g649(n1213 ,n930 ,n1131);
    nand g650(n1808 ,n1300 ,n1508);
    nand g651(n1739 ,n27[1] ,n1551);
    nor g652(n1579 ,n152 ,n1339);
    nand g653(n1852 ,n1643 ,n1559);
    nand g654(n1691 ,n56[7] ,n1341);
    nand g655(n491 ,n8[7] ,n411);
    nand g656(n1365 ,n383 ,n1200);
    or g657(n1007 ,n944 ,n943);
    nand g658(n704 ,n37[1] ,n415);
    nand g659(n277 ,n166 ,n242);
    dff g660(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1811), .Q(n26[6]));
    nor g661(n515 ,n8[0] ,n410);
    not g662(n1391 ,n1366);
    nand g663(n314 ,n5 ,n270);
    nand g664(n1423 ,n41[1] ,n1321);
    nand g665(n914 ,n695 ,n696);
    nand g666(n1626 ,n44[1] ,n1381);
    not g667(n346 ,n345);
    nand g668(n1645 ,n55[3] ,n1382);
    nand g669(n679 ,n32[4] ,n421);
    nor g670(n170 ,n22[10] ,n22[11]);
    nand g671(n1738 ,n27[2] ,n1551);
    nand g672(n1216 ,n232 ,n135);
    nand g673(n1127 ,n534 ,n847);
    or g674(n1260 ,n160 ,n1086);
    nand g675(n843 ,n46[4] ,n609);
    nor g676(n1710 ,n913 ,n1394);
    nand g677(n1211 ,n561 ,n1177);
    dff g678(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1094), .Q(n50[5]));
    nand g679(n1838 ,n1631 ,n1679);
    nand g680(n1278 ,n41[3] ,n1246);
    nand g681(n1040 ,n350 ,n889);
    not g682(n1389 ,n1364);
    dff g683(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1151), .Q(n42[6]));
    nand g684(n731 ,n36[3] ,n458);
    nor g685(n1917 ,n1864 ,n1863);
    nand g686(n1620 ,n48[7] ,n1335);
    nand g687(n1612 ,n57[0] ,n1380);
    nand g688(n635 ,n28[1] ,n413);
    nor g689(n423 ,n181 ,n363);
    nand g690(n729 ,n25[4] ,n459);
    not g691(n1536 ,n1537);
    nand g692(n1177 ,n57[4] ,n871);
    dff g693(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1950), .Q(n28[6]));
    not g694(n1082 ,n1083);
    nand g695(n1945 ,n1462 ,n1721);
    nand g696(n715 ,n33[0] ,n422);
    nand g697(n543 ,n8[2] ,n395);
    nand g698(n900 ,n56[5] ,n595);
    dff g699(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1872), .Q(n34[7]));
    nand g700(n509 ,n8[3] ,n391);
    dff g701(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2005), .Q(n35[5]));
    nand g702(n839 ,n47[1] ,n617);
    nand g703(n1074 ,n571 ,n809);
    nand g704(n1187 ,n530 ,n906);
    nand g705(n904 ,n56[2] ,n595);
    nand g706(n1947 ,n1465 ,n1724);
    dff g707(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1182), .Q(n56[6]));
    not g708(n1309 ,n1310);
    nand g709(n1516 ,n26[3] ,n1326);
    nand g710(n1597 ,n1048 ,n1390);
    nand g711(n967 ,n728 ,n686);
    nand g712(n965 ,n753 ,n674);
    nand g713(n321 ,n20[4] ,n311);
    nand g714(n1884 ,n1290 ,n1588);
    nand g715(n917 ,n733 ,n697);
    nand g716(n1497 ,n41[7] ,n1310);
    nand g717(n1607 ,n51[7] ,n1342);
    nor g718(n1228 ,n995 ,n990);
    nand g719(n1058 ,n539 ,n848);
    nand g720(n962 ,n342 ,n669);
    nand g721(n551 ,n8[1] ,n454);
    not g722(n87 ,n86);
    dff g723(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1107), .Q(n48[5]));
    nand g724(n1118 ,n580 ,n839);
    nand g725(n955 ,n306 ,n658);
    nand g726(n1750 ,n24[5] ,n1557);
    nand g727(n921 ,n703 ,n698);
    nor g728(n2117 ,n81 ,n79);
    nand g729(n2130 ,n74 ,n75);
    nor g730(n1425 ,n41[0] ,n1309);
    nor g731(n1940 ,n1570 ,n1865);
    nor g732(n1893 ,n1397 ,n1696);
    nand g733(n1531 ,n38[3] ,n1328);
    nand g734(n1666 ,n54[0] ,n1383);
    nand g735(n1304 ,n219 ,n1254);
    nand g736(n1070 ,n502 ,n807);
    or g737(n173 ,n140 ,n20[0]);
    nand g738(n251 ,n157 ,n194);
    nand g739(n184 ,n58[2] ,n163);
    nor g740(n180 ,n58[2] ,n58[3]);
    nand g741(n347 ,n39[0] ,n302);
    nand g742(n714 ,n25[7] ,n459);
    nand g743(n1188 ,n526 ,n888);
    nand g744(n1093 ,n488 ,n815);
    nand g745(n1101 ,n588 ,n822);
    nand g746(n103 ,n22[2] ,n102);
    nand g747(n1770 ,n36[6] ,n1547);
    nand g748(n1495 ,n41[5] ,n1316);
    nand g749(n932 ,n641 ,n682);
    nand g750(n138 ,n47[3] ,n1338);
    nand g751(n122 ,n22[13] ,n120);
    nand g752(n528 ,n8[2] ,n409);
    nand g753(n1478 ,n41[6] ,n1324);
    nand g754(n825 ,n49[1] ,n603);
    dff g755(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1958), .Q(n27[5]));
    nor g756(n307 ,n161 ,n277);
    nor g757(n1696 ,n28[0] ,n1548);
    nand g758(n1502 ,n30[6] ,n1330);
    dff g759(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1926), .Q(n32[0]));
    nor g760(n2051 ,n2042 ,n2029);
    nand g761(n229 ,n11[0] ,n1);
    xnor g762(n2118 ,n2123 ,n82);
    nand g763(n1073 ,n572 ,n808);
    nand g764(n743 ,n29[2] ,n423);
    nor g765(n1606 ,n165 ,n1388);
    nand g766(n2063 ,n1928 ,n2052);
    nor g767(n1939 ,n137 ,n1858);
    or g768(n1922 ,n1877 ,n1876);
    nand g769(n1467 ,n41[6] ,n1310);
    nand g770(n1881 ,n1664 ,n1586);
    nand g771(n571 ,n8[6] ,n450);
    nand g772(n1448 ,n41[6] ,n1307);
    dff g773(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n432), .Q(n22[6]));
    nand g774(n937 ,n642 ,n752);
    nand g775(n1369 ,n635 ,n1228);
    nand g776(n2058 ,n1939 ,n2057);
    nor g777(n1918 ,n1867 ,n1866);
    nand g778(n1099 ,n565 ,n820);
    nand g779(n343 ,n9[1] ,n311);
    nor g780(n1896 ,n1400 ,n1700);
    nand g781(n1067 ,n506 ,n803);
    dff g782(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1986), .Q(n32[4]));
    nor g783(n482 ,n8[0] ,n406);
    nand g784(n650 ,n31[7] ,n414);
    nor g785(n1335 ,n184 ,n1260);
    nand g786(n568 ,n8[4] ,n456);
    dff g787(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1089), .Q(n51[3]));
    nand g788(n1277 ,n41[7] ,n1251);
    nor g789(n418 ,n188 ,n361);
    nand g790(n1451 ,n41[3] ,n1307);
    nor g791(n315 ,n267 ,n299);
    nand g792(n372 ,n2111 ,n326);
    nand g793(n1033 ,n40[3] ,n872);
    nor g794(n457 ,n216 ,n360);
    nand g795(n1161 ,n318 ,n885);
    nor g796(n1017 ,n470 ,n771);
    nand g797(n2038 ,n1675 ,n1910);
    nor g798(n393 ,n260 ,n359);
    nand g799(n1137 ,n586 ,n853);
    nor g800(n492 ,n8[0] ,n449);
    not g801(n159 ,n14);
    dff g802(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1095), .Q(n50[4]));
    nand g803(n65 ,n20[2] ,n61);
    nand g804(n1580 ,n34[4] ,n1332);
    nand g805(n1457 ,n41[7] ,n1317);
    nand g806(n1501 ,n41[7] ,n1306);
    nand g807(n1298 ,n41[1] ,n1251);
    nand g808(n1658 ,n56[1] ,n1341);
    nand g809(n862 ,n43[3] ,n611);
    not g810(n190 ,n191);
    not g811(n604 ,n605);
    nand g812(n820 ,n49[7] ,n603);
    nand g813(n226 ,n14 ,n6);
    nor g814(n448 ,n216 ,n362);
    nand g815(n788 ,n21[1] ,n628);
    nand g816(n1816 ,n1285 ,n1519);
    nand g817(n1320 ,n191 ,n1254);
    nand g818(n1107 ,n531 ,n827);
    nand g819(n460 ,n263 ,n364);
    nor g820(n244 ,n154 ,n206);
    nand g821(n691 ,n25[5] ,n459);
    dff g822(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2012), .Q(n36[6]));
    nand g823(n1637 ,n54[4] ,n1383);
    nand g824(n845 ,n46[2] ,n609);
    nand g825(n1091 ,n574 ,n813);
    nand g826(n62 ,n20[1] ,n20[0]);
    nor g827(n1716 ,n962 ,n1407);
    nand g828(n959 ,n661 ,n727);
    nand g829(n439 ,n288 ,n373);
    nand g830(n578 ,n8[3] ,n403);
    nand g831(n1974 ,n1429 ,n1751);
    nand g832(n1943 ,n1460 ,n1719);
    nand g833(n1747 ,n25[1] ,n1539);
    dff g834(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1803), .Q(n30[7]));
    or g835(n1002 ,n917 ,n968);
    nor g836(n787 ,n365 ,n764);
    nand g837(n956 ,n665 ,n663);
    nand g838(n68 ,n19[1] ,n19[0]);
    nand g839(n664 ,n23[6] ,n419);
    dff g840(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1976), .Q(n9[0]));
    nand g841(n1116 ,n537 ,n837);
    buf g842(n12[5], 1'b0);
    nand g843(n432 ,n282 ,n357);
    dff g844(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1945), .Q(n29[4]));
    nand g845(n478 ,n8[3] ,n399);
    nand g846(n821 ,n49[6] ,n603);
    nand g847(n570 ,n8[5] ,n450);
    nor g848(n607 ,n140 ,n395);
    dff g849(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1108), .Q(n48[4]));
    nor g850(n625 ,n20[4] ,n460);
    nor g851(n2088 ,n95 ,n93);
    nand g852(n283 ,n22[2] ,n245);
    nand g853(n927 ,n633 ,n632);
    nand g854(n1489 ,n41[3] ,n1316);
    not g855(n1538 ,n1539);
    nand g856(n1587 ,n42[0] ,n1387);
    nor g857(n1717 ,n973 ,n1406);
    nand g858(n1683 ,n50[7] ,n1337);
    nor g859(n391 ,n259 ,n359);
    nor g860(n1899 ,n1826 ,n1825);
    nand g861(n792 ,n54[4] ,n601);
    nand g862(n355 ,n339 ,n332);
    dff g863(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1819), .Q(n38[3]));
    not g864(n81 ,n80);
    buf g865(n11[7], 1'b0);
    nor g866(n1324 ,n215 ,n1253);
    not g867(n332 ,n331);
    dff g868(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n199), .Q(n13[6]));
    nand g869(n1024 ,n41[4] ,n867);
    nand g870(n276 ,n176 ,n243);
    nand g871(n1723 ,n29[2] ,n1537);
    or g872(n1269 ,n1210 ,n1039);
    dff g873(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1091), .Q(n51[1]));
    dff g874(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1103), .Q(n49[3]));
    dff g875(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2026), .Q(n23[5]));
    nand g876(n655 ,n32[6] ,n421);
    nand g877(n1819 ,n1297 ,n1531);
    nand g878(n1777 ,n35[4] ,n1541);
    or g879(n303 ,n140 ,n273);
    dff g880(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1209), .Q(n57[2]));
    nand g881(n1615 ,n48[1] ,n1335);
    nand g882(n1934 ,n1431 ,n1754);
    nor g883(n980 ,n464 ,n778);
    nand g884(n1563 ,n46[3] ,n1340);
    nand g885(n925 ,n675 ,n699);
    dff g886(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1185), .Q(n56[2]));
    nor g887(n772 ,n44[0] ,n622);
    dff g888(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1348), .Q(n20[1]));
    nand g889(n1025 ,n41[3] ,n867);
    nand g890(n1601 ,n45[6] ,n1386);
    xnor g891(n2092 ,n21[2] ,n126);
    nand g892(n1766 ,n37[3] ,n1543);
    not g893(n618 ,n619);
    nand g894(n906 ,n55[7] ,n619);
    not g895(n453 ,n454);
    nand g896(n1804 ,n1272 ,n1502);
    not g897(n1262 ,n1261);
    nand g898(n2122 ,n2070 ,n2077);
    nand g899(n1618 ,n52[7] ,n1333);
    nand g900(n1966 ,n1468 ,n1743);
    nand g901(n268 ,n207 ,n236);
    nand g902(n1990 ,n1459 ,n1796);
    not g903(n1253 ,n1254);
    nand g904(n1203 ,n19[0] ,n1081);
    dff g905(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1113), .Q(n47[6]));
    not g906(n146 ,n39[3]);
    nand g907(n2027 ,n1432 ,n1758);
    dff g908(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1106), .Q(n48[6]));
    nor g909(n1925 ,n1441 ,n1707);
    dff g910(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1117), .Q(n47[2]));
    nor g911(n463 ,n8[0] ,n390);
    not g912(n141 ,n21[0]);
    nand g913(n856 ,n44[2] ,n623);
    dff g914(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n358), .Q(n22[0]));
    nand g915(n1870 ,n1576 ,n1524);
    nor g916(n1382 ,n217 ,n1259);
    nand g917(n1527 ,n38[7] ,n1328);
    nand g918(n922 ,n325 ,n757);
    nand g919(n1858 ,n1648 ,n1504);
    nand g920(n754 ,n30[2] ,n417);
    nand g921(n1375 ,n1026 ,n1234);
    nor g922(n1229 ,n983 ,n987);
    nand g923(n2035 ,n1919 ,n1918);
    nand g924(n1521 ,n34[6] ,n1332);
    nand g925(n1591 ,n43[0] ,n1384);
    nand g926(n1589 ,n42[6] ,n1387);
    dff g927(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1110), .Q(n48[2]));
    nand g928(n1456 ,n41[7] ,n1311);
    dff g929(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1159), .Q(n54[5]));
    nand g930(n291 ,n22[14] ,n245);
    not g931(n446 ,n447);
    nand g932(n710 ,n37[7] ,n415);
    nor g933(n1701 ,n23[0] ,n1534);
    nor g934(n1083 ,n228 ,n864);
    not g935(n223 ,n222);
    nand g936(n1877 ,n1585 ,n1662);
    nand g937(n828 ,n48[4] ,n605);
    nand g938(n1660 ,n1173 ,n1353);
    nor g939(n1698 ,n1270 ,n1399);
    nand g940(n1428 ,n41[4] ,n1311);
    nand g941(n1935 ,n1012 ,n1716);
    nand g942(n692 ,n33[3] ,n422);
    nand g943(n1484 ,n41[4] ,n1306);
    nand g944(n1684 ,n45[5] ,n1386);
    nand g945(n1762 ,n23[1] ,n1535);
    dff g946(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n988), .Q(n48[0]));
    nand g947(n368 ,n2097 ,n326);
    dff g948(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1995), .Q(n31[2]));
    nand g949(n1136 ,n517 ,n852);
    or g950(n992 ,n934 ,n938);
    nand g951(n690 ,n28[4] ,n413);
    nand g952(n2032 ,n1909 ,n1908);
    nand g953(n944 ,n645 ,n717);
    nand g954(n685 ,n23[4] ,n419);
    nand g955(n1803 ,n1291 ,n1610);
    nand g956(n1730 ,n28[3] ,n1549);
    or g957(n1010 ,n952 ,n951);
    nand g958(n1476 ,n41[2] ,n1306);
    nand g959(n746 ,n29[5] ,n423);
    nor g960(n1908 ,n1846 ,n1845);
    dff g961(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1936), .Q(n9[4]));
    nor g962(n182 ,n18[1] ,n18[2]);
    nand g963(n1996 ,n1453 ,n1802);
    nand g964(n357 ,n2102 ,n326);
    not g965(n143 ,n40[2]);
    nand g966(n673 ,n23[3] ,n419);
    nand g967(n577 ,n8[2] ,n393);
    nand g968(n1821 ,n1296 ,n1530);
    or g969(n1008 ,n945 ,n942);
    nand g970(n1385 ,n180 ,n1261);
    dff g971(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1804), .Q(n30[6]));
    nand g972(n1862 ,n1651 ,n1650);
    nor g973(n1395 ,n30[0] ,n1329);
    nand g974(n1206 ,n555 ,n1166);
    nand g975(n728 ,n38[0] ,n448);
    nand g976(n1088 ,n567 ,n811);
    nand g977(n1609 ,n50[6] ,n1337);
    nor g978(n623 ,n140 ,n403);
    nand g979(n1344 ,n719 ,n1226);
    not g980(n1332 ,n1331);
    nand g981(n1510 ,n45[4] ,n1386);
    nor g982(n270 ,n19[4] ,n246);
    dff g983(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1913), .Q(n36[0]));
    not g984(n311 ,n310);
    nand g985(n222 ,n18[2] ,n4);
    nand g986(n2017 ,n1477 ,n1766);
    nand g987(n1096 ,n478 ,n805);
    nand g988(n742 ,n29[3] ,n423);
    nand g989(n435 ,n285 ,n379);
    nand g990(n1948 ,n1464 ,n1723);
    dff g991(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2014), .Q(n36[7]));
    not g992(n1250 ,n1251);
    nand g993(n745 ,n35[3] ,n457);
    xnor g994(n2104 ,n22[8] ,n112);
    nand g995(n1095 ,n469 ,n817);
    nand g996(n1602 ,n42[2] ,n1387);
    nand g997(n1786 ,n33[3] ,n1545);
    nand g998(n1072 ,n224 ,n875);
    nand g999(n1740 ,n36[5] ,n1547);
    nand g1000(n2000 ,n1498 ,n1782);
    dff g1001(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1933), .Q(n9[6]));
    nand g1002(n1989 ,n1447 ,n1795);
    nand g1003(n1420 ,n41[5] ,n1321);
    nand g1004(n1988 ,n1446 ,n1891);
    nand g1005(n735 ,n36[5] ,n458);
    nand g1006(n1755 ,n36[7] ,n1547);
    or g1007(n67 ,n19[1] ,n19[0]);
    dff g1008(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1053), .Q(n54[4]));
    nand g1009(n1724 ,n29[1] ,n1537);
    nand g1010(n1827 ,n1298 ,n1393);
    nor g1011(n456 ,n249 ,n385);
    nor g1012(n421 ,n185 ,n361);
    nand g1013(n1657 ,n57[1] ,n1380);
    nor g1014(n253 ,n164 ,n182);
    dff g1015(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2010), .Q(n36[3]));
    nor g1016(n780 ,n11[3] ,n759);
    nand g1017(n1158 ,n60[7] ,n865);
    dff g1018(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n355), .Q(n39[0]));
    xnor g1019(n2090 ,n58[3] ,n96);
    dff g1020(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1906), .Q(n37[0]));
    not g1021(n1257 ,n1258);
    nor g1022(n2055 ,n2046 ,n2035);
    nand g1023(n546 ,n8[6] ,n454);
    not g1024(n123 ,n122);
    nand g1025(n1817 ,n1277 ,n1527);
    nand g1026(n1197 ,n321 ,n1043);
    buf g1027(n12[1], n11[1]);
    nand g1028(n1471 ,n41[2] ,n1310);
    dff g1029(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1147), .Q(n43[3]));
    nand g1030(n814 ,n50[7] ,n621);
    nand g1031(n181 ,n39[2] ,n146);
    nand g1032(n806 ,n52[3] ,n597);
    nand g1033(n1069 ,n503 ,n806);
    nand g1034(n1647 ,n1171 ,n1361);
    nor g1035(n783 ,n214 ,n760);
    nand g1036(n902 ,n49[3] ,n603);
    nand g1037(n1585 ,n49[0] ,n1334);
    nor g1038(n998 ,n489 ,n772);
    nand g1039(n212 ,n21[0] ,n7[3]);
    dff g1040(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2068), .Q(n60[5]));
    not g1041(n156 ,n21[2]);
    dff g1042(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n225), .Q(n10[1]));
    nor g1043(n1337 ,n189 ,n1256);
    buf g1044(n12[4], 1'b0);
    nand g1045(n1980 ,n1490 ,n1786);
    nand g1046(n1200 ,n19[3] ,n1081);
    nand g1047(n1062 ,n520 ,n798);
    or g1048(n1394 ,n912 ,n1371);
    nand g1049(n1828 ,n1517 ,n1620);
    nand g1050(n1564 ,n47[7] ,n1338);
    dff g1051(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1001), .Q(n43[0]));
    nand g1052(n1847 ,n1678 ,n1637);
    nand g1053(n585 ,n8[4] ,n403);
    nand g1054(n1486 ,n41[5] ,n1302);
    xnor g1055(n2084 ,n59[3] ,n88);
    dff g1056(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1969), .Q(n25[1]));
    nand g1057(n498 ,n8[4] ,n391);
    nor g1058(n352 ,n213 ,n333);
    nand g1059(n1351 ,n60[4] ,n1252);
    dff g1060(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1146), .Q(n43[4]));
    nand g1061(n1598 ,n1047 ,n1391);
    nand g1062(n1308 ,n219 ,n1258);
    nand g1063(n1946 ,n1463 ,n1722);
    nor g1064(n74 ,n19[2] ,n19[0]);
    dff g1065(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1983), .Q(n32[7]));
    nand g1066(n130 ,n40[1] ,n40[0]);
    nand g1067(n382 ,n2116 ,n328);
    nor g1068(n2052 ,n1883 ,n2048);
    dff g1069(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1376), .Q(n41[4]));
    nand g1070(n1358 ,n1203 ,n1239);
    nand g1071(n1048 ,n2114 ,n868);
    nand g1072(n1222 ,n58[3] ,n1079);
    nor g1073(n1398 ,n41[0] ,n1322);
    nand g1074(n748 ,n31[2] ,n414);
    nand g1075(n1477 ,n41[3] ,n1306);
    nand g1076(n1507 ,n30[2] ,n1330);
    nand g1077(n688 ,n34[4] ,n416);
    not g1078(n449 ,n450);
    nand g1079(n797 ,n53[4] ,n615);
    nand g1080(n1481 ,n41[2] ,n1324);
    nand g1081(n1987 ,n1445 ,n1793);
    nor g1082(n2094 ,n131 ,n129);
    nand g1083(n620 ,n1 ,n398);
    nor g1084(n1310 ,n186 ,n1263);
    nand g1085(n749 ,n27[2] ,n412);
    nor g1086(n1927 ,n1411 ,n1709);
    nand g1087(n2112 ,n68 ,n67);
    dff g1088(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n433), .Q(n22[4]));
    nand g1089(n586 ,n8[5] ,n403);
    nand g1090(n318 ,n39[2] ,n311);
    nand g1091(n2076 ,n19[1] ,n2081);
    nand g1092(n1036 ,n40[0] ,n863);
    dff g1093(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2066), .Q(n60[6]));
    nand g1094(n220 ,n18[1] ,n1);
    nor g1095(n1383 ,n217 ,n1256);
    not g1096(n616 ,n617);
    nor g1097(n458 ,n216 ,n361);
    nor g1098(n1381 ,n179 ,n1260);
    dff g1099(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n734), .Q(n11[0]));
    nand g1100(n837 ,n47[3] ,n617);
    nand g1101(n1991 ,n1448 ,n1797);
    dff g1102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1118), .Q(n47[1]));
    nor g1103(n242 ,n20[2] ,n173);
    nand g1104(n1846 ,n1520 ,n1636);
    nand g1105(n830 ,n48[2] ,n605);
    nor g1106(n1225 ,n1011 ,n1010);
    nand g1107(n576 ,n8[1] ,n393);
    nor g1108(n2054 ,n2045 ,n2032);
    nand g1109(n952 ,n656 ,n655);
    xnor g1110(n2083 ,n59[2] ,n86);
    nor g1111(n1397 ,n41[0] ,n1320);
    nand g1112(n587 ,n8[6] ,n452);
    nand g1113(n1929 ,n991 ,n1710);
    nand g1114(n1361 ,n60[3] ,n1252);
    not g1115(n1307 ,n1308);
    nand g1116(n1611 ,n57[4] ,n1380);
    dff g1117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2018), .Q(n37[4]));
    nand g1118(n1970 ,n1456 ,n1748);
    nor g1119(n415 ,n216 ,n363);
    nand g1120(n718 ,n36[0] ,n458);
    dff g1121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1817), .Q(n38[7]));
    dff g1122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1996), .Q(n31[1]));
    nand g1123(n200 ,n7[4] ,n156);
    nor g1124(n1021 ,n140 ,n955);
    nor g1125(n2085 ,n91 ,n89);
    not g1126(n1692 ,n1630);
    nand g1127(n1286 ,n41[6] ,n1246);
    nand g1128(n720 ,n37[0] ,n415);
    buf g1129(n13[3], n10[1]);
    nand g1130(n555 ,n8[5] ,n452);
    nand g1131(n547 ,n8[5] ,n454);
    nand g1132(n1124 ,n486 ,n845);
    nand g1133(n1443 ,n41[5] ,n1303);
    nand g1134(n2033 ,n1912 ,n1911);
    nand g1135(n953 ,n654 ,n720);
    nand g1136(n933 ,n343 ,n638);
    nand g1137(n1688 ,n46[6] ,n1340);
    nand g1138(n1078 ,n1 ,n869);
    nor g1139(n272 ,n169 ,n253);
    nand g1140(n1997 ,n1222 ,n1888);
    not g1141(n214 ,n213);
    nand g1142(n882 ,n15 ,n758);
    nand g1143(n651 ,n32[3] ,n421);
    nand g1144(n1490 ,n41[3] ,n1302);
    dff g1145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1058), .Q(n45[5]));
    nand g1146(n2075 ,n20[1] ,n2069);
    xor g1147(n2114 ,n19[3] ,n69);
    nand g1148(n1992 ,n1449 ,n1798);
    nand g1149(n1785 ,n33[4] ,n1545);
    nand g1150(n589 ,n8[6] ,n409);
    nand g1151(n1519 ,n26[1] ,n1326);
    buf g1152(n13[1], n10[1]);
    dff g1153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n468), .Q(n14));
    nand g1154(n1890 ,n2088 ,n1558);
    nand g1155(n508 ,n8[1] ,n405);
    nand g1156(n1379 ,n1033 ,n1194);
    or g1157(n168 ,n22[6] ,n22[7]);
    nor g1158(n2105 ,n114 ,n116);
    nand g1159(n811 ,n51[4] ,n613);
    dff g1160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1963), .Q(n25[7]));
    not g1161(n1321 ,n1322);
    nor g1162(n235 ,n177 ,n175);
    nand g1163(n1957 ,n1419 ,n1734);
    nor g1164(n1714 ,n960 ,n1405);
    xnor g1165(n387 ,n335 ,n14);
    dff g1166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1055), .Q(n54[2]));
    nor g1167(n195 ,n158 ,n59[3]);
    nand g1168(n337 ,n9[3] ,n311);
    dff g1169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1953), .Q(n28[3]));
    not g1170(n406 ,n407);
    or g1171(n1240 ,n20[0] ,n1075);
    nand g1172(n1811 ,n1280 ,n1513);
    nand g1173(n1659 ,n55[1] ,n1382);
    nand g1174(n1676 ,n43[4] ,n1384);
    dff g1175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1943), .Q(n29[6]));
    dff g1176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1948), .Q(n29[2]));
    nand g1177(n429 ,n377 ,n359);
    nand g1178(n552 ,n8[6] ,n447);
    nand g1179(n976 ,n688 ,n690);
    nor g1180(n100 ,n22[1] ,n22[0]);
    nand g1181(n112 ,n22[7] ,n111);
    xnor g1182(n2116 ,n2122 ,n80);
    nor g1183(n773 ,n43[0] ,n610);
    nand g1184(n1824 ,n1674 ,n1618);
    nand g1185(n1856 ,n1605 ,n1563);
    dff g1186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1980), .Q(n33[3]));
    not g1187(n1080 ,n1081);
    dff g1188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1920), .Q(n35[0]));
    nand g1189(n1567 ,n51[2] ,n1342);
    nand g1190(n1043 ,n2119 ,n863);
    nand g1191(n1288 ,n41[2] ,n1246);
    nand g1192(n1235 ,n41[4] ,n1077);
    nand g1193(n1826 ,n1607 ,n1564);
    nand g1194(n1453 ,n41[1] ,n1307);
    nor g1195(n419 ,n188 ,n360);
    or g1196(n1242 ,n462 ,n1038);
    nand g1197(n817 ,n50[4] ,n621);
    nand g1198(n898 ,n56[7] ,n595);
    nand g1199(n381 ,n2117 ,n328);
    nand g1200(n1746 ,n25[2] ,n1539);
    nand g1201(n1830 ,n1691 ,n1533);
    nand g1202(n2065 ,n1903 ,n2050);
    nand g1203(n938 ,n732 ,n746);
    nand g1204(n1151 ,n493 ,n876);
    or g1205(n274 ,n154 ,n263);
    or g1206(n1406 ,n971 ,n1354);
    nand g1207(n2126 ,n65 ,n64);
    nand g1208(n639 ,n28[6] ,n413);
    nand g1209(n1280 ,n41[6] ,n1244);
    xnor g1210(n2098 ,n22[2] ,n101);
    nand g1211(n1354 ,n683 ,n1223);
    dff g1212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1702), .Q(n38[0]));
    nand g1213(n1722 ,n29[3] ,n1537);
    nand g1214(n1726 ,n28[6] ,n1549);
    xnor g1215(n2095 ,n40[2] ,n130);
    nand g1216(n951 ,n722 ,n639);
    nor g1217(n266 ,n11[2] ,n257);
    not g1218(n334 ,n333);
    nand g1219(n706 ,n33[1] ,n422);
    xnor g1220(n2107 ,n22[11] ,n117);
    nand g1221(n1237 ,n41[6] ,n1077);
    dff g1222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n435), .Q(n22[11]));
    nand g1223(n2006 ,n1473 ,n1776);
    nand g1224(n1421 ,n41[4] ,n1321);
    dff g1225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1060), .Q(n53[5]));
    nand g1226(n1636 ,n52[4] ,n1333);
    not g1227(n1076 ,n1077);
    nor g1228(n611 ,n140 ,n454);
    nand g1229(n1102 ,n523 ,n823);
    nand g1230(n744 ,n38[4] ,n448);
    nand g1231(n923 ,n689 ,n691);
    nor g1232(n1543 ,n140 ,n1306);
    dff g1233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1161), .Q(n39[2]));
    nand g1234(n1339 ,n183 ,n1255);
    dff g1235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1706), .Q(n34[0]));
    dff g1236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1962), .Q(n27[2]));
    dff g1237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1954), .Q(n28[2]));
    nand g1238(n1794 ,n37[5] ,n1543);
    nand g1239(n740 ,n37[5] ,n415);
    dff g1240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1145), .Q(n43[5]));
    nand g1241(n1426 ,n41[6] ,n1311);
    nand g1242(n926 ,n42[7] ,n599);
    nand g1243(n1312 ,n187 ,n1254);
    dff g1244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1184), .Q(n56[3]));
    nand g1245(n1686 ,n43[6] ,n1384);
    nand g1246(n899 ,n56[6] ,n595);
    dff g1247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n436), .Q(n22[2]));
    nand g1248(n1357 ,n338 ,n1215);
    nand g1249(n634 ,n32[1] ,n421);
    nand g1250(n1044 ,n2116 ,n863);
    dff g1251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1346), .Q(n20[2]));
    nand g1252(n370 ,n2109 ,n326);
    nand g1253(n136 ,n461 ,n875);
    nand g1254(n1677 ,n53[4] ,n1336);
    nand g1255(n816 ,n50[5] ,n621);
    dff g1256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1017), .Q(n54[0]));
    nand g1257(n579 ,n8[3] ,n450);
    dff g1258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1070), .Q(n52[2]));
    nand g1259(n1196 ,n2094 ,n139);
    nand g1260(n908 ,n55[4] ,n619);
    nand g1261(n574 ,n8[1] ,n450);
    nor g1262(n613 ,n140 ,n450);
    nand g1263(n1622 ,n55[7] ,n1382);
    nand g1264(n798 ,n53[3] ,n615);
    nand g1265(n630 ,n23[1] ,n419);
    nand g1266(n1122 ,n485 ,n843);
    nor g1267(n172 ,n21[2] ,n7[5]);
    nand g1268(n262 ,n59[1] ,n195);
    dff g1269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1892), .Q(n29[0]));
    nand g1270(n437 ,n287 ,n367);
    nand g1271(n1652 ,n55[2] ,n1382);
    dff g1272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1140), .Q(n55[1]));
    nand g1273(n517 ,n8[6] ,n403);
    nand g1274(n1157 ,n494 ,n881);
    dff g1275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1934), .Q(n24[1]));
    nor g1276(n187 ,n40[2] ,n40[3]);
    nand g1277(n812 ,n51[3] ,n613);
    nor g1278(n1328 ,n140 ,n1251);
    nand g1279(n2124 ,n2078 ,n2071);
    nand g1280(n1745 ,n25[3] ,n1539);
    nand g1281(n342 ,n9[5] ,n311);
    nand g1282(n1953 ,n1416 ,n1730);
    nand g1283(n189 ,n58[3] ,n144);
    nand g1284(n379 ,n2107 ,n326);
    nor g1285(n2057 ,n2044 ,n2033);
    nand g1286(n963 ,n666 ,n664);
    nand g1287(n591 ,n8[7] ,n403);
    nand g1288(n474 ,n8[4] ,n411);
    dff g1289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1880), .Q(n34[3]));
    nand g1290(n846 ,n46[1] ,n609);
    dff g1291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1061), .Q(n53[4]));
    nand g1292(n1754 ,n24[1] ,n1557);
    nor g1293(n1570 ,n153 ,n1385);
    nor g1294(n1941 ,n1579 ,n1873);
    dff g1295(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1206), .Q(n57[5]));
    nand g1296(n804 ,n52[4] ,n597);
    dff g1297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1897), .Q(n23[0]));
    nor g1298(n1334 ,n184 ,n1262);
    nand g1299(n707 ,n38[1] ,n448);
    nand g1300(n1109 ,n524 ,n829);
    nand g1301(n557 ,n8[5] ,n447);
    nor g1302(n174 ,n22[12] ,n22[13]);
    buf g1303(n12[2], n11[2]);
    not g1304(n186 ,n187);
    nand g1305(n476 ,n8[5] ,n411);
    nand g1306(n1472 ,n41[1] ,n1310);
    nor g1307(n1241 ,n41[0] ,n1076);
    dff g1308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n233), .Q(n10[6]));
    nand g1309(n945 ,n718 ,n646);
    nand g1310(n256 ,n18[0] ,n214);
    nand g1311(n916 ,n693 ,n694);
    nor g1312(n996 ,n473 ,n770);
    nand g1313(n699 ,n35[2] ,n457);
    nand g1314(n1234 ,n41[3] ,n1077);
    nand g1315(n940 ,n710 ,n644);
    dff g1316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1183), .Q(n56[5]));
    nor g1317(n1919 ,n1869 ,n1868);
    dff g1318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1896), .Q(n24[0]));
    not g1319(n1327 ,n1328);
    nand g1320(n1454 ,n41[7] ,n1319);
    nor g1321(n2082 ,n87 ,n85);
    nand g1322(n1141 ,n553 ,n856);
    dff g1323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1059), .Q(n53[7]));
    nand g1324(n532 ,n8[4] ,n407);
    not g1325(n621 ,n620);
    dff g1326(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1930), .Q(n9[2]));
    nand g1327(n1981 ,n1220 ,n1890);
    nand g1328(n1865 ,n1655 ,n1654);
    dff g1329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1092), .Q(n50[7]));
    nor g1330(n397 ,n249 ,n359);
    nand g1331(n1986 ,n1444 ,n1792);
    nand g1332(n92 ,n39[2] ,n91);
    nand g1333(n1482 ,n41[2] ,n1316);
    nor g1334(n388 ,n315 ,n366);
    nand g1335(n1194 ,n2096 ,n139);
    nand g1336(n520 ,n8[3] ,n456);
    nor g1337(n1075 ,n302 ,n863);
    nand g1338(n531 ,n8[5] ,n407);
    buf g1339(n13[5], n10[7]);
    nor g1340(n120 ,n99 ,n119);
    or g1341(n1011 ,n957 ,n954);
    nand g1342(n736 ,n33[5] ,n422);
    dff g1343(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1139), .Q(n44[4]));
    dff g1344(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1822), .Q(n38[2]));
    nand g1345(n86 ,n59[1] ,n59[0]);
    nand g1346(n1111 ,n533 ,n831);
    nand g1347(n1180 ,n57[1] ,n871);
    nand g1348(n1139 ,n585 ,n854);
    nand g1349(n1100 ,n589 ,n821);
    nand g1350(n1417 ,n41[2] ,n1319);
    nand g1351(n1057 ,n576 ,n894);
    nand g1352(n2064 ,n1907 ,n2053);
    not g1353(n1301 ,n1302);
    nand g1354(n1719 ,n29[6] ,n1537);
    not g1355(n139 ,n864);
    dff g1356(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2019), .Q(n37[5]));
    nand g1357(n659 ,n27[7] ,n412);
    nand g1358(n1885 ,n1590 ,n1363);
    dff g1359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1219), .Q(n18[0]));
    nand g1360(n698 ,n33[2] ,n422);
    dff g1361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1935), .Q(n9[5]));
    nand g1362(n667 ,n27[6] ,n412);
    not g1363(n455 ,n456);
    dff g1364(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2002), .Q(n35[2]));
    nand g1365(n1028 ,n41[0] ,n867);
    nand g1366(n592 ,n8[2] ,n401);
    not g1367(n230 ,n229);
    nand g1368(n275 ,n2129 ,n247);
    dff g1369(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1096), .Q(n50[3]));
    nand g1370(n1665 ,n56[0] ,n1341);
    nor g1371(n510 ,n8[0] ,n451);
    nand g1372(n217 ,n58[2] ,n58[3]);
    nor g1373(n196 ,n140 ,n19[0]);
    nand g1374(n484 ,n8[5] ,n405);
    nand g1375(n1455 ,n41[7] ,n1321);
    nand g1376(n1596 ,n1049 ,n1389);
    dff g1377(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n309), .Q(n16));
    nand g1378(n2059 ,n1938 ,n2054);
    nand g1379(n689 ,n32[5] ,n421);
    nand g1380(n1956 ,n1455 ,n1733);
    nor g1381(n331 ,n39[0] ,n301);
    dff g1382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1827), .Q(n38[1]));
    nand g1383(n1998 ,n1486 ,n1784);
    nand g1384(n1751 ,n24[3] ,n1557);
    or g1385(n316 ,n22[0] ,n303);
    nand g1386(n915 ,n741 ,n671);
    nand g1387(n1578 ,n34[5] ,n1332);
    nand g1388(n1888 ,n2090 ,n1558);
    nor g1389(n407 ,n262 ,n359);
    nor g1390(n782 ,n53[0] ,n614);
    nand g1391(n71 ,n19[2] ,n67);
    dff g1392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n305), .Q(n10[3]));
    nand g1393(n631 ,n34[1] ,n416);
    nand g1394(n1239 ,n196 ,n1080);
    nand g1395(n1117 ,n538 ,n838);
    nand g1396(n936 ,n707 ,n706);
    nand g1397(n1661 ,n52[1] ,n1333);
    nor g1398(n1906 ,n1440 ,n1703);
    nand g1399(n254 ,n2081 ,n182);
    nand g1400(n1715 ,n1021 ,n1403);
    nand g1401(n700 ,n35[1] ,n457);
    nand g1402(n271 ,n234 ,n241);
    nand g1403(n1891 ,n32[2] ,n1553);
    dff g1404(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1019), .Q(n55[0]));
    nor g1405(n1003 ,n515 ,n774);
    nor g1406(n1608 ,n150 ,n1388);
    dff g1407(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1597), .Q(n19[3]));
    nand g1408(n469 ,n8[4] ,n399);
    not g1409(n158 ,n59[2]);
    or g1410(n304 ,n258 ,n265);
    nand g1411(n572 ,n8[7] ,n450);
    nand g1412(n442 ,n290 ,n369);
    nand g1413(n942 ,n715 ,n711);
    nand g1414(n94 ,n58[1] ,n58[0]);
    nand g1415(n833 ,n45[3] ,n607);
    not g1416(n396 ,n397);
    nand g1417(n480 ,n8[3] ,n411);
    nand g1418(n786 ,n43[2] ,n611);
    nand g1419(n1756 ,n23[7] ,n1535);
    nand g1420(n521 ,n8[7] ,n447);
    nand g1421(n755 ,n24[2] ,n418);
    nand g1422(n540 ,n8[4] ,n454);
    nand g1423(n443 ,n280 ,n380);
    nand g1424(n756 ,n27[3] ,n412);
    nand g1425(n1218 ,n19[4] ,n1079);
    not g1426(n602 ,n603);
    nand g1427(n1449 ,n41[5] ,n1307);
    nand g1428(n1685 ,n51[5] ,n1342);
    nand g1429(n893 ,n53[7] ,n615);
    nand g1430(n1364 ,n375 ,n1218);
    nand g1431(n684 ,n27[5] ,n412);
    nor g1432(n764 ,n154 ,n425);
    nand g1433(n2071 ,n20[4] ,n2069);
    nand g1434(n977 ,n640 ,n747);
    nand g1435(n1291 ,n41[7] ,n1248);
    nand g1436(n1373 ,n1028 ,n1232);
    dff g1437(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1067), .Q(n52[5]));
    nand g1438(n1802 ,n31[1] ,n1555);
    dff g1439(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1104), .Q(n49[1]));
    dff g1440(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1148), .Q(n43[2]));
    nand g1441(n1550 ,n1 ,n1322);
    nand g1442(n669 ,n31[5] ,n414);
    nand g1443(n119 ,n22[11] ,n118);
    nand g1444(n1646 ,n56[3] ,n1341);
    nand g1445(n881 ,n42[1] ,n599);
    nand g1446(n471 ,n8[2] ,n411);
    dff g1447(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1065), .Q(n52[7]));
    nand g1448(n293 ,n22[8] ,n245);
    nor g1449(n206 ,n159 ,n6);
    nand g1450(n1743 ,n25[5] ,n1539);
    nand g1451(n1818 ,n1294 ,n1528);
    nor g1452(n263 ,n159 ,n222);
    dff g1453(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1979), .Q(n33[2]));
    nand g1454(n1973 ,n1428 ,n1752);
    nor g1455(n1081 ,n345 ,n868);
    nand g1456(n964 ,n731 ,n673);
    nand g1457(n1275 ,n41[3] ,n1248);
    nor g1458(n1238 ,n510 ,n1030);
    nor g1459(n874 ,n304 ,n626);
    or g1460(n2045 ,n1640 ,n2038);
    nand g1461(n1689 ,n47[6] ,n1338);
    nand g1462(n1757 ,n23[5] ,n1535);
    nand g1463(n227 ,n59[1] ,n59[3]);
    nand g1464(n1599 ,n51[3] ,n1342);
    not g1465(n1551 ,n1550);
    not g1466(n179 ,n180);
    nand g1467(n563 ,n8[7] ,n452);
    nand g1468(n1833 ,n1689 ,n1609);
    nand g1469(n1772 ,n36[4] ,n1547);
    or g1470(n1016 ,n972 ,n915);
    not g1471(n1390 ,n1365);
    dff g1472(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1946), .Q(n29[3]));
    nand g1473(n896 ,n52[1] ,n597);
    nand g1474(n319 ,n39[3] ,n311);
    or g1475(n207 ,n156 ,n7[2]);
    dff g1476(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1947), .Q(n29[1]));
    nand g1477(n683 ,n30[4] ,n417);
    nor g1478(n178 ,n22[14] ,n22[15]);
    not g1479(n148 ,n19[4]);
    nand g1480(n1864 ,n1652 ,n1671);
    dff g1481(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1987), .Q(n32[3]));
    dff g1482(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1100), .Q(n49[6]));
    nor g1483(n774 ,n42[0] ,n598);
    nand g1484(n1822 ,n1299 ,n1575);
    dff g1485(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1072), .Q(n11[1]));
    nand g1486(n880 ,n42[2] ,n599);
    nand g1487(n350 ,n59[3] ,n346);
    nor g1488(n412 ,n181 ,n360);
    nand g1489(n1190 ,n575 ,n908);
    nand g1490(n1872 ,n1293 ,n1574);
    nor g1491(n409 ,n262 ,n385);
    nand g1492(n1094 ,n475 ,n816);
    nand g1493(n849 ,n45[4] ,n607);
    nand g1494(n1175 ,n57[6] ,n871);
    nand g1495(n861 ,n43[4] ,n611);
    dff g1496(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1062), .Q(n53[3]));
    not g1497(n98 ,n22[8]);
    nand g1498(n1511 ,n43[1] ,n1384);
    nand g1499(n1985 ,n1443 ,n1791);
    nand g1500(n549 ,n8[2] ,n454);
    nor g1501(n452 ,n259 ,n385);
    nor g1502(n1694 ,n1271 ,n1395);
    dff g1503(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1949), .Q(n28[7]));
    nand g1504(n1176 ,n511 ,n802);
    nand g1505(n1791 ,n32[5] ,n1553);
    dff g1506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1186), .Q(n56[1]));
    nand g1507(n1789 ,n32[7] ,n1553);
    nand g1508(n1944 ,n1461 ,n1720);
    dff g1509(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1105), .Q(n48[7]));
    or g1510(n983 ,n914 ,n965);
    nor g1511(n1038 ,n220 ,n787);
    not g1512(n1542 ,n1543);
    dff g1513(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1156), .Q(n42[2]));
    or g1514(n249 ,n59[2] ,n227);
    nor g1515(n166 ,n20[1] ,n20[3]);
    nor g1516(n991 ,n916 ,n964);
    not g1517(n162 ,n59[3]);
    dff g1518(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n434), .Q(n22[9]));
    nand g1519(n205 ,n22[4] ,n22[5]);
    nand g1520(n504 ,n8[4] ,n397);
    nand g1521(n310 ,n1 ,n275);
    nand g1522(n185 ,n39[3] ,n145);
    nand g1523(n1825 ,n1532 ,n1683);
    nand g1524(n1104 ,n529 ,n825);
    not g1525(n163 ,n58[3]);
    nand g1526(n497 ,n8[3] ,n405);
    nand g1527(n485 ,n8[4] ,n405);
    dff g1528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2028), .Q(n23[7]));
    nor g1529(n2031 ,n1905 ,n1904);
    nand g1530(n1348 ,n1045 ,n1266);
    nor g1531(n1029 ,n140 ,n781);
    nand g1532(n674 ,n23[2] ,n419);
    nand g1533(n1963 ,n1497 ,n1741);
    dff g1534(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1195), .Q(n21[1]));
    nor g1535(n1400 ,n41[0] ,n1312);
    nand g1536(n488 ,n8[6] ,n399);
    nand g1537(n909 ,n45[6] ,n607);
    nand g1538(n1841 ,n1632 ,n1619);
    nand g1539(n1452 ,n41[2] ,n1307);
    dff g1540(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1931), .Q(n9[1]));
    not g1541(n70 ,n69);
    buf g1542(n11[6], 1'b0);
    or g1543(n1006 ,n941 ,n940);
    nand g1544(n1414 ,n41[5] ,n1319);
    nand g1545(n1464 ,n41[2] ,n1314);
    nand g1546(n1678 ,n49[4] ,n1334);
    nand g1547(n850 ,n45[1] ,n607);
    nand g1548(n383 ,n2118 ,n328);
    nand g1549(n1889 ,n2089 ,n1558);
    nand g1550(n1273 ,n41[5] ,n1248);
    nand g1551(n590 ,n8[3] ,n452);
    dff g1552(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1964), .Q(n25[6]));
    nand g1553(n910 ,n55[2] ,n619);
    nor g1554(n1697 ,n27[0] ,n1550);
    nor g1555(n416 ,n185 ,n362);
    not g1556(n140 ,n1);
    nand g1557(n1843 ,n1614 ,n1633);
    nand g1558(n1444 ,n41[4] ,n1303);
    not g1559(n301 ,n302);
    nand g1560(n652 ,n26[7] ,n420);
    nand g1561(n1800 ,n31[3] ,n1555);
    nand g1562(n1728 ,n36[3] ,n1547);
    not g1563(n1305 ,n1306);
    nor g1564(n454 ,n251 ,n385);
    nor g1565(n981 ,n969 ,n963);
    nand g1566(n919 ,n754 ,n738);
    xnor g1567(n2110 ,n22[14] ,n122);
    nor g1568(n1558 ,n869 ,n1380);
    nand g1569(n697 ,n35[4] ,n457);
    not g1570(n193 ,n192);
    not g1571(n149 ,n22[1]);
    nand g1572(n885 ,n2086 ,n629);
    not g1573(n1392 ,n1367);
    nand g1574(n1169 ,n573 ,n795);
    nand g1575(n2005 ,n1495 ,n1778);
    nand g1576(n1283 ,n41[3] ,n1244);
    nand g1577(n763 ,n31[3] ,n414);
    nand g1578(n1663 ,n44[0] ,n1381);
    nand g1579(n1572 ,n49[1] ,n1334);
    nor g1580(n1384 ,n179 ,n1259);
    nand g1581(n645 ,n34[7] ,n416);
    nor g1582(n353 ,n18[2] ,n322);
    dff g1583(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1966), .Q(n25[5]));
    nor g1584(n427 ,n278 ,n352);
    nand g1585(n1955 ,n1418 ,n1732);
    nand g1586(n753 ,n32[2] ,n421);
    nor g1587(n335 ,n258 ,n312);
    nand g1588(n506 ,n8[5] ,n397);
    nand g1589(n1805 ,n1273 ,n1503);
    nand g1590(n668 ,n23[5] ,n419);
    nand g1591(n1155 ,n480 ,n879);
    nand g1592(n389 ,n274 ,n364);
    nor g1593(n778 ,n52[0] ,n596);
    nand g1594(n325 ,n9[2] ,n311);
    nor g1595(n125 ,n21[1] ,n21[0]);
    dff g1596(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1042), .Q(n59[1]));
    nand g1597(n935 ,n708 ,n705);
    dff g1598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2022), .Q(n23[1]));
    nand g1599(n732 ,n38[5] ,n448);
    nand g1600(n719 ,n35[0] ,n457);
    nor g1601(n93 ,n58[1] ,n58[0]);
    nand g1602(n1569 ,n53[2] ,n1336);
    nand g1603(n1059 ,n518 ,n893);
    nand g1604(n1628 ,n57[6] ,n1380);
    nand g1605(n1087 ,n58[0] ,n868);
    dff g1606(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1188), .Q(n55[6]));
    nand g1607(n1782 ,n33[7] ,n1545);
    not g1608(n157 ,n59[1]);
    nand g1609(n1769 ,n37[1] ,n1543);
    dff g1610(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1812), .Q(n26[5]));
    nand g1611(n632 ,n24[1] ,n418);
    nand g1612(n724 ,n38[6] ,n448);
    nand g1613(n1681 ,n53[5] ,n1336);
    nor g1614(n490 ,n8[0] ,n453);
    nand g1615(n1173 ,n60[0] ,n865);
    nor g1616(n114 ,n22[9] ,n113);
    nand g1617(n1855 ,n1562 ,n1599);
    nor g1618(n171 ,n21[2] ,n7[6]);
    nand g1619(n369 ,n2099 ,n326);
    nor g1620(n1223 ,n1016 ,n1002);
    dff g1621(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1112), .Q(n47[7]));
    nand g1622(n930 ,n21[3] ,n628);
    nor g1623(n169 ,n18[2] ,n2081);
    nand g1624(n216 ,n39[2] ,n39[3]);
    nor g1625(n210 ,n164 ,n140);
    nand g1626(n1874 ,n1286 ,n1521);
    nand g1627(n1355 ,n1034 ,n1243);
    nand g1628(n1931 ,n999 ,n1712);
    nand g1629(n1933 ,n981 ,n1714);
    nor g1630(n472 ,n8[0] ,n455);
    nand g1631(n637 ,n34[5] ,n416);
    nor g1632(n501 ,n8[0] ,n400);
    dff g1633(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n984), .Q(n50[0]));
    not g1634(n1256 ,n1255);
    xor g1635(n2128 ,n20[4] ,n66);
    nand g1636(n794 ,n2083 ,n627);
    nand g1637(n545 ,n8[6] ,n407);
    dff g1638(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1972), .Q(n24[5]));
    nand g1639(n2012 ,n1478 ,n1770);
    nor g1640(n208 ,n156 ,n7[1]);
    nand g1641(n2016 ,n1476 ,n1768);
    nand g1642(n1614 ,n55[5] ,n1382);
    nand g1643(n1853 ,n1581 ,n1560);
    nand g1644(n556 ,n8[7] ,n407);
    nand g1645(n232 ,n17 ,n1);
    nand g1646(n2021 ,n1501 ,n1763);
    nand g1647(n333 ,n155 ,n313);
    dff g1648(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1216), .Q(n17));
    nand g1649(n2060 ,n1937 ,n2051);
    nand g1650(n1581 ,n53[3] ,n1336);
    nand g1651(n2078 ,n19[4] ,n2081);
    dff g1652(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1378), .Q(n41[6]));
    nand g1653(n295 ,n22[15] ,n245);
    nand g1654(n505 ,n8[1] ,n397);
    nand g1655(n1673 ,n57[3] ,n1380);
    nor g1656(n1230 ,n1013 ,n1014);
    nand g1657(n751 ,n28[2] ,n413);
    nor g1658(n322 ,n147 ,n308);
    nand g1659(n351 ,n59[1] ,n346);
    nand g1660(n1130 ,n60[6] ,n865);
    nor g1661(n66 ,n20[3] ,n64);
    not g1662(n868 ,n869);
    not g1663(n1387 ,n1388);
    nor g1664(n401 ,n260 ,n385);
    nand g1665(n1767 ,n1639 ,n1692);
    or g1666(n987 ,n919 ,n918);
    nor g1667(n354 ,n226 ,n330);
    nand g1668(n1798 ,n31[5] ,n1555);
    nand g1669(n441 ,n295 ,n372);
    nand g1670(n1873 ,n1661 ,n1511);
    dff g1671(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1121), .Q(n46[5]));
    nand g1672(n1617 ,n54[7] ,n1383);
    nor g1673(n414 ,n185 ,n360);
    nand g1674(n376 ,n2103 ,n326);
    dff g1675(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1190), .Q(n55[4]));
    nand g1676(n255 ,n211 ,n200);
    nand g1677(n1243 ,n2095 ,n139);
    nand g1678(n444 ,n286 ,n368);
    nor g1679(n399 ,n248 ,n359);
    nand g1680(n1813 ,n1282 ,n1515);
    dff g1681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2017), .Q(n37[3]));
    nand g1682(n1880 ,n1278 ,n1584);
    nand g1683(n1761 ,n23[2] ,n1535);
    nor g1684(n2101 ,n107 ,n109);
    nor g1685(n467 ,n8[0] ,n398);
    nand g1686(n785 ,n21[0] ,n628);
    dff g1687(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1343), .Q(n58[0]));
    nand g1688(n239 ,n174 ,n178);
    dff g1689(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1074), .Q(n51[6]));
    dff g1690(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2023), .Q(n23[2]));
    nand g1691(n1514 ,n26[5] ,n1326);
    nand g1692(n894 ,n54[1] ,n601);
    nor g1693(n1030 ,n57[0] ,n870);
    nand g1694(n1774 ,n36[1] ,n1547);
    not g1695(n1546 ,n1547);
    nor g1696(n1004 ,n472 ,n782);
    nor g1697(n417 ,n181 ,n362);
    nand g1698(n519 ,n8[7] ,n393);
    not g1699(n595 ,n594);
    nand g1700(n1840 ,n1685 ,n1624);
    nand g1701(n2072 ,n20[3] ,n2069);
    nand g1702(n1823 ,n1617 ,n1603);
    dff g1703(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1971), .Q(n24[6]));
    dff g1704(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1101), .Q(n49[5]));
    dff g1705(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n230), .Q(n10[0]));
    not g1706(n104 ,n103);
    dff g1707(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n986), .Q(n49[0]));
    nor g1708(n313 ,n271 ,n264);
    nor g1709(n1911 ,n1853 ,n1852);
    nand g1710(n124 ,n22[14] ,n123);
    dff g1711(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1818), .Q(n38[6]));
    nor g1712(n175 ,n4 ,n2130);
    nand g1713(n827 ,n48[5] ,n605);
    nand g1714(n1718 ,n29[7] ,n1537);
    nand g1715(n2022 ,n1437 ,n1762);
    dff g1716(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1111), .Q(n48[1]));
    nand g1717(n1534 ,n1 ,n1318);
    nand g1718(n1281 ,n41[5] ,n1244);
    nand g1719(n750 ,n30[1] ,n417);
    nand g1720(n1343 ,n1086 ,n1214);
    nand g1721(n431 ,n292 ,n370);
    nand g1722(n1168 ,n498 ,n901);
    nand g1723(n836 ,n47[4] ,n617);
    dff g1724(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2004), .Q(n35[4]));
    nand g1725(n973 ,n336 ,n737);
    dff g1726(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1379), .Q(n40[3]));
    nand g1727(n968 ,n729 ,n677);
    dff g1728(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1127), .Q(n45[7]));
    not g1729(n1540 ,n1541);
    nand g1730(n1276 ,n41[2] ,n1248);
    nand g1731(n1842 ,n1681 ,n1682);
    nand g1732(n461 ,n237 ,n354);
    nand g1733(n1097 ,n512 ,n818);
    nand g1734(n1506 ,n30[3] ,n1330);
    nor g1735(n1914 ,n1857 ,n1856);
    nand g1736(n1119 ,n514 ,n840);
    not g1737(n135 ,n136);
    nand g1738(n2039 ,n1673 ,n1914);
    nand g1739(n1725 ,n28[7] ,n1549);
    nor g1740(n1252 ,n1078 ,n865);
    nand g1741(n722 ,n37[6] ,n415);
    dff g1742(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n443), .Q(n22[10]));
    nor g1743(n2030 ,n1902 ,n1901);
    nand g1744(n584 ,n8[2] ,n452);
    nand g1745(n1936 ,n997 ,n1717);
    nor g1746(n1706 ,n1267 ,n1409);
    not g1747(n1265 ,n1198);
    nand g1748(n890 ,n53[1] ,n615);
    nand g1749(n1649 ,n44[2] ,n1381);
    nand g1750(n1741 ,n25[7] ,n1539);
    not g1751(n1303 ,n1304);
    nand g1752(n493 ,n8[6] ,n411);
    nand g1753(n1474 ,n41[1] ,n1324);
    nand g1754(n2019 ,n1487 ,n1794);
    nand g1755(n1429 ,n41[3] ,n1311);
    not g1756(n1244 ,n1245);
    dff g1757(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2061), .Q(n60[1]));
    nand g1758(n1125 ,n508 ,n846);
    nand g1759(n1530 ,n38[4] ,n1328);
    not g1760(n614 ,n615);
    nand g1761(n128 ,n21[2] ,n127);
    nor g1762(n1921 ,n1871 ,n1870);
    dff g1763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2009), .Q(n36[2]));
    nand g1764(n101 ,n22[1] ,n22[0]);
    nand g1765(n1765 ,n37[4] ,n1543);
    not g1766(n392 ,n393);
    or g1767(n1923 ,n1881 ,n1879);
    nand g1768(n709 ,n29[0] ,n423);
    dff g1769(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1068), .Q(n52[4]));
    nor g1770(n63 ,n20[2] ,n61);
    nand g1771(n284 ,n22[4] ,n245);
    not g1772(n1248 ,n1249);
    nand g1773(n278 ,n1 ,n246);
    nand g1774(n800 ,n55[3] ,n619);
    nor g1775(n191 ,n143 ,n40[3]);
    nand g1776(n1121 ,n484 ,n842);
    nand g1777(n1496 ,n41[7] ,n1314);
    nand g1778(n1113 ,n552 ,n834);
    nand g1779(n1556 ,n1 ,n1312);
    nor g1780(n1937 ,n1606 ,n1830);
    dff g1781(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1981), .Q(n58[1]));
    nor g1782(n1537 ,n140 ,n1314);
    nand g1783(n323 ,n9[6] ,n311);
    nand g1784(n1619 ,n52[5] ,n1333);
    nand g1785(n966 ,n735 ,n668);
    dff g1786(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n296), .Q(n11[2]));
    nand g1787(n647 ,n30[7] ,n417);
    dff g1788(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1040), .Q(n59[3]));
    nand g1789(n1297 ,n41[3] ,n1251);
    nand g1790(n1145 ,n547 ,n860);
    dff g1791(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1821), .Q(n38[4]));
    nand g1792(n1199 ,n341 ,n1165);
    or g1793(n265 ,n18[0] ,n240);
    dff g1794(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n439), .Q(n22[12]));
    nand g1795(n1509 ,n47[4] ,n1338);
    or g1796(n1404 ,n946 ,n1368);
    nor g1797(n994 ,n465 ,n769);
    nand g1798(n878 ,n42[4] ,n599);
    nand g1799(n537 ,n8[3] ,n447);
    nand g1800(n2028 ,n1457 ,n1756);
    nand g1801(n703 ,n38[2] ,n448);
    nand g1802(n1533 ,n46[7] ,n1340);
    dff g1803(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1985), .Q(n32[5]));
    nor g1804(n766 ,n49[0] ,n602);
    nand g1805(n198 ,n18[0] ,n1);
    nand g1806(n1795 ,n32[1] ,n1553);
    nand g1807(n1664 ,n55[0] ,n1382);
    nand g1808(n1958 ,n1420 ,n1735);
    nor g1809(n1909 ,n1848 ,n1847);
    nand g1810(n1186 ,n500 ,n905);
    dff g1811(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1125), .Q(n46[1]));
    not g1812(n151 ,n2130);
    nand g1813(n626 ,n1 ,n426);
    nand g1814(n1347 ,n726 ,n1225);
    nand g1815(n1654 ,n48[2] ,n1335);
    nand g1816(n105 ,n22[3] ,n104);
    nand g1817(n1672 ,n52[6] ,n1333);
    nand g1818(n1577 ,n34[2] ,n1332);
    or g1819(n2044 ,n1647 ,n2039);
    dff g1820(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1810), .Q(n26[7]));
    dff g1821(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n982), .Q(n51[0]));
    nand g1822(n377 ,n59[0] ,n346);
    dff g1823(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1893), .Q(n28[0]));
    nor g1824(n982 ,n492 ,n776);
    nand g1825(n1528 ,n38[6] ,n1328);
    nand g1826(n855 ,n44[3] ,n623);
    nor g1827(n1707 ,n33[0] ,n1544);
    nand g1828(n1435 ,n41[3] ,n1317);
    nand g1829(n1098 ,n479 ,n819);
    dff g1830(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1960), .Q(n27[1]));
    nand g1831(n1995 ,n1452 ,n1801);
    or g1832(n775 ,n21[0] ,n626);
    nand g1833(n544 ,n8[1] ,n401);
    nand g1834(n1590 ,n46[0] ,n1340);
    nand g1835(n1860 ,n1566 ,n1604);
    nand g1836(n513 ,n8[5] ,n391);
    nand g1837(n1112 ,n521 ,n832);
    nand g1838(n1850 ,n1611 ,n1509);
    dff g1839(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1135), .Q(n44[7]));
    nor g1840(n241 ,n205 ,n168);
    nor g1841(n237 ,n18[2] ,n220);
    nand g1842(n918 ,n743 ,n755);
    nand g1843(n1132 ,n541 ,n833);
    dff g1844(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1088), .Q(n51[4]));
    nand g1845(n1192 ,n592 ,n910);
    nand g1846(n1463 ,n41[3] ,n1314);
    nor g1847(n75 ,n19[3] ,n73);
    nor g1848(n1342 ,n189 ,n1259);
    nand g1849(n536 ,n8[4] ,n447);
    nand g1850(n1460 ,n41[6] ,n1314);
    dff g1851(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1989), .Q(n32[1]));
    nand g1852(n644 ,n23[7] ,n419);
    nand g1853(n533 ,n8[1] ,n407);
    nor g1854(n1920 ,n1439 ,n1705);
    or g1855(n252 ,n141 ,n172);
    nand g1856(n1674 ,n53[7] ,n1336);
    nor g1857(n993 ,n496 ,n768);
    nor g1858(n201 ,n151 ,n4);
    nand g1859(n805 ,n50[3] ,n621);
    dff g1860(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1814), .Q(n26[3]));
    nand g1861(n487 ,n8[7] ,n397);
    dff g1862(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1993), .Q(n31[4]));
    nand g1863(n1523 ,n47[1] ,n1338);
    nand g1864(n686 ,n26[0] ,n420);
    nand g1865(n2026 ,n1433 ,n1757);
    or g1866(n2042 ,n1623 ,n2037);
    not g1867(n165 ,n42[7]);
    nand g1868(n1189 ,n525 ,n907);
    nand g1869(n877 ,n42[5] ,n599);
    nand g1870(n1820 ,n1295 ,n1529);
    nor g1871(n403 ,n261 ,n359);
    nand g1872(n654 ,n30[0] ,n417);
    nand g1873(n561 ,n8[4] ,n452);
    nor g1874(n447 ,n250 ,n385);
    dff g1875(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1955), .Q(n28[1]));
    nand g1876(n648 ,n24[7] ,n418);
    nand g1877(n1504 ,n50[3] ,n1337);
    nand g1878(n80 ,n2121 ,n2120);
    xor g1879(n2115 ,n19[4] ,n72);
    nand g1880(n701 ,n25[1] ,n459);
    nor g1881(n1713 ,n947 ,n1404);
    nor g1882(n988 ,n482 ,n767);
    nand g1883(n1329 ,n1 ,n1249);
    dff g1884(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1875), .Q(n34[5]));
    nor g1885(n267 ,n208 ,n252);
    dff g1886(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1181), .Q(n56[7]));
    nand g1887(n1758 ,n23[6] ,n1535);
    nand g1888(n972 ,n744 ,n679);
    nor g1889(n1251 ,n215 ,n1082);
    nand g1890(n215 ,n40[2] ,n40[3]);
    nand g1891(n1505 ,n30[4] ,n1330);
    not g1892(n624 ,n625);
    nand g1893(n115 ,n22[9] ,n113);
    nand g1894(n887 ,n20[3] ,n624);
    not g1895(n622 ,n623);
    nand g1896(n1459 ,n41[7] ,n1307);
    nand g1897(n1247 ,n219 ,n1083);
    dff g1898(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n998), .Q(n44[0]));
    nand g1899(n84 ,n2123 ,n83);
    nand g1900(n1105 ,n556 ,n892);
    nand g1901(n1863 ,n1568 ,n1594);
    nand g1902(n808 ,n51[7] ,n613);
    xnor g1903(n2086 ,n39[2] ,n90);
    nand g1904(n969 ,n702 ,n667);
    not g1905(n155 ,n18[0]);
    not g1906(n133 ,n134);
    nand g1907(n385 ,n59[0] ,n328);
    nor g1908(n1702 ,n1289 ,n1408);
    not g1909(n102 ,n101);
    nand g1910(n853 ,n44[5] ,n623);
    nand g1911(n734 ,n229 ,n461);
    nor g1912(n1333 ,n189 ,n1260);
    dff g1913(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n307), .Q(n10[2]));
    nand g1914(n1965 ,n1470 ,n1745);
    xnor g1915(n2093 ,n21[3] ,n128);
    nand g1916(n809 ,n51[6] ,n613);
    nand g1917(n1780 ,n35[2] ,n1541);
    nand g1918(n1183 ,n513 ,n900);
    nand g1919(n1466 ,n41[5] ,n1324);
    nor g1920(n1547 ,n140 ,n1324);
    nand g1921(n1051 ,n519 ,n789);
    dff g1922(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2000), .Q(n33[7]));
    dff g1923(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1977), .Q(n33[4]));
    dff g1924(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1128), .Q(n45[6]));
    nand g1925(n1524 ,n51[1] ,n1342);
    nand g1926(n1930 ,n989 ,n1711);
    nand g1927(n559 ,n8[3] ,n393);
    nand g1928(n1485 ,n41[6] ,n1302);
    nand g1929(n1060 ,n569 ,n796);
    not g1930(n597 ,n596);
    not g1931(n83 ,n82);
    dff g1932(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1895), .Q(n25[0]));
    dff g1933(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2024), .Q(n23[3]));
    nand g1934(n1952 ,n1415 ,n1729);
    dff g1935(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2015), .Q(n37[1]));
    nand g1936(n564 ,n8[2] ,n456);
    nand g1937(n338 ,n2127 ,n302);
    nand g1938(n1651 ,n57[2] ,n1380);
    nand g1939(n535 ,n8[6] ,n393);
    nand g1940(n929 ,n681 ,n678);
    nand g1941(n1641 ,n44[4] ,n1381);
    nand g1942(n1201 ,n19[2] ,n1081);
    nand g1943(n819 ,n50[1] ,n621);
    nor g1944(n481 ,n8[0] ,n408);
    not g1945(n1553 ,n1552);
    dff g1946(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1992), .Q(n31[5]));
    nand g1947(n1378 ,n1023 ,n1237);
    nand g1948(n960 ,n323 ,n662);
    nand g1949(n2121 ,n2076 ,n2075);
    nand g1950(n1126 ,n60[4] ,n865);
    dff g1951(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1114), .Q(n47[5]));
    nand g1952(n1845 ,n1613 ,n1680);
    not g1953(n1079 ,n1078);
    nand g1954(n1184 ,n509 ,n903);
    nand g1955(n375 ,n2119 ,n328);
    nand g1956(n1734 ,n27[6] ,n1551);
    nand g1957(n928 ,n704 ,n634);
    dff g1958(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n221), .Q(n13[7]));
    nand g1959(n2041 ,n1659 ,n1921);
    nand g1960(n1967 ,n1469 ,n1744);
    dff g1961(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n442), .Q(n22[3]));
    dff g1962(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1956), .Q(n27[7]));
    nand g1963(n1480 ,n41[3] ,n1324);
    dff g1964(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2021), .Q(n37[7]));
    dff g1965(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1806), .Q(n30[4]));
    nand g1966(n658 ,n31[0] ,n414);
    nand g1967(n1446 ,n41[2] ,n1303);
    dff g1968(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2020), .Q(n37[6]));
    nand g1969(n281 ,n22[0] ,n245);
    nand g1970(n1854 ,n1645 ,n1644);
    nand g1971(n1682 ,n49[5] ,n1334);
    nor g1972(n1705 ,n35[0] ,n1540);
    or g1973(n1905 ,n1841 ,n1840);
    nor g1974(n1708 ,n32[0] ,n1552);
    nand g1975(n888 ,n55[6] ,n619);
    nand g1976(n1153 ,n474 ,n878);
    nand g1977(n1648 ,n54[3] ,n1383);
    nand g1978(n1600 ,n1046 ,n1392);
    nand g1979(n479 ,n8[1] ,n399);
    nand g1980(n2014 ,n1499 ,n1755);
    nand g1981(n869 ,n201 ,n516);
    nand g1982(n374 ,n2105 ,n326);
    buf g1983(n12[7], 1'b0);
    nand g1984(n324 ,n9[7] ,n311);
    nand g1985(n1978 ,n1221 ,n1889);
    nor g1986(n2050 ,n1835 ,n2047);
    nand g1987(n813 ,n51[1] ,n613);
    nand g1988(n1737 ,n27[3] ,n1551);
    nand g1989(n1932 ,n1009 ,n1713);
    dff g1990(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1808), .Q(n30[1]));
    nor g1991(n1380 ,n217 ,n1262);
    nand g1992(n371 ,n2100 ,n326);
    not g1993(n1555 ,n1554);
    not g1994(n116 ,n115);
    nor g1995(n121 ,n22[13] ,n120);
    or g1996(n2068 ,n1771 ,n2064);
    or g1997(n1901 ,n1832 ,n1831);
    nor g1998(n420 ,n188 ,n362);
    not g1999(n1264 ,n1197);
    nor g2000(n1916 ,n1862 ,n1861);
    buf g2001(n629 ,n302);
    nor g2002(n1399 ,n26[0] ,n1325);
    nand g2003(n1983 ,n1458 ,n1789);
    nand g2004(n1159 ,n566 ,n791);
    nand g2005(n671 ,n24[4] ,n418);
    nand g2006(n1560 ,n45[3] ,n1386);
    nor g2007(n1907 ,n1844 ,n1843);
    nand g2008(n341 ,n2125 ,n302);
    nor g2009(n779 ,n55[0] ,n618);
    nor g2010(n298 ,n19[4] ,n276);
    nand g2011(n1388 ,n180 ,n1255);
    nand g2012(n1638 ,n48[4] ,n1335);
    dff g2013(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1162), .Q(n39[1]));
    nand g2014(n1972 ,n1427 ,n1750);
    nand g2015(n971 ,n680 ,n685);
    nand g2016(n2010 ,n1480 ,n1728);
    nand g2017(n860 ,n43[5] ,n611);
    dff g2018(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1205), .Q(n57[6]));
    nand g2019(n678 ,n28[5] ,n413);
    nand g2020(n1552 ,n1 ,n1304);
    dff g2021(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2062), .Q(n60[2]));
    nand g2022(n1493 ,n41[6] ,n1306);
    nand g2023(n642 ,n34[0] ,n416);
    dff g2024(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1809), .Q(n30[2]));
    nand g2025(n1143 ,n550 ,n858);
    nand g2026(n1951 ,n1414 ,n1727);
    nor g2027(n1545 ,n140 ,n1302);
    nor g2028(n777 ,n56[0] ,n594);
    nand g2029(n1834 ,n1595 ,n1627);
    or g2030(n73 ,n19[4] ,n19[1]);
    nor g2031(n1020 ,n6 ,n866);
    nand g2032(n1469 ,n41[4] ,n1310);
    or g2033(n990 ,n950 ,n961);
    nand g2034(n1163 ,n887 ,n958);
    nor g2035(n1928 ,n140 ,n1885);
    nand g2036(n340 ,n2128 ,n302);
    nand g2037(n680 ,n26[4] ,n420);
    nand g2038(n1110 ,n581 ,n830);
    nand g2039(n713 ,n29[7] ,n423);
    not g2040(n219 ,n218);
    nand g2041(n82 ,n2122 ,n81);
    nand g2042(n90 ,n39[1] ,n39[0]);
    dff g2043(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2001), .Q(n35[1]));
    nand g2044(n96 ,n58[2] ,n95);
    nand g2045(n1300 ,n41[1] ,n1248);
    nand g2046(n1653 ,n1170 ,n1362);
    nand g2047(n1041 ,n349 ,n794);
    nand g2048(n1209 ,n584 ,n1179);
    nand g2049(n539 ,n8[5] ,n395);
    nand g2050(n349 ,n59[2] ,n346);
    nand g2051(n1325 ,n1 ,n1245);
    nor g2052(n113 ,n98 ,n112);
    not g2053(n233 ,n232);
    nor g2054(n72 ,n19[3] ,n70);
    nand g2055(n2070 ,n19[2] ,n2081);
    nand g2056(n646 ,n32[0] ,n421);
    dff g2057(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1925), .Q(n33[0]));
    nand g2058(n1634 ,n57[5] ,n1380);
    dff g2059(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n445), .Q(n22[7]));
    nand g2060(n1150 ,n491 ,n926);
    nand g2061(n712 ,n35[7] ,n457);
    nand g2062(n725 ,n36[6] ,n458);
    nand g2063(n739 ,n35[5] ,n457);
    nand g2064(n844 ,n46[3] ,n609);
    nor g2065(n422 ,n185 ,n363);
    dff g2066(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1123), .Q(n46[3]));
    dff g2067(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2003), .Q(n35[3]));
    nand g2068(n1090 ,n562 ,n891);
    nor g2069(n234 ,n203 ,n202);
    nand g2070(n677 ,n27[4] ,n412);
    dff g2071(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1054), .Q(n54[3]));
    nand g2072(n943 ,n716 ,n714);
    nand g2073(n1416 ,n41[3] ,n1319);
    nand g2074(n1799 ,n31[4] ,n1555);
    nor g2075(n69 ,n19[2] ,n67);
    nand g2076(n1781 ,n35[1] ,n1541);
    dff g2077(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1974), .Q(n24[3]));
    nand g2078(n1775 ,n35[7] ,n1541);
    nand g2079(n1968 ,n1471 ,n1746);
    not g2080(n394 ,n395);
    nand g2081(n1979 ,n1491 ,n1787);
    nor g2082(n1077 ,n140 ,n867);
    nor g2083(n1255 ,n58[1] ,n1086);
    nor g2084(n1219 ,n140 ,n1031);
    dff g2085(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1176), .Q(n52[6]));
    dff g2086(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1093), .Q(n50[6]));
    buf g2087(n11[5], 1'b0);
    or g2088(n1902 ,n1834 ,n1833);
    nand g2089(n884 ,n2087 ,n629);
    dff g2090(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n298), .Q(n10[5]));
    not g2091(n164 ,n16);
    nor g2092(n1910 ,n1850 ,n1849);
    nand g2093(n2048 ,n1587 ,n2036);
    not g2094(n599 ,n598);
    nand g2095(n573 ,n8[6] ,n456);
    nand g2096(n1492 ,n41[1] ,n1302);
    nand g2097(n560 ,n8[4] ,n393);
    nor g2098(n2056 ,n2043 ,n2034);
    dff g2099(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1056), .Q(n55[3]));
    nand g2100(n1742 ,n25[6] ,n1539);
    nand g2101(n907 ,n55[5] ,n619);
    nand g2102(n1487 ,n41[5] ,n1306);
    nor g2103(n768 ,n47[0] ,n616);
    dff g2104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1032), .Q(n21[0]));
    nand g2105(n356 ,n2104 ,n326);
    nand g2106(n1744 ,n25[4] ,n1539);
    nand g2107(n1667 ,n55[6] ,n1382);
    nand g2108(n434 ,n294 ,n374);
    nand g2109(n1875 ,n1287 ,n1578);
    not g2110(n404 ,n405);
    nand g2111(n1583 ,n53[0] ,n1336);
    nand g2112(n2077 ,n20[2] ,n2069);
    nand g2113(n1285 ,n41[1] ,n1244);
    nor g2114(n1012 ,n970 ,n923);
    nand g2115(n1245 ,n187 ,n1083);
    nand g2116(n1415 ,n41[4] ,n1319);
    nand g2117(n2001 ,n1483 ,n1781);
    nor g2118(n1409 ,n34[0] ,n1331);
    nand g2119(n1146 ,n540 ,n861);
    nand g2120(n358 ,n281 ,n316);
    nor g2121(n176 ,n19[1] ,n19[2]);
    dff g2122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1144), .Q(n43[6]));
    nand g2123(n958 ,n2118 ,n625);
    nand g2124(n218 ,n40[3] ,n143);
    dff g2125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1142), .Q(n44[1]));
    dff g2126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1990), .Q(n31[7]));
    dff g2127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n994), .Q(n46[0]));
    nand g2128(n2025 ,n1434 ,n1759);
    dff g2129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1372), .Q(n41[7]));
    nand g2130(n1458 ,n41[7] ,n1303);
    nor g2131(n1900 ,n1829 ,n1828);
    xnor g2132(n2106 ,n22[10] ,n115);
    nand g2133(n2015 ,n1475 ,n1769);
    nand g2134(n1106 ,n545 ,n826);
    dff g2135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1207), .Q(n57[3]));
    nand g2136(n1886 ,n1592 ,n1591);
    nand g2137(n554 ,n8[1] ,n403);
    nand g2138(n1784 ,n33[5] ,n1545);
    nor g2139(n1411 ,n41[0] ,n1308);
    or g2140(n360 ,n39[1] ,n332);
    nand g2141(n974 ,n745 ,n763);
    nand g2142(n1801 ,n31[2] ,n1555);
    nor g2143(n192 ,n154 ,n4);
    or g2144(n359 ,n59[0] ,n327);
    nand g2145(n550 ,n8[7] ,n454);
    dff g2146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1929), .Q(n9[3]));
    nor g2147(n79 ,n2121 ,n2120);
    buf g2148(n12[6], 1'b0);
    not g2149(n1326 ,n1325);
    nand g2150(n1215 ,n311 ,n1163);
    nand g2151(n1656 ,n54[1] ,n1383);
    nand g2152(n954 ,n724 ,n723);
    dff g2153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1189), .Q(n55[5]));
    nand g2154(n1491 ,n41[2] ,n1302);
    nand g2155(n1068 ,n504 ,n804);
    nand g2156(n1575 ,n38[2] ,n1328);
    nand g2157(n1748 ,n24[7] ,n1557);
    nand g2158(n2129 ,n77 ,n78);
    nand g2159(n1204 ,n563 ,n1174);
    nand g2160(n1732 ,n28[1] ,n1549);
    nand g2161(n1848 ,n1677 ,n1510);
    or g2162(n188 ,n39[2] ,n39[3]);
    nand g2163(n542 ,n8[6] ,n395);
    dff g2164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1874), .Q(n34[6]));
    nand g2165(n1680 ,n50[4] ,n1337);
    nand g2166(n1071 ,n505 ,n896);
    dff g2167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1927), .Q(n31[0]));
    nand g2168(n1498 ,n41[7] ,n1302);
    dff g2169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2059), .Q(n60[4]));
    nand g2170(n1633 ,n44[5] ,n1381);
    nand g2171(n666 ,n31[6] ,n414);
    nand g2172(n1162 ,n320 ,n886);
    nand g2173(n711 ,n25[0] ,n459);
    nand g2174(n1749 ,n24[6] ,n1557);
    nor g2175(n1892 ,n1412 ,n1695);
    nor g2176(n1699 ,n25[0] ,n1538);
    dff g2177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n297), .Q(n10[4]));
    nand g2178(n1362 ,n60[2] ,n1252);
    nand g2179(n676 ,n28[3] ,n413);
    xnor g2180(n2096 ,n40[3] ,n132);
    nor g2181(n2091 ,n127 ,n125);
    not g2182(n600 ,n601);
    nor g2183(n489 ,n8[0] ,n402);
    dff g2184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1120), .Q(n46[6]));
    or g2185(n362 ,n142 ,n347);
    dff g2186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1951), .Q(n28[5]));
    dff g2187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1975), .Q(n24[2]));
    or g2188(n2067 ,n1924 ,n2063);
    not g2189(n1693 ,n1635);
    nand g2190(n1046 ,n2112 ,n868);
    nand g2191(n499 ,n8[6] ,n391);
    nand g2192(n1152 ,n476 ,n877);
    nand g2193(n665 ,n28[0] ,n413);
    nor g2194(n194 ,n59[2] ,n59[3]);
    nor g2195(n1402 ,n41[0] ,n1318);
    nand g2196(n1377 ,n1024 ,n1236);
    nand g2197(n694 ,n25[3] ,n459);
    nand g2198(n1142 ,n554 ,n857);
    nor g2199(n1226 ,n1008 ,n1005);
    dff g2200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1155), .Q(n42[3]));
    nand g2201(n1050 ,n570 ,n810);
    nand g2202(n852 ,n44[6] ,n623);
    nand g2203(n897 ,n45[2] ,n607);
    nand g2204(n1887 ,n1593 ,n1669);
    nand g2205(n834 ,n47[6] ,n617);
    nand g2206(n886 ,n2085 ,n629);
    not g2207(n153 ,n45[2]);
    nand g2208(n840 ,n46[7] ,n609);
    nor g2209(n758 ,n430 ,n428);
    nand g2210(n1488 ,n41[4] ,n1302);
    nand g2211(n1494 ,n41[4] ,n1316);
    buf g2212(n13[0], n10[0]);
    nand g2213(n883 ,n54[2] ,n601);
    or g2214(n361 ,n39[1] ,n347);
    nand g2215(n957 ,n660 ,n725);
    nand g2216(n2049 ,n1526 ,n2031);
    nand g2217(n1433 ,n41[5] ,n1317);
    not g2218(n398 ,n399);
    nand g2219(n857 ,n44[1] ,n623);
    nand g2220(n1475 ,n41[1] ,n1306);
    or g2221(n1259 ,n58[1] ,n1087);
    not g2222(n142 ,n39[1]);
    not g2223(n118 ,n117);
    not g2224(n2069 ,n2081);
    nand g2225(n1054 ,n559 ,n793);
    nand g2226(n1322 ,n191 ,n1258);
    nand g2227(n649 ,n28[7] ,n413);
    nand g2228(n1835 ,n1687 ,n1589);
    nand g2229(n660 ,n30[6] ,n417);
    or g2230(n1405 ,n959 ,n1347);
    nand g2231(n1779 ,n35[3] ,n1541);
    nand g2232(n1512 ,n26[7] ,n1326);
    not g2233(n312 ,n313);
    nor g2234(n1261 ,n160 ,n1087);
    nand g2235(n1994 ,n1451 ,n1800);
    dff g2236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1157), .Q(n42[1]));
    nand g2237(n693 ,n38[3] ,n448);
    or g2238(n76 ,n20[4] ,n20[1]);
    nor g2239(n365 ,n18[2] ,n329);
    nand g2240(n558 ,n8[1] ,n395);
    nand g2241(n1185 ,n495 ,n904);
    nor g2242(n619 ,n140 ,n401);
    nor g2243(n236 ,n21[0] ,n171);
    nand g2244(n670 ,n30[5] ,n417);
    nand g2245(n514 ,n8[7] ,n405);
    not g2246(n329 ,n330);
    nand g2247(n687 ,n31[4] ,n414);
    dff g2248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1213), .Q(n21[3]));
    nand g2249(n1573 ,n53[1] ,n1336);
    nor g2250(n1894 ,n1398 ,n1697);
    not g2251(n863 ,n864);
    nand g2252(n1594 ,n50[2] ,n1337);
    nand g2253(n1644 ,n52[3] ,n1333);
    nand g2254(n2029 ,n1899 ,n1898);
    nor g2255(n1408 ,n38[0] ,n1327);
    nor g2256(n411 ,n251 ,n359);
    dff g2257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1029), .Q(n18[2]));
    or g2258(n1086 ,n58[0] ,n869);
    or g2259(n61 ,n20[1] ,n20[0]);
    nand g2260(n941 ,n713 ,n712);
    nand g2261(n1861 ,n1567 ,n1602);
    dff g2262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2067), .Q(n60[0]));
    or g2263(n1976 ,n985 ,n1715);
    nand g2264(n854 ,n44[4] ,n623);
    nand g2265(n2061 ,n1941 ,n2055);
    nand g2266(n903 ,n56[3] ,n595);
    xnor g2267(n2099 ,n22[3] ,n103);
    nand g2268(n879 ,n42[3] ,n599);
    nand g2269(n593 ,n8[4] ,n395);
    not g2270(n1323 ,n1324);
    nor g2271(n78 ,n20[3] ,n76);
    nand g2272(n1047 ,n2113 ,n868);
    nand g2273(n829 ,n48[3] ,n605);
    nand g2274(n1727 ,n28[5] ,n1549);
    nand g2275(n475 ,n8[5] ,n399);
    dff g2276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1063), .Q(n53[2]));
    nand g2277(n1249 ,n191 ,n1083);
    dff g2278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1141), .Q(n44[2]));
    dff g2279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1957), .Q(n27[6]));
    nand g2280(n384 ,n2110 ,n326);
    nand g2281(n1231 ,n41[7] ,n1077);
    nand g2282(n1629 ,n54[5] ,n1383);
    dff g2283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n438), .Q(n22[8]));
    nand g2284(n1263 ,n40[1] ,n1084);
    dff g2285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1932), .Q(n9[7]));
    nor g2286(n89 ,n39[1] ,n39[0]);
    nand g2287(n345 ,n1 ,n314);
    not g2288(n408 ,n409);
    nand g2289(n1419 ,n41[6] ,n1321);
    nand g2290(n380 ,n2106 ,n326);
    nand g2291(n2079 ,n19[3] ,n2081);
    nand g2292(n1592 ,n47[0] ,n1338);
    dff g2293(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1153), .Q(n42[4]));
    nand g2294(n1851 ,n1642 ,n1641);
    nor g2295(n1084 ,n40[0] ,n864);
    not g2296(n1311 ,n1312);
    nand g2297(n970 ,n740 ,n684);
    nor g2298(n129 ,n40[1] ,n40[0]);
    nand g2299(n126 ,n21[1] ,n21[0]);
    nor g2300(n628 ,n278 ,n426);
    nand g2301(n889 ,n2084 ,n627);
    not g2302(n1544 ,n1545);
    nand g2303(n2023 ,n1436 ,n1761);
    nand g2304(n1236 ,n41[5] ,n1077);
    nor g2305(n425 ,n300 ,n133);
    nand g2306(n1721 ,n29[4] ,n1537);
    nand g2307(n228 ,n40[0] ,n40[1]);
    nand g2308(n1174 ,n57[7] ,n871);
    nand g2309(n975 ,n730 ,n687);
    nand g2310(n1154 ,n2091 ,n874);
    nor g2311(n243 ,n19[3] ,n197);
    or g2312(n1904 ,n1839 ,n1838);
    nand g2313(n638 ,n31[1] ,n414);
    nand g2314(n1582 ,n50[0] ,n1337);
    dff g2315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1187), .Q(n55[7]));
    nand g2316(n320 ,n39[1] ,n311);
    nand g2317(n841 ,n46[6] ,n609);
    nand g2318(n695 ,n36[2] ,n458);
    nand g2319(n950 ,n631 ,n701);
    dff g2320(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1998), .Q(n33[5]));
    nand g2321(n1171 ,n60[2] ,n865);
    nor g2322(n386 ,n258 ,n365);
    nand g2323(n1179 ,n57[2] ,n871);
    nand g2324(n1027 ,n41[1] ,n867);
    nand g2325(n562 ,n8[2] ,n450);
    nand g2326(n823 ,n49[4] ,n603);
    dff g2327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2060), .Q(n60[7]));
    nand g2328(n273 ,n256 ,n254);
    dff g2329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1805), .Q(n30[5]));
    nor g2330(n1700 ,n24[0] ,n1556);
    dff g2331(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1982), .Q(n33[1]));
    nand g2332(n1055 ,n577 ,n883);
    nand g2333(n730 ,n33[4] ,n422);
    nand g2334(n1529 ,n38[5] ,n1328);
    nand g2335(n1034 ,n40[2] ,n872);
    dff g2336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1069), .Q(n52[3]));
    nand g2337(n524 ,n8[3] ,n407);
    nand g2338(n1520 ,n51[4] ,n1342);
    nand g2339(n1796 ,n31[7] ,n1555);
    nand g2340(n708 ,n36[1] ,n458);
    nand g2341(n810 ,n51[5] ,n613);
    nand g2342(n1586 ,n51[0] ,n1342);
    nand g2343(n1103 ,n527 ,n902);
    nand g2344(n1147 ,n548 ,n862);
    not g2345(n866 ,n867);
    nand g2346(n978 ,n43[1] ,n611);
    nand g2347(n596 ,n1 ,n396);
    nand g2348(n1393 ,n38[1] ,n1328);
    xnor g2349(n2108 ,n22[12] ,n119);
    not g2350(n199 ,n198);
    nand g2351(n373 ,n2108 ,n326);
    nand g2352(n961 ,n700 ,n630);
    nand g2353(n1292 ,n41[7] ,n1244);
    nand g2354(n494 ,n8[1] ,n411);
    nand g2355(n1624 ,n46[5] ,n1340);
    nand g2356(n636 ,n27[1] ,n412);
    nand g2357(n1961 ,n1422 ,n1737);
    not g2358(n1246 ,n1247);
    dff g2359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1942), .Q(n29[7]));
    not g2360(n402 ,n403);
    nand g2361(n1720 ,n29[5] ,n1537);
    nor g2362(n470 ,n8[0] ,n392);
    dff g2363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n440), .Q(n22[14]));
    nand g2364(n947 ,n324 ,n650);
    nand g2365(n1202 ,n19[1] ,n1081);
    nand g2366(n702 ,n25[6] ,n459);
    nand g2367(n1993 ,n1450 ,n1799);
    nand g2368(n1532 ,n49[7] ,n1334);
    nand g2369(n569 ,n8[5] ,n456);
    nand g2370(n1522 ,n42[5] ,n1387);
    nor g2371(n1695 ,n29[0] ,n1536);
    nor g2372(n1897 ,n1402 ,n1701);
    dff g2373(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2006), .Q(n35[6]));
    dff g2374(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n444), .Q(n22[1]));
    dff g2375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1099), .Q(n49[7]));
    nand g2376(n2123 ,n2079 ,n2072);
    not g2377(n612 ,n613);
    dff g2378(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1137), .Q(n44[5]));
    dff g2379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n429), .Q(n59[0]));
    dff g2380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1119), .Q(n46[7]));
    nor g2381(n1009 ,n949 ,n948);
    nor g2382(n413 ,n181 ,n361);
    not g2383(n152 ,n46[1]);
    nand g2384(n1971 ,n1426 ,n1749);
    nand g2385(n801 ,n52[7] ,n597);
    nand g2386(n1022 ,n41[6] ,n867);
    nand g2387(n723 ,n35[6] ,n457);
    nand g2388(n1418 ,n41[1] ,n1319);
    or g2389(n2043 ,n1653 ,n2040);
    nand g2390(n1208 ,n583 ,n1180);
    dff g2391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1973), .Q(n24[4]));
    dff g2392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1122), .Q(n46[4]));
    nand g2393(n1191 ,n528 ,n824);
    nand g2394(n1623 ,n1130 ,n1359);
    nand g2395(n1812 ,n1281 ,n1514);
    nand g2396(n1776 ,n35[6] ,n1541);
    nor g2397(n617 ,n140 ,n447);
    nand g2398(n859 ,n43[6] ,n611);
    nand g2399(n1442 ,n41[6] ,n1303);
    nand g2400(n1690 ,n53[6] ,n1336);
    nand g2401(n1138 ,n2092 ,n874);
    nor g2402(n1440 ,n41[0] ,n1305);
    nand g2403(n946 ,n649 ,n648);
    nor g2404(n1031 ,n761 ,n783);
    nor g2405(n1403 ,n953 ,n1344);
    not g2406(n247 ,n246);
    nor g2407(n1254 ,n40[1] ,n1036);
    nand g2408(n1668 ,n48[6] ,n1335);
    nor g2409(n85 ,n59[1] ,n59[0]);
    nand g2410(n1866 ,n1572 ,n1571);
    nand g2411(n2081 ,n18[0] ,n2080);
    nand g2412(n503 ,n8[3] ,n397);
    dff g2413(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1994), .Q(n31[3]));
    nand g2414(n1879 ,n1612 ,n1663);
    nand g2415(n1508 ,n30[1] ,n1330);
    nand g2416(n211 ,n21[2] ,n7[0]);
    dff g2417(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n431), .Q(n22[13]));
    nand g2418(n1366 ,n382 ,n1201);
    nand g2419(n1131 ,n2093 ,n874);
    dff g2420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1015), .Q(n11[3]));
    nor g2421(n770 ,n45[0] ,n606);
    nand g2422(n330 ,n18[0] ,n313);
    nand g2423(n1432 ,n41[6] ,n1317);
    nor g2424(n1306 ,n215 ,n1263);
    nand g2425(n1810 ,n1292 ,n1512);
    nand g2426(n842 ,n46[5] ,n609);
    nand g2427(n213 ,n18[1] ,n18[2]);
    nand g2428(n847 ,n45[7] ,n607);
    nand g2429(n1424 ,n41[2] ,n1321);
    not g2430(n144 ,n58[2]);
    nand g2431(n1363 ,n60[0] ,n1252);
    nand g2432(n1518 ,n26[2] ,n1326);
    nand g2433(n523 ,n8[4] ,n409);
    buf g2434(n12[0], n11[0]);
endmodule
