module top (n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [2:0] n6;
    wire [63:0] n7;
    wire [7:0] n8;
    wire [19:0] n9;
    wire n10, n11, n12, n13, n14, n15, n16, n17;
    wire n18, n19, n20, n21, n22, n23, n24, n25;
    wire n26, n27, n28, n29, n30, n31, n32, n33;
    wire n34, n35, n36, n37, n38, n39, n40, n41;
    wire n42, n43, n44, n45, n46, n47, n48, n49;
    wire n50, n51, n52, n53, n54, n55, n56, n57;
    wire n58, n59, n60, n61, n62, n63, n64, n65;
    wire n66, n67, n68, n69, n70, n71, n72, n73;
    wire n74, n75, n76, n77, n78, n79, n80, n81;
    wire n82, n83, n84, n85, n86, n87, n88, n89;
    wire n90, n91, n92, n93, n94, n95, n96, n97;
    wire n98, n99, n100, n101, n102, n103, n104, n105;
    wire n106, n107, n108, n109, n110, n111, n112, n113;
    wire n114, n115, n116, n117, n118, n119, n120, n121;
    wire n122, n123, n124, n125, n126, n127, n128, n129;
    wire n130, n131, n132, n133, n134, n135, n136, n137;
    wire n138, n139, n140, n141, n142, n143, n144, n145;
    wire n146, n147, n148, n149, n150, n151, n152, n153;
    wire n154, n155, n156, n157, n158, n159, n160, n161;
    wire n162, n163, n164, n165, n166, n167, n168, n169;
    wire n170, n171, n172, n173, n174, n175, n176, n177;
    wire n178, n179, n180, n181, n182, n183, n184, n185;
    wire n186, n187, n188, n189, n190, n191, n192, n193;
    wire n194, n195, n196, n197, n198, n199, n200, n201;
    wire n202, n203, n204, n205, n206, n207, n208, n209;
    wire n210, n211, n212, n213, n214, n215, n216, n217;
    wire n218, n219, n220, n221, n222, n223, n224, n225;
    wire n226, n227, n228, n229, n230, n231, n232, n233;
    wire n234, n235, n236, n237, n238, n239, n240, n241;
    wire n242, n243, n244, n245, n246, n247, n248, n249;
    wire n250, n251, n252, n253, n254, n255, n256, n257;
    wire n258, n259, n260, n261, n262, n263, n264, n265;
    wire n266, n267, n268, n269, n270, n271, n272, n273;
    wire n274, n275, n276, n277, n278, n279, n280, n281;
    wire n282, n283, n284, n285, n286, n287, n288, n289;
    wire n290, n291, n292, n293, n294, n295, n296, n297;
    wire n298, n299, n300, n301, n302, n303, n304, n305;
    wire n306, n307, n308, n309, n310, n311, n312, n313;
    wire n314, n315, n316, n317, n318, n319, n320, n321;
    wire n322, n323, n324, n325, n326, n327, n328, n329;
    wire n330, n331, n332, n333, n334, n335, n336, n337;
    wire n338, n339, n340, n341, n342, n343, n344, n345;
    wire n346, n347, n348, n349, n350, n351, n352, n353;
    wire n354, n355, n356, n357, n358, n359, n360, n361;
    wire n362, n363, n364, n365, n366, n367, n368, n369;
    wire n370, n371, n372, n373, n374, n375, n376, n377;
    wire n378, n379, n380, n381, n382, n383, n384, n385;
    wire n386, n387, n388, n389, n390, n391, n392, n393;
    wire n394, n395, n396, n397, n398, n399, n400, n401;
    wire n402, n403, n404, n405, n406, n407, n408, n409;
    wire n410, n411, n412, n413, n414, n415, n416, n417;
    wire n418, n419, n420, n421, n422, n423, n424, n425;
    wire n426, n427, n428, n429, n430, n431, n432, n433;
    wire n434, n435, n436, n437, n438, n439, n440, n441;
    wire n442, n443, n444, n445, n446, n447, n448, n449;
    wire n450, n451, n452, n453, n454, n455, n456, n457;
    wire n458, n459, n460, n461, n462, n463, n464, n465;
    wire n466, n467, n468, n469, n470, n471, n472, n473;
    wire n474, n475, n476, n477, n478, n479, n480, n481;
    wire n482, n483, n484, n485, n486, n487, n488, n489;
    wire n490, n491, n492, n493, n494, n495, n496, n497;
    wire n498, n499, n500, n501, n502, n503, n504, n505;
    wire n506, n507, n508, n509, n510, n511, n512, n513;
    wire n514, n515, n516, n517, n518, n519, n520, n521;
    wire n522, n523, n524, n525, n526, n527, n528, n529;
    wire n530, n531, n532, n533, n534, n535, n536, n537;
    wire n538, n539, n540, n541, n542, n543, n544, n545;
    wire n546, n547, n548, n549, n550, n551, n552, n553;
    wire n554, n555, n556, n557, n558, n559, n560, n561;
    wire n562, n563, n564, n565, n566, n567, n568, n569;
    wire n570, n571, n572, n573, n574, n575, n576, n577;
    wire n578, n579, n580, n581, n582, n583, n584, n585;
    wire n586, n587, n588, n589, n590, n591, n592, n593;
    wire n594, n595, n596, n597, n598, n599, n600, n601;
    wire n602, n603, n604, n605, n606, n607, n608, n609;
    wire n610, n611, n612, n613, n614, n615, n616, n617;
    wire n618, n619, n620, n621, n622, n623, n624, n625;
    wire n626, n627, n628, n629, n630, n631, n632, n633;
    wire n634, n635, n636, n637, n638, n639, n640, n641;
    wire n642, n643, n644, n645, n646, n647, n648, n649;
    wire n650, n651, n652, n653, n654, n655, n656, n657;
    wire n658, n659, n660, n661, n662, n663, n664, n665;
    wire n666, n667, n668, n669, n670, n671, n672, n673;
    wire n674, n675, n676, n677, n678, n679, n680, n681;
    wire n682, n683, n684, n685, n686, n687, n688, n689;
    wire n690, n691, n692, n693, n694, n695, n696, n697;
    wire n698, n699, n700, n701, n702, n703, n704, n705;
    wire n706, n707, n708, n709, n710, n711, n712, n713;
    wire n714, n715, n716, n717, n718, n719, n720, n721;
    wire n722, n723, n724, n725, n726, n727, n728, n729;
    wire n730, n731, n732, n733, n734, n735, n736, n737;
    wire n738, n739, n740, n741, n742, n743, n744, n745;
    wire n746, n747, n748, n749, n750, n751, n752, n753;
    wire n754, n755, n756, n757, n758, n759, n760, n761;
    wire n762, n763, n764, n765, n766, n767, n768, n769;
    wire n770, n771, n772, n773, n774, n775, n776, n777;
    wire n778, n779, n780, n781, n782, n783, n784, n785;
    wire n786, n787, n788, n789, n790, n791, n792, n793;
    wire n794, n795, n796, n797, n798, n799, n800, n801;
    wire n802, n803, n804, n805, n806, n807, n808, n809;
    wire n810, n811, n812, n813, n814, n815, n816, n817;
    wire n818, n819, n820, n821, n822, n823, n824, n825;
    wire n826, n827, n828, n829, n830, n831, n832, n833;
    wire n834, n835, n836, n837, n838, n839, n840, n841;
    wire n842, n843, n844, n845, n846, n847, n848, n849;
    wire n850, n851, n852, n853, n854, n855, n856, n857;
    wire n858, n859, n860, n861, n862, n863, n864, n865;
    wire n866, n867, n868, n869, n870, n871, n872, n873;
    wire n874, n875, n876, n877, n878, n879, n880, n881;
    wire n882, n883, n884, n885, n886, n887, n888, n889;
    wire n890, n891, n892, n893, n894, n895, n896, n897;
    wire n898, n899, n900, n901, n902, n903, n904, n905;
    wire n906, n907, n908, n909, n910, n911, n912, n913;
    wire n914, n915, n916, n917, n918, n919, n920, n921;
    wire n922, n923, n924, n925, n926, n927, n928, n929;
    wire n930, n931, n932, n933, n934, n935, n936, n937;
    wire n938, n939, n940, n941, n942, n943, n944, n945;
    wire n946, n947, n948, n949, n950, n951, n952, n953;
    wire n954, n955, n956, n957, n958, n959, n960, n961;
    wire n962, n963, n964, n965, n966, n967, n968, n969;
    wire n970, n971, n972, n973, n974, n975, n976, n977;
    wire n978, n979, n980, n981, n982, n983, n984, n985;
    wire n986, n987, n988, n989, n990, n991, n992, n993;
    wire n994, n995, n996, n997, n998, n999, n1000, n1001;
    wire n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009;
    wire n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017;
    wire n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
    wire n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
    wire n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041;
    wire n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049;
    wire n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057;
    wire n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065;
    wire n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073;
    wire n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081;
    wire n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089;
    wire n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097;
    wire n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105;
    wire n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113;
    wire n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121;
    wire n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129;
    wire n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137;
    wire n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145;
    wire n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153;
    wire n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161;
    wire n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169;
    wire n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177;
    wire n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185;
    wire n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193;
    wire n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201;
    wire n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209;
    wire n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217;
    wire n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225;
    wire n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233;
    wire n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241;
    wire n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249;
    wire n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257;
    wire n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265;
    wire n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273;
    wire n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281;
    wire n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289;
    wire n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297;
    wire n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305;
    wire n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313;
    wire n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321;
    wire n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329;
    wire n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;
    wire n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345;
    wire n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353;
    wire n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;
    wire n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369;
    wire n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377;
    wire n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385;
    wire n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393;
    wire n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401;
    wire n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409;
    wire n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417;
    wire n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425;
    wire n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433;
    wire n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441;
    wire n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449;
    wire n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457;
    wire n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465;
    wire n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473;
    wire n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481;
    wire n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489;
    wire n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497;
    wire n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505;
    wire n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513;
    wire n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521;
    wire n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529;
    wire n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537;
    wire n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545;
    wire n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553;
    wire n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561;
    wire n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569;
    wire n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577;
    wire n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585;
    wire n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593;
    wire n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601;
    wire n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609;
    wire n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617;
    wire n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625;
    wire n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633;
    wire n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641;
    wire n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649;
    wire n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657;
    wire n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665;
    wire n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673;
    wire n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681;
    wire n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689;
    wire n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697;
    wire n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705;
    wire n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713;
    wire n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721;
    wire n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729;
    wire n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737;
    wire n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745;
    wire n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753;
    wire n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761;
    wire n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769;
    wire n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777;
    wire n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785;
    wire n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793;
    wire n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801;
    wire n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809;
    wire n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817;
    wire n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825;
    wire n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833;
    wire n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;
    wire n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849;
    wire n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857;
    wire n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865;
    wire n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873;
    wire n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881;
    wire n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889;
    wire n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897;
    wire n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905;
    wire n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913;
    wire n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921;
    wire n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929;
    wire n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937;
    wire n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945;
    wire n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953;
    wire n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961;
    wire n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969;
    wire n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977;
    wire n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985;
    wire n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993;
    wire n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001;
    wire n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009;
    wire n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017;
    wire n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025;
    wire n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033;
    wire n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041;
    wire n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049;
    wire n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057;
    wire n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065;
    wire n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073;
    wire n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081;
    wire n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089;
    wire n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097;
    wire n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105;
    wire n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113;
    wire n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121;
    wire n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129;
    wire n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137;
    wire n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145;
    wire n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153;
    wire n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161;
    wire n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169;
    wire n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177;
    wire n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185;
    wire n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193;
    wire n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201;
    wire n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209;
    wire n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217;
    wire n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225;
    wire n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233;
    wire n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241;
    wire n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249;
    wire n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257;
    wire n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265;
    wire n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273;
    wire n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281;
    wire n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289;
    wire n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297;
    wire n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305;
    wire n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313;
    wire n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321;
    wire n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329;
    wire n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337;
    wire n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345;
    wire n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353;
    wire n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361;
    wire n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369;
    wire n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377;
    wire n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385;
    wire n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393;
    wire n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401;
    wire n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409;
    wire n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417;
    wire n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425;
    wire n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433;
    wire n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441;
    wire n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449;
    wire n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457;
    wire n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465;
    wire n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473;
    wire n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481;
    wire n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489;
    wire n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497;
    wire n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505;
    wire n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513;
    wire n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521;
    wire n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529;
    wire n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537;
    wire n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545;
    wire n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553;
    wire n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561;
    wire n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569;
    wire n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577;
    wire n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585;
    wire n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593;
    wire n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601;
    wire n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609;
    wire n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617;
    wire n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625;
    wire n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633;
    wire n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641;
    wire n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649;
    wire n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657;
    wire n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665;
    wire n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673;
    wire n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681;
    wire n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689;
    wire n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697;
    wire n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705;
    wire n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713;
    wire n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721;
    wire n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729;
    wire n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737;
    wire n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745;
    wire n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753;
    wire n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761;
    wire n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769;
    wire n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777;
    wire n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785;
    wire n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793;
    wire n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801;
    wire n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809;
    wire n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817;
    wire n2818, n2819;
    nand g0(n1159 ,n2324 ,n650);
    xnor g1(n2337 ,n74 ,n192);
    or g2(n912 ,n452 ,n586);
    nand g3(n1008 ,n4[17] ,n565);
    nand g4(n2741 ,n4[53] ,n2736);
    nand g5(n1085 ,n2350 ,n651);
    nand g6(n2189 ,n2[4] ,n6[1]);
    nand g7(n2220 ,n2042 ,n3[9]);
    xor g8(n2308 ,n2436 ,n2372);
    nor g9(n1708 ,n1027 ,n1518);
    nand g10(n1990 ,n1385 ,n1833);
    nor g11(n1837 ,n1034 ,n1770);
    nand g12(n1061 ,n364 ,n476);
    nand g13(n1981 ,n1376 ,n1824);
    nand g14(n1341 ,n741 ,n1271);
    nand g15(n2050 ,n2[16] ,n6[1]);
    xnor g16(n2350 ,n130 ,n218);
    nand g17(n2655 ,n2654 ,n2653);
    nand g18(n1912 ,n1134 ,n1663);
    nand g19(n2651 ,n2647 ,n2646);
    nand g20(n2398 ,n2121 ,n2120);
    or g21(n524 ,n3[36] ,n465);
    nor g22(n1884 ,n1025 ,n1769);
    not g23(n2662 ,n2661);
    nand g24(n2408 ,n2216 ,n2211);
    xnor g25(n2360 ,n122 ,n238);
    xnor g26(n96 ,n2469 ,n2405);
    nand g27(n1580 ,n2[106] ,n1259);
    nand g28(n2421 ,n2193 ,n2185);
    nor g29(n2250 ,n2576 ,n2578);
    nor g30(n2697 ,n2507 ,n2692);
    nor g31(n177 ,n131 ,n176);
    or g32(n14 ,n2437 ,n2373);
    nor g33(n31 ,n2490 ,n2426);
    or g34(n2653 ,n4[29] ,n2649);
    nor g35(n648 ,n7[7] ,n462);
    nand g36(n853 ,n427 ,n568);
    nand g37(n2146 ,n2[82] ,n6[1]);
    nand g38(n1939 ,n1164 ,n1691);
    not g39(n271 ,n270);
    nand g40(n1781 ,n1327 ,n1395);
    nand g41(n399 ,n2324 ,n274);
    nand g42(n989 ,n347 ,n513);
    nand g43(n956 ,n354 ,n491);
    nand g44(n2579 ,n4[7] ,n2578);
    nor g45(n216 ,n19 ,n215);
    nand g46(n2462 ,n2141 ,n2073);
    or g47(n2793 ,n9[5] ,n1);
    nand g48(n374 ,n2337 ,n273);
    nand g49(n2112 ,n2[107] ,n6[1]);
    nor g50(n2615 ,n4[18] ,n2613);
    nand g51(n1444 ,n706 ,n1234);
    nor g52(n810 ,n5[12] ,n621);
    xnor g53(n85 ,n2460 ,n2396);
    nand g54(n447 ,n2246 ,n312);
    nand g55(n1527 ,n844 ,n1332);
    nor g56(n2756 ,n2755 ,n2754);
    nor g57(n1601 ,n841 ,n1411);
    nand g58(n625 ,n7[31] ,n461);
    nand g59(n2676 ,n2673 ,n2672);
    nor g60(n2727 ,n2509 ,n2724);
    nand g61(n2179 ,n2043 ,n3[56]);
    nand g62(n623 ,n7[23] ,n461);
    nor g63(n2531 ,n2516 ,n4[11]);
    or g64(n1381 ,n2[108] ,n1263);
    nand g65(n1777 ,n1586 ,n1047);
    xor g66(n2807 ,n2[2] ,n9[2]);
    nand g67(n2188 ,n2[34] ,n6[1]);
    or g68(n576 ,n4[40] ,n464);
    nand g69(n866 ,n4[19] ,n565);
    nand g70(n1117 ,n2[42] ,n560);
    nand g71(n1056 ,n4[30] ,n647);
    nand g72(n404 ,n2321 ,n274);
    or g73(n301 ,n293 ,n300);
    or g74(n772 ,n2327 ,n623);
    nor g75(n172 ,n44 ,n171);
    nand g76(n2614 ,n4[17] ,n2610);
    nand g77(n1570 ,n2[117] ,n1258);
    nand g78(n1310 ,n3[14] ,n915);
    xnor g79(n77 ,n2481 ,n2417);
    not g80(n275 ,n276);
    not g81(n2553 ,n2552);
    xnor g82(n2341 ,n96 ,n200);
    nand g83(n2725 ,n2723 ,n2724);
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1876), .Q(n3[59]));
    nand g85(n2025 ,n1354 ,n1802);
    nor g86(n2744 ,n2733 ,n2740);
    or g87(n688 ,n2[58] ,n630);
    nor g88(n41 ,n2445 ,n2381);
    nand g89(n1214 ,n5[42] ,n912);
    nand g90(n1590 ,n2[96] ,n1256);
    nand g91(n397 ,n2348 ,n274);
    or g92(n1365 ,n2[68] ,n1265);
    nand g93(n1500 ,n798 ,n1305);
    nor g94(n836 ,n5[52] ,n644);
    nor g95(n34 ,n2472 ,n2408);
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1975), .Q(n4[62]));
    nand g97(n1944 ,n1169 ,n1696);
    nor g98(n22 ,n2442 ,n2378);
    nand g99(n1301 ,n3[20] ,n909);
    nand g100(n1026 ,n343 ,n593);
    nand g101(n2452 ,n2142 ,n2126);
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1911), .Q(n3[34]));
    nor g103(n522 ,n7[7] ,n451);
    nand g104(n1577 ,n2[109] ,n1259);
    nand g105(n1212 ,n5[43] ,n912);
    nand g106(n1564 ,n2[123] ,n1257);
    or g107(n845 ,n5[2] ,n631);
    nand g108(n1041 ,n398 ,n570);
    xnor g109(n2627 ,n4[21] ,n2622);
    nand g110(n2467 ,n2141 ,n2079);
    nand g111(n2140 ,n7[7] ,n2043);
    nand g112(n406 ,n2281 ,n312);
    nand g113(n2430 ,n2057 ,n2061);
    nand g114(n1239 ,n5[33] ,n922);
    or g115(n1362 ,n2[70] ,n1265);
    xnor g116(n75 ,n2482 ,n2418);
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2807), .Q(n7[23]));
    nand g118(n1192 ,n5[59] ,n914);
    nor g119(n242 ,n57 ,n241);
    nor g120(n1841 ,n1041 ,n1774);
    nand g121(n2053 ,n2[81] ,n6[1]);
    or g122(n923 ,n456 ,n620);
    nand g123(n1092 ,n2[57] ,n562);
    nand g124(n1086 ,n2[61] ,n562);
    nand g125(n2715 ,n2714 ,n2713);
    nand g126(n2215 ,n2[111] ,n6[1]);
    nand g127(n996 ,n317 ,n613);
    nand g128(n352 ,n2358 ,n274);
    nor g129(n2712 ,n2711 ,n2708);
    or g130(n546 ,n3[27] ,n466);
    nand g131(n2599 ,n2543 ,n2597);
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2788), .Q(n9[3]));
    nor g133(n2764 ,n4[58] ,n2762);
    nand g134(n1475 ,n753 ,n1279);
    not g135(n2540 ,n2539);
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1985), .Q(n4[52]));
    xnor g137(n105 ,n2484 ,n2420);
    nand g138(n1483 ,n763 ,n1286);
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1990), .Q(n4[47]));
    nand g140(n402 ,n2302 ,n273);
    nand g141(n2170 ,n2042 ,n3[0]);
    nand g142(n964 ,n397 ,n609);
    nand g143(n1124 ,n2336 ,n652);
    or g144(n542 ,n3[29] ,n466);
    or g145(n538 ,n4[22] ,n468);
    not g146(n2785 ,n9[10]);
    nand g147(n1031 ,n400 ,n475);
    or g148(n1719 ,n1334 ,n1528);
    nand g149(n1999 ,n1394 ,n1842);
    or g150(n1368 ,n2[65] ,n1265);
    nand g151(n1486 ,n768 ,n1291);
    or g152(n552 ,n3[22] ,n468);
    nor g153(n2635 ,n2557 ,n2634);
    nor g154(n247 ,n92 ,n246);
    or g155(n2706 ,n4[43] ,n2702);
    nor g156(n51 ,n2494 ,n2430);
    or g157(n2581 ,n4[8] ,n2580);
    nand g158(n462 ,n308 ,n380);
    xor g159(n2813 ,n2[6] ,n9[6]);
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1969), .Q(n3[51]));
    nor g161(n1833 ,n1028 ,n1766);
    xnor g162(n2332 ,n85 ,n182);
    nand g163(n1180 ,n2[3] ,n657);
    nor g164(n1851 ,n1059 ,n1786);
    nand g165(n875 ,n4[15] ,n558);
    nand g166(n1019 ,n387 ,n618);
    nand g167(n2122 ,n2[78] ,n6[1]);
    or g168(n533 ,n3[34] ,n465);
    nor g169(n1598 ,n826 ,n1408);
    nor g170(n150 ,n54 ,n149);
    nand g171(n2435 ,n2173 ,n2144);
    nand g172(n1040 ,n4[39] ,n656);
    xnor g173(n95 ,n2438 ,n2374);
    nand g174(n2493 ,n2242 ,n2151);
    nand g175(n2141 ,n7[31] ,n2043);
    nor g176(n234 ,n23 ,n233);
    xnor g177(n2363 ,n132 ,n244);
    nand g178(n2002 ,n1398 ,n1845);
    or g179(n615 ,n4[36] ,n465);
    nand g180(n859 ,n393 ,n545);
    nand g181(n419 ,n2263 ,n273);
    nand g182(n1081 ,n2352 ,n651);
    nand g183(n1980 ,n1375 ,n1823);
    nand g184(n638 ,n7[31] ,n450);
    not g185(n2786 ,n9[19]);
    or g186(n1360 ,n2[72] ,n1262);
    nor g187(n1603 ,n799 ,n1413);
    xor g188(n2294 ,n2734 ,n4[50]);
    nand g189(n1959 ,n1121 ,n1710);
    nand g190(n1784 ,n1592 ,n1056);
    not g191(n2702 ,n2701);
    nor g192(n233 ,n97 ,n232);
    nor g193(n1815 ,n906 ,n1748);
    nand g194(n2458 ,n2142 ,n2105);
    nand g195(n2108 ,n2042 ,n3[44]);
    nand g196(n1960 ,n1180 ,n1711);
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1945), .Q(n5[12]));
    nor g198(n712 ,n5[63] ,n645);
    nor g199(n250 ,n32 ,n249);
    nand g200(n624 ,n7[15] ,n461);
    nand g201(n392 ,n2255 ,n273);
    nand g202(n2660 ,n2659 ,n2658);
    nand g203(n327 ,n2253 ,n312);
    xnor g204(n73 ,n2499 ,n2435);
    xnor g205(n106 ,n2443 ,n2379);
    nand g206(n2163 ,n2[74] ,n6[1]);
    nand g207(n2461 ,n2141 ,n2066);
    nor g208(n1687 ,n797 ,n1501);
    nand g209(n1534 ,n2[89] ,n1252);
    nand g210(n1552 ,n2[71] ,n1255);
    nor g211(n2246 ,n2569 ,n2571);
    nand g212(n1455 ,n1210 ,n1198);
    nand g213(n2099 ,n2043 ,n3[23]);
    nand g214(n2031 ,n1348 ,n1796);
    nor g215(n166 ,n17 ,n165);
    xnor g216(n111 ,n2446 ,n2382);
    nand g217(n391 ,n2354 ,n274);
    or g218(n1379 ,n2[117] ,n1264);
    nand g219(n2064 ,n2[85] ,n6[1]);
    nand g220(n951 ,n446 ,n519);
    nand g221(n2686 ,n7[39] ,n2683);
    not g222(n2721 ,n2720);
    nor g223(n1844 ,n995 ,n1777);
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1887), .Q(n5[34]));
    nand g225(n1315 ,n3[2] ,n911);
    nor g226(n2705 ,n2704 ,n2701);
    not g227(n2527 ,n4[1]);
    nand g228(n2208 ,n2[50] ,n6[1]);
    nor g229(n2593 ,n2592 ,n2590);
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1923), .Q(n5[20]));
    nor g231(n203 ,n101 ,n202);
    nand g232(n1451 ,n718 ,n1241);
    nand g233(n1270 ,n3[38] ,n918);
    nand g234(n1525 ,n719 ,n1323);
    nand g235(n417 ,n2310 ,n311);
    nor g236(n202 ,n18 ,n201);
    nand g237(n2463 ,n2141 ,n2069);
    nand g238(n1324 ,n5[9] ,n913);
    nand g239(n376 ,n2335 ,n274);
    nand g240(n2487 ,n2243 ,n2132);
    or g241(n1361 ,n2[71] ,n1265);
    nor g242(n30 ,n2448 ,n2384);
    nand g243(n1160 ,n2[18] ,n628);
    nand g244(n1281 ,n5[23] ,n916);
    or g245(n829 ,n2[0] ,n632);
    or g246(n742 ,n2[37] ,n643);
    nor g247(n183 ,n85 ,n182);
    xnor g248(n107 ,n2472 ,n2408);
    nor g249(n157 ,n113 ,n156);
    nor g250(n692 ,n5[39] ,n641);
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2787), .Q(n9[12]));
    nand g252(n2410 ,n2234 ,n2229);
    nand g253(n384 ,n2279 ,n274);
    nand g254(n1562 ,n2[125] ,n1257);
    nand g255(n2225 ,n2[11] ,n6[1]);
    or g256(n798 ,n2[17] ,n634);
    nor g257(n1694 ,n999 ,n1506);
    nand g258(n1184 ,n2[0] ,n657);
    nand g259(n433 ,n2261 ,n312);
    nand g260(n2000 ,n1396 ,n1843);
    nand g261(n2417 ,n2123 ,n2115);
    nand g262(n1731 ,n1541 ,n868);
    nand g263(n962 ,n430 ,n585);
    not g264(n311 ,n276);
    nand g265(n1189 ,n2309 ,n648);
    not g266(n1190 ,n1064);
    nor g267(n1824 ,n1015 ,n1757);
    nand g268(n1243 ,n3[45] ,n921);
    nor g269(n1659 ,n746 ,n1470);
    nand g270(n2074 ,n2[94] ,n6[1]);
    dff g271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2030), .Q(n4[19]));
    xnor g272(n2334 ,n81 ,n186);
    nand g273(n2107 ,n2[105] ,n6[1]);
    nand g274(n2390 ,n2095 ,n2058);
    not g275(n2757 ,n2756);
    or g276(n608 ,n3[13] ,n467);
    nand g277(n1245 ,n3[43] ,n921);
    or g278(n706 ,n2343 ,n627);
    xnor g279(n2261 ,n2612 ,n4[17]);
    nor g280(n188 ,n59 ,n187);
    nand g281(n2124 ,n2[17] ,n6[1]);
    nand g282(n1046 ,n4[26] ,n647);
    nand g283(n357 ,n2252 ,n273);
    nand g284(n622 ,n7[47] ,n461);
    nand g285(n1064 ,n2308 ,n648);
    nand g286(n967 ,n373 ,n529);
    nand g287(n1550 ,n2[73] ,n1254);
    nand g288(n854 ,n4[25] ,n647);
    nand g289(n1311 ,n5[12] ,n913);
    nand g290(n2763 ,n4[57] ,n2760);
    not g291(n2513 ,n4[18]);
    nand g292(n2098 ,n2[101] ,n6[1]);
    nand g293(n972 ,n4[33] ,n656);
    dff g294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2789), .Q(n9[8]));
    or g295(n661 ,n2339 ,n625);
    nor g296(n2801 ,n2781 ,n1);
    nor g297(n1252 ,n7[31] ,n907);
    nand g298(n1901 ,n1123 ,n1652);
    nor g299(n187 ,n81 ,n186);
    not g300(n2778 ,n9[2]);
    nand g301(n336 ,n2362 ,n311);
    nand g302(n2213 ,n2[68] ,n6[1]);
    nor g303(n249 ,n104 ,n248);
    dff g304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1877), .Q(n3[58]));
    nand g305(n1579 ,n2[107] ,n1259);
    nor g306(n1647 ,n959 ,n1458);
    xnor g307(n2268 ,n2558 ,n2634);
    nand g308(n2191 ,n2043 ,n3[34]);
    nand g309(n1891 ,n1110 ,n1641);
    not g310(n907 ,n908);
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1864), .Q(n5[46]));
    or g312(n913 ,n452 ,n547);
    or g313(n738 ,n2310 ,n629);
    or g314(n1394 ,n2[102] ,n1251);
    dff g315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1914), .Q(n5[24]));
    or g316(n487 ,n4[6] ,n469);
    xnor g317(n2362 ,n84 ,n242);
    nand g318(n431 ,n2343 ,n311);
    nand g319(n2077 ,n2[92] ,n6[1]);
    not g320(n2693 ,n2692);
    nand g321(n1238 ,n3[48] ,n923);
    nor g322(n2701 ,n4[42] ,n2699);
    nor g323(n726 ,n5[31] ,n638);
    xor g324(n2264 ,n2624 ,n4[20]);
    nor g325(n820 ,n5[0] ,n631);
    nand g326(n2455 ,n2142 ,n2056);
    nor g327(n170 ,n40 ,n169);
    nor g328(n65 ,n2492 ,n2428);
    nand g329(n1289 ,n3[27] ,n917);
    nand g330(n1519 ,n686 ,n1320);
    nand g331(n1130 ,n2[36] ,n559);
    or g332(n508 ,n3[55] ,n470);
    nand g333(n2546 ,n4[12] ,n7[15]);
    or g334(n302 ,n6[0] ,n301);
    or g335(n747 ,n2[35] ,n643);
    nand g336(n1515 ,n825 ,n1287);
    nor g337(n1259 ,n7[47] ,n907);
    nand g338(n1195 ,n5[56] ,n914);
    nand g339(n1529 ,n727 ,n1335);
    nand g340(n1750 ,n1561 ,n1060);
    nand g341(n2001 ,n1397 ,n1844);
    nand g342(n1148 ,n2[25] ,n556);
    nand g343(n1078 ,n2355 ,n651);
    nand g344(n341 ,n2366 ,n312);
    nand g345(n1582 ,n2[104] ,n1259);
    nor g346(n1700 ,n819 ,n1511);
    nand g347(n1317 ,n5[8] ,n913);
    nand g348(n943 ,n348 ,n511);
    nand g349(n1316 ,n3[9] ,n915);
    nand g350(n1957 ,n1179 ,n1708);
    nand g351(n1513 ,n724 ,n1316);
    dff g352(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2029), .Q(n4[18]));
    nand g353(n2184 ,n2[3] ,n6[1]);
    nand g354(n1892 ,n1111 ,n1643);
    nand g355(n1047 ,n4[36] ,n656);
    nand g356(n1978 ,n1374 ,n1821);
    nor g357(n1664 ,n756 ,n1475);
    nand g358(n899 ,n330 ,n490);
    nand g359(n953 ,n4[31] ,n647);
    not g360(n279 ,n2503);
    not g361(n2584 ,n2583);
    nor g362(n716 ,n5[33] ,n641);
    or g363(n1369 ,n2[64] ,n1265);
    nand g364(n1193 ,n5[58] ,n914);
    xor g365(n2269 ,n2639 ,n4[25]);
    nand g366(n472 ,n306 ,n381);
    nor g367(n1613 ,n676 ,n1423);
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1857), .Q(n5[55]));
    nand g369(n2049 ,n2042 ,n3[39]);
    nand g370(n2211 ,n2[36] ,n6[1]);
    nand g371(n1125 ,n2[39] ,n559);
    nand g372(n140 ,n71 ,n139);
    nor g373(n196 ,n68 ,n195);
    nor g374(n2529 ,n2507 ,n4[46]);
    nor g375(n246 ,n12 ,n245);
    nand g376(n2625 ,n2526 ,n2622);
    or g377(n139 ,n95 ,n138);
    nand g378(n1286 ,n3[28] ,n917);
    or g379(n695 ,n2346 ,n627);
    nand g380(n1004 ,n340 ,n514);
    nor g381(n2722 ,n2721 ,n2718);
    nand g382(n1224 ,n3[5] ,n911);
    or g383(n677 ,n2351 ,n622);
    nand g384(n2103 ,n2[39] ,n6[1]);
    nand g385(n445 ,n2254 ,n275);
    nand g386(n1573 ,n2[114] ,n1258);
    nand g387(n2626 ,n4[21] ,n2623);
    nor g388(n219 ,n130 ,n218);
    or g389(n610 ,n3[14] ,n467);
    nor g390(n154 ,n41 ,n153);
    nand g391(n2414 ,n2072 ,n2068);
    nand g392(n1883 ,n1095 ,n1628);
    nor g393(n19 ,n2476 ,n2412);
    buf g394(n6[2] ,n2040);
    nor g395(n1816 ,n927 ,n1749);
    nor g396(n68 ,n2466 ,n2402);
    nor g397(n1690 ,n803 ,n1502);
    nand g398(n1467 ,n740 ,n1270);
    dff g399(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1889), .Q(n3[48]));
    nor g400(n1618 ,n932 ,n1428);
    nor g401(n2534 ,n2517 ,n7[63]);
    nand g402(n2665 ,n2662 ,n2663);
    dff g403(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1920), .Q(n3[28]));
    nand g404(n2621 ,n4[19] ,n2617);
    nor g405(n769 ,n5[20] ,n636);
    nand g406(n1217 ,n3[61] ,n924);
    nor g407(n169 ,n123 ,n168);
    nand g408(n1769 ,n1578 ,n1032);
    nand g409(n1909 ,n1131 ,n1660);
    nand g410(n2227 ,n2[51] ,n6[1]);
    nand g411(n2425 ,n2071 ,n2067);
    nor g412(n2623 ,n2522 ,n2621);
    nand g413(n1141 ,n2[29] ,n556);
    nand g414(n307 ,n2039 ,n303);
    xnor g415(n2371 ,n73 ,n260);
    nand g416(n1218 ,n3[60] ,n924);
    nand g417(n892 ,n357 ,n544);
    dff g418(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1930), .Q(n3[23]));
    or g419(n2672 ,n4[35] ,n2668);
    nand g420(n2438 ,n2140 ,n2230);
    nand g421(n2234 ,n2042 ,n3[38]);
    nand g422(n1854 ,n1063 ,n1599);
    or g423(n566 ,n4[14] ,n467);
    nor g424(n38 ,n2460 ,n2396);
    or g425(n504 ,n3[57] ,n463);
    nand g426(n2532 ,n4[11] ,n2516);
    nand g427(n409 ,n2244 ,n273);
    nand g428(n993 ,n324 ,n597);
    dff g429(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1935), .Q(n5[16]));
    nand g430(n1755 ,n1565 ,n865);
    or g431(n1363 ,n2[69] ,n1265);
    nor g432(n1670 ,n761 ,n1482);
    nor g433(n1632 ,n937 ,n1443);
    nand g434(n1965 ,n1184 ,n1717);
    nand g435(n2085 ,n2[96] ,n6[1]);
    nand g436(n1112 ,n2340 ,n653);
    dff g437(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1950), .Q(n3[9]));
    nand g438(n2078 ,n2042 ,n3[15]);
    nand g439(n2083 ,n2[88] ,n6[1]);
    nand g440(n1302 ,n3[19] ,n909);
    nand g441(n1738 ,n1548 ,n885);
    nor g442(n2583 ,n7[15] ,n2581);
    nand g443(n1531 ,n849 ,n1339);
    nand g444(n428 ,n2258 ,n273);
    nand g445(n1000 ,n404 ,n608);
    not g446(n2743 ,n2742);
    nand g447(n383 ,n2274 ,n275);
    nand g448(n2066 ,n2[89] ,n6[1]);
    xor g449(n2811 ,n2[7] ,n9[7]);
    xor g450(n2299 ,n4[55] ,n2752);
    nand g451(n1449 ,n715 ,n1239);
    nand g452(n1266 ,n7[63] ,n908);
    nor g453(n678 ,n304 ,n619);
    nand g454(n1989 ,n1384 ,n1832);
    nor g455(n1721 ,n722 ,n1529);
    dff g456(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1993), .Q(n4[44]));
    or g457(n785 ,n2325 ,n623);
    or g458(n2789 ,n9[9] ,n1);
    nand g459(n1237 ,n3[49] ,n923);
    nand g460(n2556 ,n4[32] ,n7[39]);
    not g461(n2709 ,n2708);
    or g462(n1403 ,n2[95] ,n1260);
    nand g463(n2168 ,n2[0] ,n6[1]);
    or g464(n1370 ,n2[114] ,n1264);
    nand g465(n2420 ,n2176 ,n2166);
    nor g466(n1639 ,n950 ,n1450);
    nor g467(n1812 ,n899 ,n1745);
    nand g468(n2669 ,n2666 ,n2664);
    dff g469(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2017), .Q(n4[6]));
    nand g470(n1961 ,n1178 ,n1712);
    nor g471(n666 ,n5[49] ,n644);
    nand g472(n896 ,n345 ,n487);
    nand g473(n994 ,n4[59] ,n564);
    or g474(n2664 ,n4[33] ,n2663);
    nand g475(n1752 ,n1562 ,n887);
    nor g476(n721 ,n5[32] ,n641);
    nand g477(n1548 ,n2[75] ,n1254);
    nand g478(n2152 ,n2[122] ,n6[1]);
    nand g479(n1052 ,n366 ,n579);
    or g480(n536 ,n3[33] ,n465);
    nand g481(n1566 ,n2[121] ,n1257);
    nand g482(n2707 ,n4[43] ,n2704);
    or g483(n545 ,n4[23] ,n468);
    nand g484(n2036 ,n1342 ,n1791);
    nand g485(n1104 ,n2343 ,n653);
    nor g486(n381 ,n305 ,n314);
    nand g487(n1303 ,n3[40] ,n921);
    nand g488(n2379 ,n2207 ,n2206);
    nand g489(n1894 ,n1113 ,n1692);
    nand g490(n313 ,n6[0] ,n308);
    nand g491(n1418 ,n663 ,n1202);
    nand g492(n1541 ,n2[82] ,n1253);
    dff g493(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2810), .Q(n7[39]));
    nand g494(n2037 ,n1388 ,n1790);
    nand g495(n1516 ,n728 ,n1268);
    nor g496(n2729 ,n2727 ,n2726);
    not g497(n281 ,n2506);
    nand g498(n2150 ,n2[47] ,n6[1]);
    nor g499(n194 ,n11 ,n193);
    nor g500(n1685 ,n788 ,n1495);
    xnor g501(n129 ,n2456 ,n2392);
    nor g502(n2671 ,n2670 ,n2667);
    dff g503(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2024), .Q(n4[13]));
    xnor g504(n119 ,n2475 ,n2411);
    nand g505(n1059 ,n333 ,n498);
    dff g506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1872), .Q(n3[62]));
    or g507(n1372 ,n2[127] ,n1266);
    nand g508(n2607 ,n4[16] ,n2605);
    or g509(n2787 ,n9[13] ,n1);
    dff g510(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1785), .Q(n5[3]));
    nand g511(n1867 ,n1080 ,n1612);
    dff g512(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1871), .Q(n3[63]));
    nand g513(n1951 ,n1070 ,n1700);
    or g514(n563 ,n454 ,n380);
    nand g515(n444 ,n2284 ,n311);
    nor g516(n254 ,n70 ,n253);
    dff g517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2008), .Q(n4[29]));
    nor g518(n2732 ,n2524 ,n2728);
    or g519(n729 ,n2[43] ,n640);
    nand g520(n1982 ,n1377 ,n1825);
    nand g521(n2228 ,n2[65] ,n6[1]);
    nand g522(n1586 ,n2[100] ,n1256);
    dff g523(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2011), .Q(n4[0]));
    dff g524(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2025), .Q(n4[14]));
    nand g525(n326 ,n2260 ,n312);
    nor g526(n1809 ,n893 ,n1742);
    nand g527(n1862 ,n1073 ,n1607);
    nand g528(n1968 ,n1188 ,n1722);
    nand g529(n1861 ,n1072 ,n1606);
    nand g530(n634 ,n7[23] ,n471);
    or g531(n656 ,n455 ,n380);
    nand g532(n1945 ,n1168 ,n1695);
    nand g533(n1751 ,n1593 ,n942);
    nand g534(n1973 ,n1100 ,n1631);
    nand g535(n1441 ,n700 ,n1231);
    xnor g536(n2316 ,n124 ,n150);
    nand g537(n2465 ,n2141 ,n2063);
    nand g538(n2156 ,n2[60] ,n6[1]);
    nand g539(n1077 ,n2315 ,n648);
    xnor g540(n2365 ,n104 ,n248);
    nand g541(n959 ,n356 ,n523);
    nor g542(n1642 ,n726 ,n1456);
    nand g543(n1492 ,n782 ,n1296);
    nor g544(n1691 ,n997 ,n1503);
    nand g545(n1151 ,n2326 ,n650);
    nor g546(n244 ,n31 ,n243);
    nand g547(n443 ,n2308 ,n311);
    nor g548(n1619 ,n685 ,n1429);
    nand g549(n1744 ,n1554 ,n897);
    or g550(n670 ,n2365 ,n646);
    nand g551(n2024 ,n1355 ,n1803);
    nand g552(n1484 ,n764 ,n1288);
    nand g553(n1914 ,n1135 ,n1664);
    nor g554(n48 ,n2464 ,n2400);
    nand g555(n1136 ,n2[32] ,n559);
    dff g556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1866), .Q(n5[47]));
    nand g557(n1783 ,n1591 ,n953);
    xnor g558(n116 ,n2487 ,n2423);
    or g559(n697 ,n2355 ,n622);
    dff g560(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n448), .Q(n2040));
    dff g561(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n285), .Q(n8[3]));
    or g562(n667 ,n2356 ,n626);
    nand g563(n636 ,n7[23] ,n450);
    nor g564(n165 ,n120 ,n164);
    nor g565(n1710 ,n904 ,n1520);
    nor g566(n379 ,n1 ,n313);
    dff g567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2033), .Q(n4[22]));
    nor g568(n1820 ,n1007 ,n1753);
    nand g569(n1294 ,n3[24] ,n917);
    not g570(n2728 ,n2727);
    nand g571(n1153 ,n2[22] ,n628);
    xnor g572(n112 ,n2497 ,n2433);
    nand g573(n1205 ,n3[4] ,n911);
    not g574(n91 ,n90);
    or g575(n531 ,n3[35] ,n465);
    nand g576(n2404 ,n2171 ,n2167);
    or g577(n523 ,n3[43] ,n464);
    or g578(n2685 ,n2551 ,n2682);
    nand g579(n295 ,n8[0] ,n8[1]);
    or g580(n822 ,n2317 ,n624);
    not g581(n283 ,n2500);
    nand g582(n2018 ,n1361 ,n1809);
    dff g583(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2805), .Q(n9[14]));
    dff g584(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1919), .Q(n5[22]));
    nor g585(n286 ,n279 ,n1);
    nand g586(n1524 ,n835 ,n1206);
    dff g587(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2021), .Q(n4[10]));
    nand g588(n1758 ,n1568 ,n1016);
    nor g589(n689 ,n5[47] ,n635);
    nand g590(n364 ,n2272 ,n275);
    or g591(n744 ,n2[36] ,n643);
    nand g592(n1908 ,n1130 ,n1658);
    nor g593(n292 ,n281 ,n1);
    nand g594(n1268 ,n3[6] ,n911);
    nand g595(n2071 ,n2043 ,n3[53]);
    nand g596(n1956 ,n1177 ,n1706);
    nand g597(n2555 ,n4[56] ,n7[63]);
    or g598(n1718 ,n1333 ,n1532);
    dff g599(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1989), .Q(n4[48]));
    nand g600(n1208 ,n5[46] ,n912);
    or g601(n918 ,n455 ,n620);
    nand g602(n2008 ,n1405 ,n1851);
    nor g603(n838 ,n5[30] ,n638);
    nand g604(n1158 ,n2[19] ,n628);
    nand g605(n1122 ,n2337 ,n652);
    nand g606(n1073 ,n2358 ,n654);
    nand g607(n1907 ,n1129 ,n1659);
    nand g608(n349 ,n2275 ,n274);
    nor g609(n1400 ,n840 ,n1329);
    nand g610(n437 ,n2256 ,n311);
    nand g611(n2580 ,n7[7] ,n2579);
    dff g612(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1836), .Q(n3[54]));
    nand g613(n407 ,n2286 ,n311);
    dff g614(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1868), .Q(n5[44]));
    nand g615(n426 ,n2356 ,n312);
    xnor g616(n2345 ,n110 ,n208);
    nand g617(n1970 ,n1101 ,n1633);
    nor g618(n717 ,n5[48] ,n644);
    nand g619(n2106 ,n2043 ,n3[54]);
    nand g620(n1053 ,n4[50] ,n658);
    or g621(n766 ,n2[27] ,n637);
    nor g622(n651 ,n7[47] ,n462);
    xnor g623(n102 ,n2452 ,n2388);
    nor g624(n556 ,n7[31] ,n472);
    xnor g625(n2500 ,n8[7] ,n272);
    nand g626(n1788 ,n1550 ,n889);
    nand g627(n2586 ,n2582 ,n2581);
    xor g628(n2277 ,n2665 ,n4[33]);
    or g629(n614 ,n3[18] ,n468);
    nor g630(n191 ,n76 ,n190);
    nand g631(n2663 ,n2537 ,n2660);
    nor g632(n649 ,n7[15] ,n462);
    or g633(n515 ,n3[50] ,n470);
    nor g634(n1680 ,n985 ,n1492);
    nor g635(n288 ,n282 ,n1);
    not g636(n266 ,n265);
    nand g637(n2724 ,n4[48] ,n2722);
    nor g638(n10 ,n2483 ,n2419);
    nor g639(n160 ,n30 ,n159);
    nand g640(n2710 ,n2707 ,n2706);
    dff g641(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1998), .Q(n4[39]));
    nand g642(n2173 ,n2043 ,n3[63]);
    nand g643(n2133 ,n2[116] ,n6[1]);
    nand g644(n2070 ,n2[20] ,n6[1]);
    nand g645(n2205 ,n2043 ,n3[62]);
    nand g646(n138 ,n14 ,n137);
    nor g647(n40 ,n2453 ,n2389);
    nor g648(n252 ,n51 ,n251);
    nand g649(n932 ,n441 ,n499);
    xnor g650(n2354 ,n75 ,n226);
    xnor g651(n108 ,n2486 ,n2422);
    nor g652(n2746 ,n4[51] ,n2738);
    nand g653(n904 ,n319 ,n580);
    nor g654(n184 ,n38 ,n183);
    nand g655(n1853 ,n1176 ,n1598);
    nor g656(n2678 ,n2677 ,n2674);
    nand g657(n1865 ,n1076 ,n1609);
    nor g658(n1703 ,n1013 ,n1513);
    dff g659(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1892), .Q(n3[46]));
    nor g660(n1678 ,n984 ,n1490);
    nand g661(n991 ,n395 ,n616);
    nand g662(n1060 ,n4[63] ,n564);
    dff g663(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2019), .Q(n4[8]));
    nand g664(n1102 ,n2[52] ,n561);
    nand g665(n2186 ,n2043 ,n3[3]);
    nor g666(n146 ,n21 ,n145);
    not g667(n2675 ,n2674);
    nand g668(n2478 ,n2138 ,n2109);
    or g669(n481 ,n3[9] ,n467);
    dff g670(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1861), .Q(n5[51]));
    nor g671(n18 ,n2469 ,n2405);
    xnor g672(n126 ,n2454 ,n2390);
    nand g673(n2695 ,n2507 ,n2691);
    nand g674(n1746 ,n1556 ,n900);
    dff g675(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2007), .Q(n4[30]));
    nand g676(n2689 ,n4[39] ,n2685);
    xnor g677(n115 ,n2474 ,n2410);
    nand g678(n1054 ,n390 ,n535);
    nor g679(n1611 ,n804 ,n1421);
    or g680(n613 ,n3[17] ,n468);
    nand g681(n928 ,n351 ,n489);
    nand g682(n2231 ,n2[12] ,n6[1]);
    nand g683(n2128 ,n2043 ,n3[27]);
    nand g684(n975 ,n328 ,n537);
    not g685(n2523 ,n4[58]);
    xnor g686(n2357 ,n97 ,n232);
    nand g687(n2730 ,n2524 ,n2726);
    nor g688(n2592 ,n2521 ,n2589);
    or g689(n1354 ,n2[78] ,n1262);
    nand g690(n1216 ,n3[62] ,n924);
    nor g691(n1852 ,n1061 ,n1787);
    nor g692(n178 ,n53 ,n177);
    nand g693(n643 ,n7[39] ,n471);
    nand g694(n1773 ,n1582 ,n1037);
    xnor g695(n2364 ,n92 ,n246);
    nand g696(n1013 ,n418 ,n481);
    nand g697(n961 ,n432 ,n525);
    nand g698(n2716 ,n2545 ,n2715);
    nor g699(n32 ,n2493 ,n2429);
    xnor g700(n2342 ,n101 ,n202);
    nand g701(n1902 ,n1124 ,n1654);
    nand g702(n1182 ,n2313 ,n648);
    nand g703(n1232 ,n3[52] ,n923);
    nor g704(n11 ,n2465 ,n2401);
    or g705(n518 ,n4[21] ,n468);
    or g706(n811 ,n2[13] ,n633);
    nand g707(n1456 ,n661 ,n1246);
    nor g708(n1790 ,n853 ,n1723);
    nand g709(n891 ,n4[8] ,n558);
    nand g710(n1976 ,n1373 ,n1819);
    dff g711(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1933), .Q(n3[20]));
    nand g712(n2138 ,n7[47] ,n2043);
    or g713(n817 ,n2366 ,n646);
    xnor g714(n2307 ,n2776 ,n4[63]);
    nand g715(n2393 ,n2082 ,n2076);
    nor g716(n210 ,n29 ,n209);
    nand g717(n416 ,n2282 ,n311);
    nand g718(n860 ,n4[22] ,n565);
    nor g719(n209 ,n110 ,n208);
    or g720(n664 ,n2[4] ,n632);
    nand g721(n900 ,n4[3] ,n563);
    nand g722(n1940 ,n1163 ,n1690);
    dff g723(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1967), .Q(n5[62]));
    nand g724(n2159 ,n2[125] ,n6[1]);
    nand g725(n2003 ,n1399 ,n1846);
    nand g726(n1186 ,n2371 ,n655);
    xnor g727(n2313 ,n103 ,n144);
    nor g728(n238 ,n35 ,n237);
    or g729(n846 ,n2340 ,n627);
    nand g730(n321 ,n2280 ,n311);
    xnor g731(n87 ,n2468 ,n2404);
    or g732(n2790 ,n9[8] ,n1);
    not g733(n2736 ,n2735);
    nand g734(n2116 ,n2[109] ,n6[1]);
    xnor g735(n2352 ,n83 ,n222);
    dff g736(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1928), .Q(n5[19]));
    nor g737(n1683 ,n989 ,n1494);
    or g738(n711 ,n2342 ,n627);
    nand g739(n1997 ,n1392 ,n1840);
    xnor g740(n74 ,n2465 ,n2401);
    xnor g741(n109 ,n2445 ,n2381);
    nand g742(n1741 ,n1551 ,n891);
    or g743(n575 ,n3[3] ,n469);
    nand g744(n1565 ,n2[122] ,n1257);
    nor g745(n212 ,n61 ,n211);
    nor g746(n152 ,n24 ,n151);
    nand g747(n857 ,n411 ,n602);
    nand g748(n389 ,n2365 ,n274);
    or g749(n828 ,n5[4] ,n631);
    nand g750(n1167 ,n2[14] ,n557);
    nand g751(n322 ,n2259 ,n275);
    nor g752(n1823 ,n1012 ,n1756);
    nand g753(n1422 ,n673 ,n1209);
    nand g754(n2214 ,n2043 ,n3[8]);
    nor g755(n1635 ,n946 ,n1446);
    nand g756(n1530 ,n672 ,n1337);
    xnor g757(n110 ,n2473 ,n2409);
    or g758(n501 ,n3[60] ,n463);
    nor g759(n240 ,n43 ,n239);
    nor g760(n173 ,n128 ,n172);
    dff g761(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1898), .Q(n3[42]));
    nor g762(n45 ,n2477 ,n2413);
    nand g763(n949 ,n329 ,n516);
    not g764(n274 ,n276);
    nand g765(n2400 ,n2135 ,n2134);
    nand g766(n1287 ,n3[7] ,n911);
    nand g767(n1314 ,n3[10] ,n915);
    or g768(n700 ,n2344 ,n627);
    nand g769(n375 ,n2336 ,n273);
    nand g770(n1930 ,n1152 ,n1680);
    nor g771(n159 ,n114 ,n158);
    not g772(n2571 ,n2570);
    nand g773(n2771 ,n2770 ,n2769);
    nand g774(n2240 ,n2[61] ,n6[1]);
    nand g775(n1262 ,n7[15] ,n908);
    nand g776(n340 ,n2306 ,n311);
    dff g777(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n290), .Q(n8[6]));
    nand g778(n1528 ,n738 ,n1331);
    not g779(n2519 ,n4[28]);
    nor g780(n49 ,n2471 ,n2407);
    or g781(n1373 ,n2[125] ,n1266);
    nand g782(n1209 ,n5[45] ,n912);
    xnor g783(n2815 ,n9[11] ,n9[15]);
    nand g784(n862 ,n318 ,n518);
    not g785(n312 ,n276);
    nand g786(n1920 ,n1143 ,n1671);
    nor g787(n305 ,n6[0] ,n303);
    nand g788(n1009 ,n414 ,n483);
    nand g789(n974 ,n339 ,n536);
    or g790(n1364 ,n2[124] ,n1266);
    nand g791(n362 ,n2296 ,n312);
    nor g792(n58 ,n2479 ,n2415);
    or g793(n590 ,n4[25] ,n466);
    dff g794(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2799), .Q(n9[9]));
    or g795(n509 ,n4[41] ,n464);
    or g796(n737 ,n2319 ,n624);
    nand g797(n2424 ,n2054 ,n2046);
    not g798(n2642 ,n2641);
    nand g799(n2442 ,n2140 ,n2197);
    nand g800(n1111 ,n2[46] ,n560);
    nand g801(n2428 ,n2179 ,n2160);
    nand g802(n1132 ,n2333 ,n652);
    nor g803(n765 ,n5[21] ,n636);
    nand g804(n2402 ,n2154 ,n2153);
    nor g805(n1665 ,n975 ,n1477);
    nand g806(n1207 ,n5[47] ,n912);
    or g807(n1399 ,n2[98] ,n1251);
    nand g808(n1936 ,n1160 ,n1688);
    nand g809(n1103 ,n2[51] ,n561);
    nand g810(n1163 ,n2322 ,n649);
    xnor g811(n134 ,n2479 ,n2415);
    xnor g812(n2326 ,n126 ,n170);
    nand g813(n2703 ,n2700 ,n2699);
    nand g814(n1296 ,n3[23] ,n909);
    nor g815(n70 ,n2495 ,n2431);
    nand g816(n2549 ,n4[0] ,n7[7]);
    dff g817(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1991), .Q(n4[46]));
    nor g818(n235 ,n108 ,n234);
    or g819(n2620 ,n4[19] ,n2616);
    or g820(n1382 ,n2[115] ,n1264);
    nand g821(n1464 ,n736 ,n1303);
    nand g822(n1581 ,n2[105] ,n1259);
    dff g823(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1943), .Q(n3[14]));
    nand g824(n1868 ,n1081 ,n1613);
    nand g825(n2497 ,n2242 ,n2159);
    nand g826(n1730 ,n1540 ,n866);
    nand g827(n1408 ,n843 ,n1192);
    nand g828(n884 ,n4[41] ,n639);
    nand g829(n2100 ,n2[54] ,n6[1]);
    nor g830(n557 ,n7[15] ,n472);
    nor g831(n213 ,n119 ,n212);
    nand g832(n2217 ,n2043 ,n3[57]);
    nor g833(n1255 ,n7[7] ,n907);
    nand g834(n1419 ,n667 ,n1204);
    or g835(n1358 ,n2[74] ,n1262);
    dff g836(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2000), .Q(n4[37]));
    nand g837(n1025 ,n342 ,n604);
    nand g838(n1496 ,n794 ,n1299);
    xnor g839(n103 ,n2441 ,n2377);
    xnor g840(n2331 ,n136 ,n180);
    or g841(n1347 ,n2[85] ,n1261);
    nand g842(n1116 ,n2[43] ,n560);
    nor g843(n186 ,n39 ,n185);
    not g844(n261 ,n8[4]);
    nand g845(n1917 ,n1138 ,n1667);
    nor g846(n56 ,n2458 ,n2394);
    nor g847(n2803 ,n2779 ,n1);
    nand g848(n1786 ,n1594 ,n938);
    or g849(n577 ,n4[35] ,n465);
    nand g850(n2125 ,n2[55] ,n6[1]);
    nand g851(n2207 ,n2043 ,n3[7]);
    xor g852(n2812 ,n2[5] ,n9[5]);
    nand g853(n1943 ,n1167 ,n1694);
    nor g854(n1609 ,n717 ,n1419);
    nand g855(n137 ,n72 ,n91);
    nand g856(n434 ,n2264 ,n273);
    nand g857(n1532 ,n684 ,n1336);
    nand g858(n1129 ,n2334 ,n652);
    nand g859(n1558 ,n2[65] ,n1255);
    nor g860(n25 ,n2481 ,n2417);
    nand g861(n1293 ,n3[25] ,n917);
    or g862(n555 ,n4[15] ,n467);
    nor g863(n2798 ,n2783 ,n1);
    nand g864(n2582 ,n4[8] ,n2580);
    dff g865(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1858), .Q(n5[54]));
    nand g866(n950 ,n426 ,n517);
    nand g867(n2091 ,n2042 ,n3[43]);
    nand g868(n1933 ,n1157 ,n1684);
    nand g869(n1888 ,n1109 ,n1640);
    nand g870(n1506 ,n809 ,n1310);
    or g871(n537 ,n3[32] ,n465);
    xor g872(n2266 ,n2630 ,n4[22]);
    nand g873(n2564 ,n2555 ,n2540);
    nand g874(n1753 ,n1563 ,n1002);
    nand g875(n1726 ,n1536 ,n895);
    nand g876(n1462 ,n733 ,n1250);
    or g877(n751 ,n2[33] ,n643);
    nand g878(n2714 ,n4[45] ,n2711);
    nand g879(n1264 ,n7[55] ,n908);
    nand g880(n1114 ,n2[44] ,n560);
    nor g881(n2733 ,n4[50] ,n2730);
    nand g882(n1488 ,n770 ,n1293);
    nand g883(n2431 ,n2117 ,n2093);
    nand g884(n2045 ,n2[77] ,n6[1]);
    nor g885(n606 ,n7[39] ,n451);
    nand g886(n2447 ,n2143 ,n2080);
    or g887(n724 ,n2[9] ,n633);
    xnor g888(n2353 ,n77 ,n224);
    nor g889(n1660 ,n971 ,n1472);
    nand g890(n337 ,n2292 ,n275);
    nand g891(n1188 ,n2369 ,n655);
    nand g892(n2392 ,n2094 ,n2070);
    nand g893(n2484 ,n2243 ,n2210);
    not g894(n2551 ,n2550);
    nand g895(n1880 ,n1094 ,n1626);
    not g896(n2696 ,n2695);
    nand g897(n1491 ,n779 ,n1295);
    or g898(n612 ,n3[16] ,n468);
    nand g899(n2060 ,n2[87] ,n6[1]);
    xor g900(n2272 ,n2651 ,n4[28]);
    nand g901(n2372 ,n2170 ,n2168);
    nand g902(n1263 ,n7[47] ,n908);
    nand g903(n2443 ,n2140 ,n2137);
    nand g904(n1323 ,n3[1] ,n911);
    nand g905(n2223 ,n2042 ,n3[10]);
    xor g906(n2282 ,n4[38] ,n2681);
    nor g907(n304 ,n2039 ,n303);
    nor g908(n2541 ,n4[24] ,n7[31]);
    nand g909(n276 ,n298 ,n306);
    or g910(n2734 ,n2732 ,n2731);
    nor g911(n259 ,n89 ,n258);
    nand g912(n469 ,n7[7] ,n379);
    nand g913(n405 ,n2319 ,n273);
    nand g914(n879 ,n4[13] ,n558);
    nand g915(n1260 ,n7[31] ,n908);
    nand g916(n2082 ,n2043 ,n3[21]);
    nand g917(n1897 ,n1118 ,n1649);
    nand g918(n1075 ,n2[1] ,n657);
    nand g919(n2176 ,n2042 ,n3[48]);
    nand g920(n2180 ,n2[72] ,n6[1]);
    nand g921(n942 ,n4[62] ,n564);
    or g922(n910 ,n452 ,n522);
    nand g923(n1438 ,n696 ,n1227);
    nand g924(n1886 ,n1106 ,n1636);
    or g925(n813 ,n2320 ,n624);
    nand g926(n2171 ,n2042 ,n3[32]);
    or g927(n800 ,n2[8] ,n633);
    or g928(n818 ,n2[59] ,n630);
    nand g929(n1490 ,n777 ,n1294);
    nor g930(n189 ,n78 ,n188);
    dff g931(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1952), .Q(n5[9]));
    nand g932(n1859 ,n1069 ,n1604);
    nand g933(n2046 ,n2[52] ,n6[1]);
    nand g934(n1772 ,n1581 ,n884);
    nand g935(n1213 ,n3[63] ,n924);
    or g936(n553 ,n3[62] ,n463);
    or g937(n544 ,n4[8] ,n467);
    nand g938(n2148 ,n2042 ,n3[29]);
    dff g939(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1907), .Q(n5[26]));
    nand g940(n365 ,n2364 ,n311);
    dff g941(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2038), .Q(n4[27]));
    dff g942(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1949), .Q(n3[10]));
    nand g943(n1733 ,n1543 ,n873);
    nor g944(n2745 ,n2552 ,n2741);
    nand g945(n296 ,n8[2] ,n8[3]);
    nand g946(n874 ,n435 ,n538);
    nand g947(n323 ,n2285 ,n275);
    nor g948(n1668 ,n977 ,n1480);
    nor g949(n168 ,n15 ,n167);
    nand g950(n1561 ,n2[127] ,n1257);
    xnor g951(n2335 ,n78 ,n188);
    nor g952(n185 ,n86 ,n184);
    nor g953(n1695 ,n810 ,n1507);
    nand g954(n1134 ,n2[33] ,n559);
    nand g955(n2380 ,n2214 ,n2212);
    nor g956(n15 ,n2452 ,n2388);
    nor g957(n1831 ,n955 ,n1764);
    or g958(n475 ,n4[45] ,n464);
    or g959(n795 ,n2[18] ,n634);
    nand g960(n1300 ,n3[21] ,n909);
    or g961(n617 ,n3[20] ,n468);
    xnor g962(n2292 ,n2509 ,n2725);
    nor g963(n141 ,n98 ,n140);
    or g964(n786 ,n2[22] ,n634);
    dff g965(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1716), .Q(n5[0]));
    nand g966(n1106 ,n2[49] ,n561);
    nand g967(n966 ,n4[51] ,n658);
    nand g968(n2160 ,n2[56] ,n6[1]);
    nand g969(n2065 ,n2043 ,n3[19]);
    or g970(n713 ,n2360 ,n626);
    nor g971(n1655 ,n967 ,n1467);
    nor g972(n2644 ,n2512 ,n2640);
    nand g973(n934 ,n4[48] ,n658);
    or g974(n2646 ,n4[27] ,n2642);
    dff g975(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2016), .Q(n4[5]));
    or g976(n299 ,n295 ,n296);
    nand g977(n978 ,n374 ,n542);
    nand g978(n1272 ,n3[37] ,n918);
    nor g979(n1838 ,n957 ,n1771);
    nand g980(n334 ,n2309 ,n275);
    nand g981(n1756 ,n1566 ,n880);
    nand g982(n2014 ,n1366 ,n1813);
    nor g983(n669 ,n5[61] ,n645);
    nand g984(n1958 ,n1077 ,n1709);
    nand g985(n1028 ,n331 ,n493);
    xnor g986(n2312 ,n100 ,n142);
    nand g987(n2681 ,n2680 ,n2679);
    or g988(n763 ,n2[28] ,n637);
    nor g989(n650 ,n7[23] ,n462);
    xnor g990(n2561 ,n7[31] ,n4[30]);
    nand g991(n2468 ,n2139 ,n2085);
    nor g992(n1644 ,n807 ,n1505);
    nand g993(n629 ,n7[7] ,n461);
    or g994(n764 ,n2329 ,n623);
    nand g995(n1592 ,n2[94] ,n1252);
    nor g996(n1663 ,n974 ,n1476);
    nand g997(n1048 ,n4[45] ,n639);
    nand g998(n348 ,n2361 ,n274);
    nor g999(n310 ,n297 ,n306);
    nor g1000(n54 ,n2443 ,n2379);
    nand g1001(n2533 ,n7[63] ,n2517);
    nor g1002(n180 ,n56 ,n179);
    nand g1003(n1535 ,n2[88] ,n1252);
    nand g1004(n1522 ,n847 ,n1328);
    nor g1005(n193 ,n74 ,n192);
    or g1006(n672 ,n2369 ,n646);
    or g1007(n1355 ,n2[77] ,n1262);
    nand g1008(n345 ,n2250 ,n273);
    nand g1009(n979 ,n375 ,n543);
    nor g1010(n547 ,n7[15] ,n451);
    nand g1011(n344 ,n2293 ,n274);
    nand g1012(n325 ,n2313 ,n274);
    nand g1013(n1734 ,n1544 ,n875);
    nor g1014(n47 ,n2498 ,n2434);
    nand g1015(n2433 ,n2052 ,n2240);
    nand g1016(n1295 ,n5[18] ,n916);
    nor g1017(n550 ,n7[23] ,n451);
    nand g1018(n2634 ,n2632 ,n2633);
    or g1019(n691 ,n2[57] ,n630);
    dff g1020(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1597), .Q(n5[60]));
    nand g1021(n1094 ,n2[56] ,n562);
    xnor g1022(n2336 ,n76 ,n190);
    nor g1023(n1686 ,n991 ,n1498);
    nand g1024(n2101 ,n2[44] ,n6[1]);
    or g1025(n1383 ,n2[113] ,n1264);
    nor g1026(n2594 ,n2531 ,n2593);
    nand g1027(n1222 ,n3[57] ,n924);
    nor g1028(n1604 ,n734 ,n1414);
    nand g1029(n901 ,n4[28] ,n647);
    xor g1030(n2559 ,n7[63] ,n4[62]);
    nor g1031(n2674 ,n4[36] ,n2672);
    or g1032(n551 ,n3[23] ,n468);
    nor g1033(n43 ,n2488 ,n2424);
    nor g1034(n268 ,n261 ,n267);
    nand g1035(n1863 ,n1074 ,n1608);
    xor g1036(n2304 ,n2771 ,n4[60]);
    or g1037(n825 ,n2[7] ,n632);
    nor g1038(n27 ,n2486 ,n2422);
    dff g1039(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2790), .Q(n9[7]));
    or g1040(n1356 ,n2[76] ,n1262);
    nand g1041(n1194 ,n5[57] ,n914);
    dff g1042(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2806), .Q(n7[31]));
    or g1043(n1374 ,n2[123] ,n1266);
    nand g1044(n883 ,n437 ,n611);
    nand g1045(n1539 ,n2[84] ,n1253);
    or g1046(n782 ,n2[23] ,n634);
    nor g1047(n1797 ,n867 ,n1730);
    nand g1048(n293 ,n8[6] ,n8[7]);
    nand g1049(n2488 ,n2243 ,n2133);
    nor g1050(n671 ,n5[57] ,n645);
    or g1051(n495 ,n4[18] ,n468);
    xnor g1052(n125 ,n2477 ,n2413);
    or g1053(n1380 ,n2[126] ,n1266);
    xor g1054(n2809 ,n2[0] ,n9[0]);
    nand g1055(n2636 ,n2541 ,n2634);
    nor g1056(n306 ,n2039 ,n302);
    dff g1057(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1865), .Q(n5[48]));
    nand g1058(n2413 ,n2059 ,n2118);
    nand g1059(n1244 ,n3[44] ,n921);
    nand g1060(n1560 ,n2[113] ,n1258);
    nor g1061(n562 ,n7[63] ,n472);
    nand g1062(n2483 ,n2138 ,n2215);
    nand g1063(n1329 ,n839 ,n1174);
    nor g1064(n460 ,n7[47] ,n378);
    nor g1065(n1711 ,n1033 ,n1522);
    nand g1066(n2388 ,n2145 ,n2050);
    nor g1067(n2575 ,n2528 ,n2574);
    nor g1068(n2677 ,n2525 ,n2673);
    nor g1069(n791 ,n5[16] ,n636);
    xnor g1070(n122 ,n2488 ,n2424);
    nor g1071(n221 ,n134 ,n220);
    nand g1072(n1499 ,n795 ,n1340);
    or g1073(n521 ,n4[58] ,n463);
    nand g1074(n2456 ,n2142 ,n2111);
    or g1075(n579 ,n4[33] ,n465);
    nor g1076(n2796 ,n2777 ,n1);
    nor g1077(n1650 ,n962 ,n1461);
    nand g1078(n1903 ,n1126 ,n1656);
    xnor g1079(n120 ,n2451 ,n2387);
    dff g1080(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1938), .Q(n5[15]));
    nand g1081(n2080 ,n2[75] ,n6[1]);
    nand g1082(n2166 ,n2[48] ,n6[1]);
    nor g1083(n1803 ,n881 ,n1736);
    or g1084(n1468 ,n2[91] ,n1260);
    nand g1085(n1415 ,n713 ,n1199);
    nor g1086(n61 ,n2474 ,n2410);
    xnor g1087(n2265 ,n2627 ,n2623);
    nand g1088(n2739 ,n2536 ,n2733);
    nand g1089(n350 ,n2328 ,n312);
    nand g1090(n1200 ,n5[51] ,n920);
    nand g1091(n2093 ,n2[59] ,n6[1]);
    or g1092(n506 ,n4[60] ,n463);
    nor g1093(n2670 ,n2511 ,n2666);
    dff g1094(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1931), .Q(n3[22]));
    nand g1095(n1725 ,n1535 ,n856);
    nand g1096(n2381 ,n2220 ,n2218);
    nor g1097(n1666 ,n976 ,n1478);
    or g1098(n513 ,n3[21] ,n468);
    nand g1099(n1288 ,n5[21] ,n916);
    xnor g1100(n117 ,n2449 ,n2385);
    nand g1101(n2426 ,n2106 ,n2100);
    or g1102(n516 ,n3[49] ,n470);
    nand g1103(n2389 ,n2055 ,n2124);
    nand g1104(n464 ,n7[47] ,n379);
    nand g1105(n1276 ,n5[25] ,n919);
    nand g1106(n2385 ,n2088 ,n2239);
    nand g1107(n2030 ,n1349 ,n1797);
    nand g1108(n418 ,n2317 ,n311);
    nand g1109(n2545 ,n4[46] ,n2507);
    nand g1110(n2630 ,n2626 ,n2625);
    nand g1111(n1305 ,n3[17] ,n909);
    dff g1112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2037), .Q(n4[26]));
    dff g1113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1999), .Q(n4[38]));
    nor g1114(n657 ,n7[7] ,n472);
    nand g1115(n1051 ,n436 ,n541);
    nor g1116(n39 ,n2461 ,n2397);
    xnor g1117(n2284 ,n2694 ,n7[47]);
    or g1118(n741 ,n2335 ,n625);
    nand g1119(n2105 ,n2[86] ,n6[1]);
    xnor g1120(n2339 ,n82 ,n196);
    nand g1121(n1545 ,n2[78] ,n1254);
    nand g1122(n976 ,n316 ,n540);
    nor g1123(n797 ,n5[15] ,n621);
    nand g1124(n1575 ,n2[111] ,n1259);
    nor g1125(n1829 ,n963 ,n1762);
    xnor g1126(n2251 ,n4[7] ,n2577);
    nand g1127(n1931 ,n1153 ,n1682);
    nand g1128(n1265 ,n7[7] ,n908);
    nor g1129(n1807 ,n890 ,n1788);
    or g1130(n762 ,n2[29] ,n637);
    nand g1131(n2233 ,n2042 ,n3[12]);
    or g1132(n580 ,n3[4] ,n469);
    nand g1133(n2127 ,n2[113] ,n6[1]);
    dff g1134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1863), .Q(n5[49]));
    dff g1135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1885), .Q(n3[50]));
    nand g1136(n1869 ,n1085 ,n1617);
    nand g1137(n1921 ,n1145 ,n1673);
    dff g1138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1953), .Q(n3[8]));
    nor g1139(n776 ,n5[50] ,n644);
    or g1140(n2723 ,n4[48] ,n2722);
    nand g1141(n332 ,n2359 ,n275);
    nand g1142(n938 ,n4[29] ,n647);
    nand g1143(n1084 ,n2[62] ,n562);
    nor g1144(n2602 ,n4[15] ,n2599);
    dff g1145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n678), .Q(n2039));
    nor g1146(n2622 ,n4[20] ,n2620);
    nand g1147(n1210 ,n5[0] ,n910);
    nand g1148(n876 ,n322 ,n555);
    nand g1149(n1896 ,n1116 ,n1647);
    nand g1150(n1875 ,n1087 ,n1619);
    dff g1151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1900), .Q(n5[29]));
    nor g1152(n1606 ,n659 ,n1416);
    nor g1153(n823 ,n5[58] ,n645);
    nor g1154(n253 ,n99 ,n252);
    nor g1155(n174 ,n46 ,n173);
    nand g1156(n997 ,n399 ,n612);
    nand g1157(n2486 ,n2243 ,n2204);
    dff g1158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2005), .Q(n4[32]));
    xor g1159(n2808 ,n2[1] ,n9[1]);
    nor g1160(n2539 ,n4[56] ,n7[63]);
    nand g1161(n1191 ,n850 ,n1062);
    nor g1162(n55 ,n2482 ,n2418);
    nand g1163(n1069 ,n2361 ,n654);
    nand g1164(n1280 ,n3[32] ,n918);
    nand g1165(n1477 ,n755 ,n1280);
    xnor g1166(n136 ,n2459 ,n2395);
    not g1167(n2783 ,n9[14]);
    nand g1168(n309 ,n6[0] ,n303);
    nand g1169(n314 ,n277 ,n309);
    nand g1170(n1022 ,n371 ,n595);
    dff g1171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2794), .Q(n9[15]));
    nand g1172(n1505 ,n806 ,n1308);
    or g1173(n1716 ,n830 ,n1455);
    nor g1174(n2502 ,n269 ,n271);
    nand g1175(n1967 ,n1187 ,n1721);
    nor g1176(n908 ,n309 ,n619);
    or g1177(n581 ,n4[30] ,n466);
    nand g1178(n1764 ,n1560 ,n944);
    or g1179(n1406 ,n2[92] ,n1260);
    nor g1180(n1198 ,n820 ,n1190);
    nand g1181(n1430 ,n832 ,n1218);
    nand g1182(n1877 ,n1090 ,n1623);
    or g1183(n584 ,n4[27] ,n466);
    nand g1184(n2136 ,n2043 ,n3[55]);
    xnor g1185(n2346 ,n115 ,n210);
    not g1186(n2637 ,n2636);
    dff g1187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1954), .Q(n3[7]));
    nand g1188(n1860 ,n1071 ,n1605);
    nand g1189(n1204 ,n5[48] ,n920);
    nand g1190(n970 ,n358 ,n524);
    nor g1191(n217 ,n125 ,n216);
    nand g1192(n2554 ,n4[14] ,n4[13]);
    or g1193(n827 ,n2[5] ,n632);
    nor g1194(n1629 ,n952 ,n1440);
    nand g1195(n346 ,n2360 ,n274);
    nand g1196(n2183 ,n2043 ,n3[33]);
    nor g1197(n1847 ,n1052 ,n1780);
    nand g1198(n2449 ,n2143 ,n2045);
    nand g1199(n955 ,n344 ,n589);
    nand g1200(n1925 ,n1148 ,n1676);
    nor g1201(n837 ,n5[5] ,n631);
    dff g1202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n289), .Q(n8[7]));
    nand g1203(n2235 ,n2043 ,n3[24]);
    dff g1204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1918), .Q(n3[29]));
    dff g1205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1946), .Q(n3[12]));
    nand g1206(n272 ,n8[6] ,n271);
    xor g1207(n2278 ,n2669 ,n4[34]);
    nor g1208(n1621 ,n690 ,n1433);
    dff g1209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2027), .Q(n4[16]));
    dff g1210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1932), .Q(n3[21]));
    nand g1211(n2418 ,n2194 ,n2131);
    nand g1212(n1215 ,n5[41] ,n912);
    or g1213(n503 ,n3[52] ,n470);
    nand g1214(n1770 ,n1579 ,n1058);
    nor g1215(n28 ,n2446 ,n2382);
    nand g1216(n1164 ,n2[16] ,n628);
    nor g1217(n2631 ,n2629 ,n2628);
    or g1218(n583 ,n4[11] ,n467);
    nand g1219(n1864 ,n1079 ,n1611);
    nor g1220(n1617 ,n682 ,n1426);
    or g1221(n595 ,n4[53] ,n470);
    or g1222(n2737 ,n4[51] ,n2733);
    nor g1223(n1669 ,n978 ,n1481);
    nand g1224(n941 ,n359 ,n508);
    nand g1225(n2069 ,n2[91] ,n6[1]);
    nor g1226(n754 ,n5[55] ,n644);
    xor g1227(n2810 ,n2[4] ,n9[4]);
    or g1228(n663 ,n2357 ,n626);
    nand g1229(n906 ,n424 ,n494);
    nand g1230(n2683 ,n4[38] ,n2681);
    nand g1231(n1322 ,n5[6] ,n910);
    not g1232(n2759 ,n2758);
    nand g1233(n852 ,n442 ,n584);
    or g1234(n512 ,n4[31] ,n466);
    nand g1235(n2406 ,n2191 ,n2188);
    xnor g1236(n128 ,n2455 ,n2391);
    or g1237(n528 ,n3[5] ,n469);
    nand g1238(n1199 ,n5[52] ,n920);
    nand g1239(n1428 ,n683 ,n1217);
    or g1240(n478 ,n3[10] ,n467);
    not g1241(n2509 ,n7[55]);
    nand g1242(n358 ,n2344 ,n274);
    nor g1243(n163 ,n118 ,n162);
    nor g1244(n1830 ,n1026 ,n1763);
    nand g1245(n1919 ,n1142 ,n1670);
    nand g1246(n328 ,n2340 ,n312);
    nand g1247(n2474 ,n2139 ,n2051);
    nand g1248(n1173 ,n2[9] ,n557);
    nand g1249(n2029 ,n1350 ,n1798);
    nand g1250(n1549 ,n2[74] ,n1254);
    nand g1251(n400 ,n2289 ,n275);
    dff g1252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2015), .Q(n4[4]));
    nand g1253(n2086 ,n2[43] ,n6[1]);
    nand g1254(n1234 ,n5[35] ,n922);
    nor g1255(n26 ,n2478 ,n2414);
    nand g1256(n1229 ,n5[37] ,n922);
    nor g1257(n251 ,n121 ,n250);
    dff g1258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1875), .Q(n5[41]));
    nand g1259(n398 ,n2283 ,n274);
    dff g1260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1963), .Q(n3[2]));
    nand g1261(n1923 ,n1147 ,n1675);
    nor g1262(n148 ,n22 ,n147);
    nand g1263(n2104 ,n2[24] ,n6[1]);
    xnor g1264(n2321 ,n117 ,n160);
    nand g1265(n1447 ,n711 ,n1236);
    dff g1266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1966), .Q(n5[63]));
    nor g1267(n821 ,n5[8] ,n621);
    dff g1268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1941), .Q(n3[15]));
    nand g1269(n2020 ,n1359 ,n1807);
    nand g1270(n2567 ,n2547 ,n2535);
    nand g1271(n858 ,n4[27] ,n647);
    or g1272(n2606 ,n4[16] ,n2605);
    nand g1273(n888 ,n4[10] ,n558);
    nand g1274(n1241 ,n3[47] ,n921);
    nand g1275(n2399 ,n2128 ,n2209);
    or g1276(n1357 ,n2[75] ,n1262);
    nand g1277(n2473 ,n2139 ,n2098);
    or g1278(n775 ,n2363 ,n626);
    or g1279(n565 ,n459 ,n380);
    nand g1280(n414 ,n2303 ,n312);
    nand g1281(n347 ,n2329 ,n275);
    nand g1282(n2044 ,n2[15] ,n6[1]);
    xnor g1283(n2349 ,n125 ,n216);
    nand g1284(n626 ,n7[55] ,n461);
    nor g1285(n2755 ,n4[55] ,n2753);
    nand g1286(n894 ,n4[6] ,n563);
    nand g1287(n1410 ,n670 ,n1194);
    nand g1288(n2481 ,n2138 ,n2116);
    nor g1289(n262 ,n8[1] ,n8[0]);
    nand g1290(n2219 ,n2043 ,n3[50]);
    or g1291(n570 ,n4[39] ,n465);
    nor g1292(n2754 ,n2509 ,n2752);
    not g1293(n2784 ,n9[3]);
    or g1294(n1401 ,n2[97] ,n1251);
    nor g1295(n237 ,n116 ,n236);
    nand g1296(n968 ,n370 ,n532);
    or g1297(n684 ,n2309 ,n629);
    dff g1298(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1948), .Q(n5[11]));
    nor g1299(n676 ,n5[44] ,n635);
    nand g1300(n2374 ,n2182 ,n2181);
    nand g1301(n871 ,n326 ,n473);
    nand g1302(n878 ,n428 ,n566);
    dff g1303(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2001), .Q(n4[36]));
    xor g1304(n2288 ,n2710 ,n4[44]);
    nand g1305(n1138 ,n2331 ,n650);
    nand g1306(n1333 ,n680 ,n1189);
    nand g1307(n1963 ,n1181 ,n1713);
    nand g1308(n2153 ,n2[30] ,n6[1]);
    nor g1309(n231 ,n105 ,n230);
    nor g1310(n1848 ,n1054 ,n1782);
    nand g1311(n1995 ,n1390 ,n1838);
    nand g1312(n1233 ,n3[51] ,n923);
    nor g1313(n2726 ,n7[55] ,n2723);
    or g1314(n802 ,n2[16] ,n634);
    nand g1315(n2557 ,n4[24] ,n7[31]);
    nand g1316(n1748 ,n1558 ,n1043);
    nand g1317(n2432 ,n2187 ,n2156);
    xor g1318(n2291 ,n2719 ,n4[47]);
    nand g1319(n2027 ,n1352 ,n1800);
    nor g1320(n451 ,n379 ,n311);
    nand g1321(n1929 ,n1154 ,n1685);
    nor g1322(n1254 ,n7[15] ,n907);
    nand g1323(n646 ,n7[63] ,n461);
    or g1324(n449 ,n306 ,n379);
    or g1325(n609 ,n3[40] ,n464);
    xnor g1326(n2333 ,n86 ,n184);
    dff g1327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1902), .Q(n5[28]));
    nand g1328(n2035 ,n1344 ,n1792);
    nand g1329(n2751 ,n4[54] ,n2745);
    nand g1330(n2416 ,n2108 ,n2101);
    nand g1331(n2384 ,n2233 ,n2231);
    nand g1332(n872 ,n433 ,n480);
    nand g1333(n2096 ,n2[100] ,n6[1]);
    or g1334(n1376 ,n2[120] ,n1266);
    xor g1335(n2270 ,n2643 ,n4[26]);
    nand g1336(n2656 ,n2561 ,n2655);
    nand g1337(n2395 ,n2099 ,n2097);
    nand g1338(n2115 ,n2[45] ,n6[1]);
    nand g1339(n2057 ,n2042 ,n3[58]);
    nand g1340(n1740 ,n1469 ,n858);
    or g1341(n535 ,n4[32] ,n465);
    nand g1342(n2102 ,n2[103] ,n6[1]);
    nand g1343(n343 ,n2294 ,n312);
    nor g1344(n526 ,n7[63] ,n451);
    nand g1345(n1166 ,n2321 ,n649);
    or g1346(n1351 ,n2[81] ,n1261);
    xnor g1347(n130 ,n2478 ,n2414);
    nand g1348(n2475 ,n2139 ,n2102);
    nand g1349(n1018 ,n385 ,n596);
    nand g1350(n2167 ,n2[32] ,n6[1]);
    nand g1351(n1312 ,n3[13] ,n915);
    nand g1352(n1551 ,n2[72] ,n1254);
    nand g1353(n2378 ,n2202 ,n2201);
    or g1354(n718 ,n2[47] ,n640);
    nor g1355(n1713 ,n1035 ,n1523);
    nand g1356(n1589 ,n2[97] ,n1256);
    xnor g1357(n2293 ,n2729 ,n4[49]);
    or g1358(n591 ,n3[6] ,n469);
    nor g1359(n2718 ,n4[47] ,n2716);
    nor g1360(n1649 ,n838 ,n1459);
    dff g1361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2803), .Q(n9[5]));
    nand g1362(n990 ,n350 ,n617);
    nand g1363(n1416 ,n693 ,n1200);
    nor g1364(n1806 ,n981 ,n1739);
    nor g1365(n218 ,n45 ,n217);
    nor g1366(n1658 ,n970 ,n1471);
    dff g1367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2004), .Q(n4[33]));
    nand g1368(n856 ,n4[24] ,n647);
    nand g1369(n1452 ,n720 ,n1242);
    nor g1370(n655 ,n7[63] ,n462);
    nor g1371(n534 ,n7[31] ,n451);
    nor g1372(n167 ,n102 ,n166);
    nor g1373(n2805 ,n2780 ,n1);
    dff g1374(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1929), .Q(n5[17]));
    nand g1375(n2023 ,n1356 ,n1804);
    dff g1376(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2792), .Q(n9[16]));
    nand g1377(n1546 ,n2[77] ,n1254);
    or g1378(n801 ,n2322 ,n624);
    nand g1379(n388 ,n2330 ,n275);
    nand g1380(n2239 ,n2[13] ,n6[1]);
    nand g1381(n2819 ,n2816 ,n2818);
    or g1382(n725 ,n2[44] ,n640);
    nand g1383(n881 ,n369 ,n477);
    nand g1384(n1413 ,n752 ,n1196);
    nor g1385(n162 ,n33 ,n161);
    nand g1386(n387 ,n2316 ,n312);
    nand g1387(n1044 ,n4[37] ,n656);
    xnor g1388(n2361 ,n127 ,n240);
    not g1389(n2514 ,n4[42]);
    nor g1390(n709 ,n5[34] ,n641);
    nand g1391(n1461 ,n732 ,n1249);
    nor g1392(n2605 ,n2602 ,n2604);
    nor g1393(n1846 ,n1051 ,n1779);
    nand g1394(n2550 ,n7[39] ,n2510);
    nand g1395(n1137 ,n2[31] ,n556);
    nand g1396(n1574 ,n2[112] ,n1258);
    dff g1397(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2791), .Q(n9[11]));
    or g1398(n921 ,n460 ,n620);
    nor g1399(n2610 ,n2518 ,n2607);
    nand g1400(n1942 ,n1166 ,n1644);
    nand g1401(n2113 ,n2042 ,n3[25]);
    nand g1402(n1074 ,n2357 ,n654);
    nand g1403(n890 ,n327 ,n554);
    nor g1404(n1256 ,n7[39] ,n907);
    nand g1405(n1327 ,n5[4] ,n910);
    nand g1406(n1308 ,n5[13] ,n913);
    nand g1407(n2411 ,n2049 ,n2103);
    nand g1408(n316 ,n2339 ,n273);
    nand g1409(n2132 ,n2[115] ,n6[1]);
    xor g1410(n2305 ,n2774 ,n4[61]);
    or g1411(n727 ,n2370 ,n646);
    xor g1412(n2290 ,n4[46] ,n2715);
    nand g1413(n1964 ,n1075 ,n1714);
    nand g1414(n2226 ,n2042 ,n3[11]);
    nand g1415(n1593 ,n2[126] ,n1257);
    nor g1416(n256 ,n64 ,n255);
    nor g1417(n453 ,n7[15] ,n378);
    or g1418(n517 ,n3[48] ,n470);
    dff g1419(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1855), .Q(n5[57]));
    or g1420(n745 ,n2334 ,n625);
    nand g1421(n1766 ,n1575 ,n925);
    nor g1422(n1627 ,n941 ,n1438);
    or g1423(n482 ,n4[10] ,n467);
    nor g1424(n2708 ,n4[44] ,n2706);
    nor g1425(n35 ,n2487 ,n2423);
    nor g1426(n743 ,n5[27] ,n638);
    nor g1427(n699 ,n5[37] ,n641);
    nand g1428(n1176 ,n2367 ,n655);
    nand g1429(n2157 ,n2[76] ,n6[1]);
    nor g1430(n2691 ,n4[40] ,n2690);
    nand g1431(n1145 ,n2[27] ,n556);
    nand g1432(n2476 ,n2138 ,n2236);
    nand g1433(n1029 ,n421 ,n588);
    nand g1434(n627 ,n7[39] ,n461);
    nand g1435(n1273 ,n5[26] ,n919);
    nor g1436(n682 ,n5[42] ,n635);
    nand g1437(n1274 ,n3[36] ,n918);
    dff g1438(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2793), .Q(n9[4]));
    nor g1439(n1845 ,n1049 ,n1778);
    nor g1440(n1395 ,n831 ,n1325);
    nor g1441(n1817 ,n1001 ,n1750);
    nand g1442(n1016 ,n4[55] ,n658);
    nand g1443(n1948 ,n1171 ,n1697);
    nor g1444(n1799 ,n872 ,n1732);
    not g1445(n278 ,n2501);
    nand g1446(n1339 ,n5[60] ,n914);
    or g1447(n568 ,n4[26] ,n466);
    or g1448(n806 ,n2321 ,n624);
    dff g1449(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2035), .Q(n4[24]));
    nand g1450(n1953 ,n1140 ,n1704);
    nand g1451(n931 ,n337 ,n587);
    nand g1452(n2195 ,n2[117] ,n6[1]);
    nand g1453(n1187 ,n2370 ,n655);
    nand g1454(n330 ,n2248 ,n275);
    xor g1455(n2274 ,n4[30] ,n2655);
    not g1456(n619 ,n620);
    nor g1457(n12 ,n2491 ,n2427);
    nor g1458(n824 ,n5[7] ,n631);
    nand g1459(n1509 ,n812 ,n1313);
    nand g1460(n1924 ,n1146 ,n1674);
    xnor g1461(n2303 ,n2768 ,n4[59]);
    nand g1462(n1542 ,n2[81] ,n1253);
    or g1463(n1346 ,n2[86] ,n1261);
    nor g1464(n42 ,n2468 ,n2404);
    or g1465(n696 ,n2[55] ,n642);
    nand g1466(n395 ,n2327 ,n275);
    or g1467(n835 ,n2313 ,n629);
    nor g1468(n452 ,n1 ,n315);
    nand g1469(n1179 ,n2[5] ,n657);
    nand g1470(n2154 ,n2042 ,n3[30]);
    nand g1471(n880 ,n4[57] ,n564);
    xnor g1472(n2344 ,n107 ,n206);
    nor g1473(n190 ,n62 ,n189);
    dff g1474(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1904), .Q(n3[39]));
    or g1475(n519 ,n3[47] ,n464);
    nand g1476(n1759 ,n1569 ,n1055);
    nor g1477(n1791 ,n855 ,n1724);
    nand g1478(n1261 ,n7[23] ,n908);
    nand g1479(n1175 ,n2[11] ,n557);
    nand g1480(n998 ,n401 ,n582);
    nand g1481(n2143 ,n7[15] ,n2042);
    nand g1482(n1110 ,n2[47] ,n560);
    nand g1483(n855 ,n429 ,n590);
    or g1484(n1390 ,n2[106] ,n1263);
    nor g1485(n2768 ,n2767 ,n2764);
    nand g1486(n1299 ,n5[16] ,n916);
    nand g1487(n2446 ,n2143 ,n2163);
    xnor g1488(n2367 ,n99 ,n252);
    or g1489(n708 ,n2[50] ,n642);
    nand g1490(n1336 ,n5[1] ,n910);
    nand g1491(n424 ,n2245 ,n311);
    nand g1492(n2595 ,n2532 ,n2594);
    nand g1493(n72 ,n2436 ,n2372);
    nand g1494(n1494 ,n789 ,n1300);
    nand g1495(n2051 ,n2[102] ,n6[1]);
    nor g1496(n1692 ,n956 ,n1454);
    nand g1497(n1881 ,n1093 ,n1624);
    nand g1498(n2062 ,n2[19] ,n6[1]);
    nand g1499(n1034 ,n413 ,n598);
    xnor g1500(n90 ,n2437 ,n2373);
    xnor g1501(n2253 ,n2587 ,n4[9]);
    xnor g1502(n93 ,n2496 ,n2432);
    nand g1503(n1002 ,n4[60] ,n564);
    or g1504(n474 ,n3[44] ,n464);
    not g1505(n2731 ,n2730);
    or g1506(n1353 ,n2[79] ,n1262);
    or g1507(n2750 ,n2565 ,n2747);
    or g1508(n740 ,n2[38] ,n643);
    nand g1509(n2692 ,n4[40] ,n2690);
    nand g1510(n633 ,n7[15] ,n471);
    nand g1511(n645 ,n7[63] ,n450);
    nand g1512(n898 ,n338 ,n488);
    or g1513(n1352 ,n2[80] ,n1261);
    or g1514(n448 ,n310 ,n379);
    nand g1515(n2482 ,n2138 ,n2119);
    nor g1516(n1634 ,n945 ,n1445);
    nand g1517(n2386 ,n2169 ,n2084);
    nand g1518(n1487 ,n767 ,n1290);
    nor g1519(n164 ,n60 ,n163);
    or g1520(n771 ,n2347 ,n627);
    nand g1521(n1003 ,n420 ,n569);
    nand g1522(n2477 ,n2138 ,n2107);
    nor g1523(n831 ,n2312 ,n629);
    xnor g1524(n81 ,n2462 ,n2398);
    nand g1525(n412 ,n2262 ,n273);
    nand g1526(n2480 ,n2138 ,n2114);
    nand g1527(n1857 ,n1067 ,n1602);
    nor g1528(n200 ,n42 ,n199);
    or g1529(n768 ,n2[26] ,n637);
    dff g1530(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1994), .Q(n4[43]));
    xnor g1531(n2358 ,n108 ,n234);
    nand g1532(n1177 ,n2316 ,n649);
    xnor g1533(n2366 ,n121 ,n250);
    or g1534(n2795 ,n9[1] ,n1);
    nand g1535(n1927 ,n1150 ,n1678);
    nor g1536(n1602 ,n754 ,n1412);
    or g1537(n665 ,n2318 ,n624);
    nand g1538(n2237 ,n2042 ,n3[51]);
    nand g1539(n333 ,n2273 ,n312);
    or g1540(n915 ,n453 ,n620);
    nand g1541(n1988 ,n1383 ,n1831);
    nor g1542(n1707 ,n947 ,n1516);
    nand g1543(n2114 ,n2[108] ,n6[1]);
    nand g1544(n1520 ,n664 ,n1205);
    nand g1545(n1482 ,n760 ,n1284);
    nand g1546(n372 ,n2338 ,n312);
    nand g1547(n373 ,n2346 ,n312);
    or g1548(n2776 ,n2559 ,n2775);
    nand g1549(n1297 ,n3[22] ,n909);
    or g1550(n603 ,n4[56] ,n463);
    dff g1551(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1718), .Q(n5[1]));
    nand g1552(n1057 ,n383 ,n581);
    nand g1553(n1006 ,n405 ,n607);
    nand g1554(n1156 ,n2317 ,n649);
    nand g1555(n1421 ,n662 ,n1208);
    nor g1556(n2800 ,n2784 ,n1);
    dff g1557(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1940), .Q(n5[14]));
    nand g1558(n2552 ,n4[52] ,n4[51]);
    not g1559(n2521 ,n4[10]);
    xnor g1560(n88 ,n2471 ,n2407);
    nand g1561(n1485 ,n766 ,n1289);
    nand g1562(n1765 ,n1574 ,n934);
    nand g1563(n1095 ,n2346 ,n653);
    nand g1564(n1282 ,n3[31] ,n917);
    nor g1565(n1705 ,n968 ,n1515);
    not g1566(n378 ,n379);
    or g1567(n2791 ,n9[12] ,n1);
    nand g1568(n1996 ,n1391 ,n1839);
    or g1569(n668 ,n2[63] ,n630);
    dff g1570(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1960), .Q(n3[3]));
    xnor g1571(n2355 ,n80 ,n228);
    nor g1572(n50 ,n2456 ,n2392);
    dff g1573(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1980), .Q(n4[57]));
    nand g1574(n885 ,n4[11] ,n558);
    or g1575(n300 ,n294 ,n299);
    nor g1576(n2576 ,n4[6] ,n2575);
    nand g1577(n1147 ,n2328 ,n650);
    nand g1578(n1787 ,n1595 ,n901);
    nor g1579(n1662 ,n973 ,n1474);
    buf g1580(n6[1] ,n2039);
    nand g1581(n2436 ,n2140 ,n2165);
    nand g1582(n2405 ,n2183 ,n2178);
    nand g1583(n1885 ,n1105 ,n1635);
    nand g1584(n2445 ,n2143 ,n2081);
    nand g1585(n2224 ,n2043 ,n3[37]);
    nor g1586(n458 ,n7[31] ,n378);
    nand g1587(n1780 ,n1589 ,n972);
    nand g1588(n1309 ,n3[15] ,n915);
    nor g1589(n2617 ,n2513 ,n2614);
    xnor g1590(n2505 ,n8[2] ,n263);
    nor g1591(n260 ,n47 ,n259);
    nand g1592(n356 ,n2351 ,n274);
    nand g1593(n868 ,n4[18] ,n565);
    nand g1594(n470 ,n7[55] ,n379);
    not g1595(n298 ,n297);
    xnor g1596(n2317 ,n109 ,n152);
    dff g1597(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1879), .Q(n5[40]));
    nand g1598(n1325 ,n828 ,n1183);
    nor g1599(n826 ,n5[59] ,n645);
    nand g1600(n2624 ,n2621 ,n2620);
    not g1601(n2779 ,n9[6]);
    nand g1602(n1905 ,n1127 ,n1655);
    or g1603(n748 ,n2333 ,n625);
    or g1604(n497 ,n3[51] ,n470);
    xnor g1605(n127 ,n2489 ,n2425);
    dff g1606(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1915), .Q(n3[31]));
    nand g1607(n1123 ,n2[40] ,n560);
    nand g1608(n2471 ,n2139 ,n2092);
    dff g1609(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n292), .Q(n8[1]));
    nor g1610(n2569 ,n4[2] ,n2568);
    nand g1611(n2055 ,n2042 ,n3[17]);
    not g1612(n2544 ,n2543);
    nor g1613(n248 ,n65 ,n247);
    nand g1614(n1050 ,n4[34] ,n656);
    nor g1615(n456 ,n7[55] ,n378);
    nand g1616(n873 ,n4[16] ,n565);
    nand g1617(n965 ,n386 ,n527);
    dff g1618(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1973), .Q(n3[53]));
    or g1619(n477 ,n4[13] ,n467);
    xnor g1620(n2297 ,n2750 ,n4[53]);
    nor g1621(n197 ,n82 ,n196);
    nor g1622(n2661 ,n2556 ,n2660);
    xnor g1623(n131 ,n2457 ,n2393);
    nor g1624(n161 ,n117 ,n160);
    nand g1625(n2460 ,n2141 ,n2083);
    nand g1626(n2182 ,n2043 ,n3[2]);
    nand g1627(n1508 ,n811 ,n1312);
    nand g1628(n1889 ,n1108 ,n1639);
    nand g1629(n351 ,n2371 ,n275);
    xnor g1630(n2325 ,n123 ,n168);
    nor g1631(n455 ,n7[39] ,n378);
    xnor g1632(n99 ,n2495 ,n2431);
    nor g1633(n2650 ,n2519 ,n2647);
    nand g1634(n1181 ,n2[2] ,n657);
    nand g1635(n958 ,n355 ,n474);
    nand g1636(n2236 ,n2[104] ,n6[1]);
    nand g1637(n1588 ,n2[98] ,n1256);
    or g1638(n2639 ,n2635 ,n2637);
    not g1639(n2043 ,n2041);
    dff g1640(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2012), .Q(n4[1]));
    nor g1641(n1789 ,n852 ,n1740);
    nand g1642(n1526 ,n829 ,n1326);
    nor g1643(n2760 ,n2555 ,n2757);
    not g1644(n2780 ,n9[15]);
    nand g1645(n2230 ,n2[66] ,n6[1]);
    nor g1646(n1699 ,n1006 ,n1510);
    xnor g1647(n123 ,n2453 ,n2389);
    nand g1648(n1313 ,n3[12] ,n915);
    nand g1649(n1407 ,n822 ,n1324);
    nand g1650(n2019 ,n1360 ,n1808);
    nand g1651(n1435 ,n771 ,n1223);
    nand g1652(n1335 ,n5[62] ,n914);
    nand g1653(n1099 ,n2345 ,n653);
    dff g1654(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2002), .Q(n4[35]));
    or g1655(n1597 ,n1191 ,n1531);
    nand g1656(n2178 ,n2[33] ,n6[1]);
    nor g1657(n1832 ,n931 ,n1765);
    dff g1658(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1942), .Q(n5[13]));
    nand g1659(n2600 ,n4[15] ,n2597);
    nand g1660(n1497 ,n792 ,n1301);
    nand g1661(n926 ,n4[0] ,n563);
    nor g1662(n761 ,n5[22] ,n636);
    not g1663(n2522 ,n4[20]);
    nor g1664(n2506 ,n264 ,n262);
    nor g1665(n156 ,n28 ,n155);
    nand g1666(n1536 ,n2[87] ,n1253);
    nor g1667(n1646 ,n721 ,n1453);
    nand g1668(n1131 ,n2[35] ,n559);
    nor g1669(n1712 ,n833 ,n1521);
    nor g1670(n158 ,n63 ,n157);
    nor g1671(n1625 ,n939 ,n1434);
    nand g1672(n2072 ,n2042 ,n3[42]);
    nand g1673(n1143 ,n2[28] ,n556);
    nand g1674(n2747 ,n2740 ,n2737);
    or g1675(n543 ,n3[28] ,n466);
    nand g1676(n1267 ,n5[28] ,n919);
    or g1677(n2794 ,n9[16] ,n1);
    nand g1678(n267 ,n8[3] ,n266);
    nor g1679(n1258 ,n7[55] ,n907);
    or g1680(n683 ,n2[61] ,n630);
    dff g1681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1987), .Q(n4[50]));
    xnor g1682(n121 ,n2494 ,n2430);
    nor g1683(n2817 ,n2815 ,n2814);
    nand g1684(n1154 ,n2325 ,n650);
    or g1685(n558 ,n453 ,n380);
    nand g1686(n1737 ,n1547 ,n882);
    not g1687(n2518 ,n7[23]);
    nand g1688(n2383 ,n2226 ,n2225);
    or g1689(n549 ,n3[24] ,n466);
    nand g1690(n1063 ,n2366 ,n655);
    or g1691(n832 ,n2[60] ,n630);
    nand g1692(n1206 ,n5[5] ,n910);
    or g1693(n922 ,n452 ,n606);
    nor g1694(n560 ,n7[47] ,n472);
    nand g1695(n2120 ,n2[26] ,n6[1]);
    nand g1696(n1470 ,n745 ,n1273);
    nand g1697(n1278 ,n3[33] ,n918);
    nand g1698(n1776 ,n1585 ,n1044);
    not g1699(n2524 ,n4[49]);
    nand g1700(n1139 ,n2[30] ,n556);
    nor g1701(n2608 ,n7[23] ,n2606);
    not g1702(n2511 ,n4[34]);
    dff g1703(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n286), .Q(n8[4]));
    nand g1704(n897 ,n4[5] ,n563);
    nand g1705(n2682 ,n2548 ,n2681);
    dff g1706(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1968), .Q(n5[61]));
    nand g1707(n2090 ,n2042 ,n3[22]);
    nand g1708(n2063 ,n2[93] ,n6[1]);
    nor g1709(n269 ,n8[5] ,n268);
    or g1710(n2638 ,n4[25] ,n2636);
    nand g1711(n1878 ,n1092 ,n1625);
    nand g1712(n1762 ,n1572 ,n966);
    nand g1713(n948 ,n349 ,n512);
    nor g1714(n840 ,n2311 ,n629);
    xnor g1715(n2263 ,n2619 ,n4[19]);
    nand g1716(n2200 ,n2[57] ,n6[1]);
    nand g1717(n2084 ,n2[14] ,n6[1]);
    nand g1718(n355 ,n2352 ,n312);
    nand g1719(n861 ,n4[21] ,n565);
    nor g1720(n2628 ,n4[22] ,n2625);
    nand g1721(n2654 ,n4[29] ,n2650);
    xnor g1722(n2245 ,n4[1] ,n2549);
    or g1723(n479 ,n3[26] ,n466);
    nand g1724(n1947 ,n1175 ,n1699);
    nand g1725(n2375 ,n2186 ,n2184);
    nor g1726(n20 ,n2470 ,n2406);
    nand g1727(n2162 ,n2042 ,n3[31]);
    or g1728(n1404 ,n2[94] ,n1260);
    nand g1729(n2010 ,n1372 ,n1817);
    nand g1730(n1432 ,n688 ,n1221);
    nor g1731(n206 ,n49 ,n205);
    nand g1732(n1001 ,n353 ,n578);
    nand g1733(n992 ,n396 ,n614);
    not g1734(n308 ,n307);
    nand g1735(n2241 ,n2[29] ,n6[1]);
    nand g1736(n1427 ,n739 ,n1216);
    nor g1737(n2601 ,n2554 ,n2600);
    nand g1738(n1007 ,n439 ,n506);
    nand g1739(n2218 ,n2[9] ,n6[1]);
    nand g1740(n637 ,n7[31] ,n471);
    or g1741(n681 ,n2350 ,n622);
    nor g1742(n144 ,n69 ,n143);
    or g1743(n686 ,n2315 ,n629);
    or g1744(n618 ,n3[8] ,n467);
    nand g1745(n360 ,n2331 ,n311);
    nand g1746(n903 ,n4[2] ,n563);
    or g1747(n736 ,n2[40] ,n640);
    nand g1748(n1518 ,n827 ,n1224);
    nand g1749(n1760 ,n1570 ,n1020);
    nand g1750(n1503 ,n802 ,n1307);
    nand g1751(n1174 ,n2311 ,n648);
    nand g1752(n889 ,n4[9] ,n558);
    or g1753(n919 ,n452 ,n534);
    or g1754(n489 ,n3[63] ,n463);
    nor g1755(n239 ,n122 ,n238);
    nor g1756(n1822 ,n1011 ,n1755);
    or g1757(n790 ,n2361 ,n626);
    or g1758(n916 ,n452 ,n550);
    nand g1759(n945 ,n332 ,n497);
    or g1760(n1386 ,n2[110] ,n1263);
    dff g1761(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1964), .Q(n3[1]));
    nand g1762(n432 ,n2350 ,n311);
    xnor g1763(n2320 ,n114 ,n158);
    nand g1764(n1043 ,n4[1] ,n563);
    or g1765(n602 ,n4[24] ,n466);
    nand g1766(n1767 ,n1576 ,n870);
    nand g1767(n1039 ,n444 ,n576);
    nor g1768(n819 ,n5[10] ,n621);
    nor g1769(n841 ,n5[56] ,n645);
    or g1770(n911 ,n454 ,n620);
    nand g1771(n2076 ,n2[21] ,n6[1]);
    not g1772(n2597 ,n2596);
    nand g1773(n2047 ,n2[98] ,n6[1]);
    or g1774(n909 ,n459 ,n620);
    nor g1775(n153 ,n109 ,n152);
    or g1776(n793 ,n2[19] ,n634);
    nand g1777(n1072 ,n2359 ,n654);
    nand g1778(n1495 ,n785 ,n1298);
    nand g1779(n902 ,n363 ,n492);
    nor g1780(n243 ,n84 ,n242);
    or g1781(n569 ,n3[12] ,n467);
    nand g1782(n2429 ,n2217 ,n2200);
    nand g1783(n2574 ,n4[4] ,n2573);
    nand g1784(n1033 ,n425 ,n575);
    nand g1785(n1557 ,n2[66] ,n1255);
    nor g1786(n290 ,n278 ,n1);
    nand g1787(n335 ,n2314 ,n274);
    nand g1788(n2448 ,n2143 ,n2157);
    nand g1789(n1979 ,n1343 ,n1822);
    nand g1790(n2657 ,n4[30] ,n2655);
    nor g1791(n702 ,n5[36] ,n641);
    nor g1792(n1673 ,n980 ,n1485);
    nor g1793(n1612 ,n674 ,n1422);
    not g1794(n2538 ,n2537);
    nor g1795(n33 ,n2449 ,n2385);
    nor g1796(n1631 ,n943 ,n1442);
    nand g1797(n2172 ,n2[124] ,n6[1]);
    nor g1798(n561 ,n7[55] ,n472);
    or g1799(n1388 ,n2[90] ,n1260);
    dff g1800(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2022), .Q(n4[11]));
    nand g1801(n1227 ,n3[55] ,n923);
    or g1802(n483 ,n4[59] ,n463);
    nand g1803(n1985 ,n1371 ,n1828);
    nand g1804(n1993 ,n1381 ,n1884);
    nor g1805(n1698 ,n1003 ,n1509);
    nor g1806(n2585 ,n2516 ,n2582);
    nand g1807(n1521 ,n842 ,n1322);
    nand g1808(n1732 ,n1542 ,n1008);
    nand g1809(n2193 ,n2043 ,n3[49]);
    dff g1810(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1996), .Q(n4[41]));
    nand g1811(n631 ,n7[7] ,n450);
    nand g1812(n1168 ,n2320 ,n649);
    nand g1813(n1076 ,n2356 ,n654);
    dff g1814(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1853), .Q(n5[59]));
    nand g1815(n1994 ,n1389 ,n1837);
    nand g1816(n1543 ,n2[80] ,n1253);
    nand g1817(n1120 ,n2[41] ,n560);
    nand g1818(n1172 ,n2[10] ,n557);
    nand g1819(n2489 ,n2243 ,n2195);
    nand g1820(n940 ,n365 ,n505);
    nand g1821(n1249 ,n3[41] ,n921);
    nand g1822(n1987 ,n1370 ,n1830);
    nor g1823(n799 ,n5[54] ,n644);
    xnor g1824(n2328 ,n129 ,n174);
    or g1825(n1402 ,n2[96] ,n1251);
    nand g1826(n1739 ,n1549 ,n888);
    dff g1827(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2034), .Q(n4[23]));
    nand g1828(n393 ,n2267 ,n312);
    nand g1829(n438 ,n2295 ,n311);
    nand g1830(n1157 ,n2[20] ,n628);
    nor g1831(n1605 ,n836 ,n1415);
    nand g1832(n641 ,n7[39] ,n450);
    dff g1833(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2014), .Q(n4[3]));
    nand g1834(n2121 ,n2042 ,n3[26]);
    nand g1835(n2187 ,n2043 ,n3[60]);
    not g1836(n2765 ,n2764);
    not g1837(n277 ,n1);
    nand g1838(n1768 ,n1577 ,n1048);
    nand g1839(n1949 ,n1172 ,n1701);
    nand g1840(n995 ,n321 ,n615);
    or g1841(n484 ,n3[58] ,n463);
    nor g1842(n214 ,n37 ,n213);
    nor g1843(n1637 ,n707 ,n1444);
    or g1844(n1378 ,n2[118] ,n1264);
    nor g1845(n69 ,n2440 ,n2376);
    nand g1846(n1119 ,n2[7] ,n657);
    nand g1847(n1493 ,n786 ,n1297);
    dff g1848(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1873), .Q(n3[61]));
    nor g1849(n67 ,n2467 ,n2403);
    nand g1850(n439 ,n2304 ,n273);
    nand g1851(n1291 ,n3[26] ,n917);
    nand g1852(n635 ,n7[47] ,n450);
    nand g1853(n1248 ,n3[42] ,n921);
    or g1854(n1342 ,n2[89] ,n1260);
    nand g1855(n1024 ,n362 ,n594);
    nand g1856(n1283 ,n3[30] ,n917);
    dff g1857(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1781), .Q(n5[4]));
    or g1858(n604 ,n4[44] ,n464);
    nand g1859(n1895 ,n1114 ,n1645);
    nand g1860(n1005 ,n406 ,n573);
    nand g1861(n315 ,n307 ,n276);
    nand g1862(n2028 ,n1351 ,n1799);
    nand g1863(n980 ,n376 ,n546);
    nor g1864(n2568 ,n2527 ,n2549);
    nand g1865(n1096 ,n2[55] ,n561);
    nor g1866(n2711 ,n2515 ,n2707);
    nor g1867(n659 ,n5[51] ,n644);
    nand g1868(n2770 ,n4[59] ,n2767);
    or g1869(n2792 ,n9[17] ,n1);
    or g1870(n1397 ,n2[100] ,n1251);
    dff g1871(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1921), .Q(n3[27]));
    nand g1872(n2169 ,n2042 ,n3[14]);
    nor g1873(n52 ,n2480 ,n2416);
    dff g1874(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2026), .Q(n4[15]));
    nand g1875(n642 ,n7[55] ,n471);
    nor g1876(n830 ,n2308 ,n629);
    not g1877(n2777 ,n9[7]);
    nand g1878(n1977 ,n1364 ,n1820);
    or g1879(n485 ,n3[1] ,n469);
    nor g1880(n289 ,n283 ,n1);
    or g1881(n600 ,n3[2] ,n469);
    or g1882(n755 ,n2[32] ,n643);
    or g1883(n1385 ,n2[111] ,n1263);
    nor g1884(n459 ,n7[23] ,n378);
    nor g1885(n2799 ,n2785 ,n1);
    or g1886(n693 ,n2359 ,n626);
    or g1887(n1343 ,n2[122] ,n1266);
    xnor g1888(n101 ,n2470 ,n2406);
    not g1889(n2042 ,n2041);
    nand g1890(n1431 ,n818 ,n1219);
    nand g1891(n423 ,n2251 ,n311);
    nand g1892(n2472 ,n2139 ,n2096);
    or g1893(n492 ,n4[3] ,n469);
    nand g1894(n1962 ,n1182 ,n1715);
    nor g1895(n44 ,n2454 ,n2390);
    nor g1896(n1653 ,n965 ,n1466);
    nand g1897(n1062 ,n2368 ,n655);
    nand g1898(n1594 ,n2[93] ,n1252);
    dff g1899(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1926), .Q(n5[35]));
    nor g1900(n1641 ,n951 ,n1451);
    nand g1901(n1183 ,n2312 ,n648);
    dff g1902(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1936), .Q(n3[18]));
    nand g1903(n2016 ,n1363 ,n1811);
    or g1904(n2769 ,n4[59] ,n2765);
    nand g1905(n1591 ,n2[95] ,n1252);
    not g1906(n2773 ,n2772);
    nand g1907(n1450 ,n714 ,n1238);
    nor g1908(n2619 ,n2617 ,n2615);
    dff g1909(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1880), .Q(n3[56]));
    nand g1910(n869 ,n412 ,n495);
    nor g1911(n155 ,n111 ,n154);
    nor g1912(n37 ,n2475 ,n2411);
    nor g1913(n230 ,n10 ,n229);
    dff g1914(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2032), .Q(n4[21]));
    xnor g1915(n84 ,n2490 ,n2426);
    nand g1916(n2005 ,n1402 ,n1848);
    or g1917(n507 ,n4[19] ,n468);
    nand g1918(n886 ,n392 ,n583);
    nand g1919(n1185 ,n2310 ,n648);
    dff g1920(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2797), .Q(n9[17]));
    or g1921(n1396 ,n2[101] ,n1251);
    nand g1922(n2022 ,n1357 ,n1805);
    nor g1923(n182 ,n13 ,n181);
    nand g1924(n1876 ,n1089 ,n1622);
    or g1925(n511 ,n3[53] ,n470);
    or g1926(n2658 ,n4[31] ,n2656);
    or g1927(n502 ,n3[30] ,n466);
    nand g1928(n446 ,n2355 ,n275);
    nand g1929(n2034 ,n1345 ,n1793);
    nand g1930(n2563 ,n2556 ,n2538);
    nand g1931(n939 ,n389 ,n504);
    nor g1932(n1253 ,n7[23] ,n907);
    nor g1933(n2543 ,n4[14] ,n4[13]);
    nand g1934(n2033 ,n1346 ,n1794);
    nor g1935(n2648 ,n4[28] ,n2646);
    nand g1936(n988 ,n4[7] ,n563);
    or g1937(n1377 ,n2[119] ,n1264);
    nand g1938(n1882 ,n1096 ,n1627);
    nand g1939(n411 ,n2268 ,n273);
    nor g1940(n255 ,n93 ,n254);
    xnor g1941(n2287 ,n2705 ,n4[43]);
    or g1942(n2679 ,n4[37] ,n2675);
    nand g1943(n1269 ,n3[39] ,n918);
    nor g1944(n2645 ,n2644 ,n2641);
    or g1945(n491 ,n3[45] ,n464);
    nor g1946(n2537 ,n4[32] ,n7[39]);
    nand g1947(n985 ,n360 ,n551);
    nand g1948(n363 ,n2247 ,n311);
    xnor g1949(n2281 ,n2678 ,n4[37]);
    or g1950(n498 ,n4[29] ,n466);
    nor g1951(n59 ,n2462 ,n2398);
    dff g1952(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2813), .Q(n7[55]));
    nand g1953(n1433 ,n687 ,n1220);
    or g1954(n812 ,n2[12] ,n633);
    nor g1955(n807 ,n5[13] ,n621);
    nand g1956(n1587 ,n2[99] ,n1256);
    not g1957(n273 ,n276);
    nand g1958(n1950 ,n1173 ,n1703);
    nand g1959(n2216 ,n2043 ,n3[36]);
    nand g1960(n2175 ,n2[123] ,n6[1]);
    or g1961(n703 ,n2[34] ,n643);
    nor g1962(n1636 ,n949 ,n1448);
    or g1963(n1384 ,n2[112] ,n1264);
    nor g1964(n1675 ,n769 ,n1487);
    nand g1965(n342 ,n2288 ,n312);
    nand g1966(n1771 ,n1580 ,n1021);
    nor g1967(n2694 ,n2691 ,n2693);
    nor g1968(n1818 ,n1004 ,n1751);
    nand g1969(n1049 ,n384 ,n577);
    nand g1970(n440 ,n2318 ,n311);
    nor g1971(n303 ,n2040 ,n301);
    nand g1972(n1952 ,n1156 ,n1702);
    nand g1973(n2017 ,n1362 ,n1810);
    dff g1974(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1978), .Q(n4[59]));
    xnor g1975(n2338 ,n79 ,n194);
    nand g1976(n1271 ,n5[27] ,n919);
    or g1977(n842 ,n2314 ,n629);
    or g1978(n773 ,n2[56] ,n630);
    nand g1979(n371 ,n2297 ,n312);
    nor g1980(n1835 ,n1031 ,n1768);
    nand g1981(n1969 ,n1103 ,n1634);
    nor g1982(n1645 ,n958 ,n1457);
    nand g1983(n2199 ,n2[35] ,n6[1]);
    dff g1984(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2003), .Q(n4[34]));
    nand g1985(n410 ,n2367 ,n311);
    nand g1986(n1334 ,n845 ,n1185);
    dff g1987(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1893), .Q(n5[31]));
    nand g1988(n408 ,n2300 ,n311);
    nor g1989(n223 ,n83 ,n222);
    dff g1990(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1912), .Q(n3[33]));
    nand g1991(n2387 ,n2078 ,n2044);
    nor g1992(n679 ,n5[43] ,n635);
    nor g1993(n774 ,n5[19] ,n636);
    nand g1994(n2192 ,n2[118] ,n6[1]);
    nor g1995(n2738 ,n2736 ,n2733);
    nand g1996(n1563 ,n2[124] ,n1257);
    nand g1997(n887 ,n4[61] ,n564);
    nand g1998(n2011 ,n1369 ,n1816);
    dff g1999(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1899), .Q(n3[41]));
    dff g2000(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2010), .Q(n4[63]));
    dff g2001(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1983), .Q(n4[54]));
    nand g2002(n2577 ,n4[6] ,n2575);
    or g2003(n730 ,n2[42] ,n640);
    nor g2004(n1798 ,n869 ,n1731);
    nand g2005(n2666 ,n4[33] ,n2661);
    nor g2006(n226 ,n25 ,n225);
    or g2007(n541 ,n4[34] ,n465);
    xor g2008(n2258 ,n4[14] ,n2598);
    nand g2009(n864 ,n434 ,n571);
    nand g2010(n1107 ,n2342 ,n653);
    not g2011(n264 ,n263);
    not g2012(n2508 ,n7[39]);
    nor g2013(n1821 ,n1009 ,n1754);
    nand g2014(n2123 ,n2043 ,n3[45]);
    dff g2015(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1719), .Q(n5[2]));
    xor g2016(n2254 ,n2591 ,n4[10]);
    nand g2017(n294 ,n8[4] ,n8[5]);
    nand g2018(n2139 ,n7[39] ,n2042);
    dff g2019(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1859), .Q(n5[53]));
    nand g2020(n1036 ,n323 ,n509);
    nand g2021(n870 ,n4[46] ,n639);
    nand g2022(n1228 ,n3[54] ,n923);
    nand g2023(n2647 ,n4[27] ,n2644);
    nand g2024(n354 ,n2353 ,n275);
    nor g2025(n1720 ,n712 ,n1527);
    nand g2026(n401 ,n2323 ,n274);
    or g2027(n490 ,n4[4] ,n469);
    nand g2028(n1463 ,n783 ,n1317);
    or g2029(n660 ,n2358 ,n626);
    nand g2030(n2494 ,n2242 ,n2152);
    nand g2031(n1736 ,n1546 ,n879);
    xnor g2032(n2322 ,n118 ,n162);
    nor g2033(n833 ,n5[6] ,n631);
    nand g2034(n1236 ,n5[34] ,n922);
    or g2035(n739 ,n2[62] ,n630);
    nand g2036(n1277 ,n3[34] ,n918);
    dff g2037(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1977), .Q(n4[60]));
    nor g2038(n2587 ,n2585 ,n2583);
    nand g2039(n1478 ,n758 ,n1282);
    nand g2040(n2633 ,n7[23] ,n2631);
    nor g2041(n1814 ,n905 ,n1747);
    nand g2042(n1038 ,n334 ,n485);
    nand g2043(n2126 ,n2[80] ,n6[1]);
    nor g2044(n2761 ,n2760 ,n2759);
    nand g2045(n1596 ,n742 ,n1272);
    nand g2046(n2242 ,n7[63] ,n2043);
    nand g2047(n1032 ,n4[44] ,n639);
    dff g2048(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1895), .Q(n3[44]));
    or g2049(n809 ,n2[14] ,n633);
    dff g2050(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1939), .Q(n3[16]));
    nor g2051(n2704 ,n2514 ,n2700);
    or g2052(n815 ,n2[2] ,n632);
    nand g2053(n2094 ,n2042 ,n3[20]);
    nand g2054(n2766 ,n2763 ,n2762);
    nor g2055(n694 ,n5[38] ,n641);
    not g2056(n2687 ,n2686);
    dff g2057(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1979), .Q(n4[58]));
    dff g2058(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2028), .Q(n4[17]));
    nand g2059(n1118 ,n2338 ,n652);
    or g2060(n1344 ,n2[88] ,n1260);
    nand g2061(n1161 ,n2323 ,n649);
    dff g2062(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1962), .Q(n5[5]));
    dff g2063(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1982), .Q(n4[55]));
    xnor g2064(n2504 ,n8[3] ,n265);
    nand g2065(n2144 ,n2[63] ,n6[1]);
    or g2066(n1387 ,n2[109] ,n1263);
    xnor g2067(n100 ,n2440 ,n2376);
    not g2068(n2510 ,n4[38]);
    dff g2069(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1961), .Q(n5[6]));
    nand g2070(n385 ,n2298 ,n274);
    or g2071(n2535 ,n4[61] ,n4[60]);
    or g2072(n2713 ,n4[45] ,n2709);
    dff g2073(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1909), .Q(n3[35]));
    nor g2074(n2590 ,n4[10] ,n2588);
    nand g2075(n1775 ,n1584 ,n1042);
    nor g2076(n287 ,n284 ,n1);
    dff g2077(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2798), .Q(n9[13]));
    nand g2078(n1067 ,n2363 ,n654);
    nand g2079(n265 ,n8[2] ,n264);
    nor g2080(n176 ,n50 ,n175);
    or g2081(n847 ,n2[3] ,n632);
    nand g2082(n2059 ,n2042 ,n3[41]);
    nand g2083(n1890 ,n1112 ,n1646);
    nand g2084(n1476 ,n751 ,n1278);
    nand g2085(n973 ,n367 ,n533);
    nand g2086(n2492 ,n2242 ,n2149);
    nand g2087(n954 ,n391 ,n520);
    nand g2088(n2185 ,n2[49] ,n6[1]);
    nor g2089(n36 ,n2497 ,n2433);
    nand g2090(n1595 ,n2[92] ,n1252);
    nand g2091(n429 ,n2269 ,n273);
    nand g2092(n1502 ,n801 ,n1306);
    nor g2093(n1813 ,n902 ,n1746);
    nand g2094(n1974 ,n1151 ,n1679);
    nand g2095(n1105 ,n2[50] ,n561);
    nor g2096(n734 ,n5[53] ,n644);
    nand g2097(n2087 ,n2[97] ,n6[1]);
    nor g2098(n225 ,n77 ,n224);
    nor g2099(n192 ,n48 ,n191);
    xnor g2100(n2267 ,n4[23] ,n2631);
    dff g2101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1970), .Q(n5[36]));
    dff g2102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1905), .Q(n3[38]));
    nand g2103(n1874 ,n1088 ,n1620);
    xnor g2104(n2285 ,n2698 ,n4[41]);
    not g2105(n2528 ,n4[5]);
    nand g2106(n2566 ,n2546 ,n2530);
    nand g2107(n1870 ,n1082 ,n1614);
    nand g2108(n2485 ,n2243 ,n2127);
    dff g2109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1937), .Q(n3[17]));
    nand g2110(n1972 ,n1099 ,n1630);
    or g2111(n719 ,n2[1] ,n632);
    xnor g2112(n2247 ,n4[3] ,n2570);
    nand g2113(n1472 ,n747 ,n1275);
    nand g2114(n2201 ,n2[6] ,n6[1]);
    or g2115(n759 ,n2[30] ,n637);
    dff g2116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n287), .Q(n8[2]));
    nand g2117(n2088 ,n2042 ,n3[13]);
    nand g2118(n863 ,n4[20] ,n565);
    nand g2119(n1906 ,n1128 ,n1657);
    nand g2120(n430 ,n2349 ,n273);
    nand g2121(n1922 ,n1144 ,n1672);
    nor g2122(n1722 ,n669 ,n1530);
    nand g2123(n929 ,n4[4] ,n563);
    nand g2124(n1858 ,n1068 ,n1603);
    nor g2125(n628 ,n7[23] ,n472);
    nor g2126(n1599 ,n823 ,n1409);
    nand g2127(n1934 ,n1158 ,n1686);
    nand g2128(n1454 ,n723 ,n1243);
    nand g2129(n2437 ,n2140 ,n2228);
    or g2130(n1405 ,n2[93] ,n1260);
    or g2131(n1349 ,n2[83] ,n1261);
    nand g2132(n2596 ,n2566 ,n2594);
    nand g2133(n2009 ,n1406 ,n1852);
    nand g2134(n933 ,n415 ,n501);
    or g2135(n647 ,n458 ,n380);
    nand g2136(n1065 ,n2365 ,n655);
    nor g2137(n1689 ,n996 ,n1500);
    or g2138(n2295 ,n2744 ,n2746);
    nor g2139(n227 ,n75 ,n226);
    nand g2140(n1887 ,n1107 ,n1638);
    or g2141(n767 ,n2328 ,n623);
    dff g2142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1997), .Q(n4[40]));
    nand g2143(n1937 ,n1162 ,n1689);
    nand g2144(n2038 ,n1468 ,n1789);
    nand g2145(n2439 ,n2140 ,n2232);
    nand g2146(n1898 ,n1117 ,n1648);
    nand g2147(n2058 ,n2[18] ,n6[1]);
    nand g2148(n2081 ,n2[73] ,n6[1]);
    nand g2149(n1458 ,n729 ,n1245);
    nand g2150(n1453 ,n846 ,n1240);
    nand g2151(n1080 ,n2353 ,n651);
    or g2152(n2632 ,n4[23] ,n2631);
    xnor g2153(n2370 ,n89 ,n258);
    or g2154(n808 ,n2364 ,n646);
    nand g2155(n2119 ,n2[110] ,n6[1]);
    nor g2156(n1654 ,n780 ,n1465);
    nand g2157(n1899 ,n1120 ,n1650);
    nand g2158(n1203 ,n5[10] ,n913);
    not g2159(n2041 ,n6[2]);
    nor g2160(n1648 ,n961 ,n1460);
    nand g2161(n2464 ,n2141 ,n2077);
    xnor g2162(n2501 ,n8[6] ,n270);
    xnor g2163(n2560 ,n2516 ,n4[13]);
    nor g2164(n1626 ,n940 ,n1436);
    nand g2165(n2130 ,n2042 ,n3[40]);
    nand g2166(n1761 ,n1571 ,n1023);
    nor g2167(n1681 ,n791 ,n1496);
    xnor g2168(n78 ,n2463 ,n2399);
    or g2169(n710 ,n2[49] ,n642);
    nand g2170(n2118 ,n2[41] ,n6[1]);
    nor g2171(n1709 ,n824 ,n1519);
    nand g2172(n1728 ,n1538 ,n861);
    nand g2173(n2111 ,n2[84] ,n6[1]);
    nand g2174(n331 ,n2291 ,n274);
    nand g2175(n1155 ,n2[21] ,n628);
    dff g2176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1986), .Q(n4[51]));
    or g2177(n816 ,n2[11] ,n633);
    nand g2178(n1900 ,n1122 ,n1651);
    or g2179(n1350 ,n2[82] ,n1261);
    nand g2180(n2453 ,n2142 ,n2053);
    not g2181(n2520 ,n4[22]);
    nand g2182(n621 ,n7[15] ,n450);
    nand g2183(n2422 ,n2219 ,n2208);
    or g2184(n539 ,n4[61] ,n463);
    nand g2185(n1585 ,n2[101] ,n1256);
    nand g2186(n2490 ,n2243 ,n2192);
    nor g2187(n1600 ,n671 ,n1410);
    xnor g2188(n135 ,n2442 ,n2378);
    nor g2189(n1826 ,n1018 ,n1759);
    nand g2190(n963 ,n438 ,n592);
    nand g2191(n2659 ,n7[31] ,n2657);
    or g2192(n567 ,n4[57] ,n463);
    or g2193(n505 ,n3[56] ,n463);
    nand g2194(n2073 ,n2[90] ,n6[1]);
    or g2195(n2762 ,n4[57] ,n2758);
    nand g2196(n1135 ,n2332 ,n652);
    xnor g2197(n2368 ,n93 ,n254);
    or g2198(n499 ,n3[61] ,n463);
    dff g2199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1906), .Q(n3[37]));
    or g2200(n1393 ,n2[103] ,n1251);
    xor g2201(n2286 ,n2703 ,n4[42]);
    nor g2202(n756 ,n5[24] ,n638);
    xor g2203(n2260 ,n2611 ,n7[23]);
    nand g2204(n2222 ,n2[10] ,n6[1]);
    dff g2205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1878), .Q(n3[57]));
    dff g2206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2009), .Q(n4[28]));
    nand g2207(n867 ,n419 ,n507);
    nor g2208(n1834 ,n1029 ,n1767);
    nand g2209(n1504 ,n805 ,n1309);
    nand g2210(n1014 ,n4[56] ,n564);
    not g2211(n2517 ,n4[60]);
    nand g2212(n2415 ,n2091 ,n2086);
    nand g2213(n466 ,n7[31] ,n379);
    nand g2214(n361 ,n2345 ,n274);
    dff g2215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1916), .Q(n3[30]));
    nand g2216(n2450 ,n2143 ,n2122);
    not g2217(n2609 ,n2608);
    nand g2218(n1015 ,n408 ,n603);
    nand g2219(n1567 ,n2[120] ,n1257);
    or g2220(n611 ,n4[12] ,n467);
    nand g2221(n2470 ,n2139 ,n2047);
    nand g2222(n1434 ,n691 ,n1222);
    nor g2223(n211 ,n115 ,n210);
    nor g2224(n204 ,n20 ,n203);
    nand g2225(n2210 ,n2[112] ,n6[1]);
    not g2226(n2573 ,n2572);
    nand g2227(n1501 ,n796 ,n1304);
    nand g2228(n2673 ,n4[35] ,n2670);
    nor g2229(n781 ,n5[18] ,n636);
    nor g2230(n1652 ,n964 ,n1464);
    nand g2231(n467 ,n7[15] ,n379);
    nand g2232(n1556 ,n2[67] ,n1255);
    nand g2233(n2643 ,n2640 ,n2638);
    nand g2234(n2562 ,n2554 ,n2544);
    not g2235(n2516 ,n7[15]);
    or g2236(n554 ,n4[9] ,n467);
    nor g2237(n1622 ,n935 ,n1431);
    nor g2238(n2742 ,n4[53] ,n2739);
    or g2239(n587 ,n4[48] ,n470);
    nor g2240(n2748 ,n2745 ,n2742);
    xor g2241(n2310 ,n95 ,n138);
    or g2242(n616 ,n3[19] ,n468);
    nand g2243(n1481 ,n762 ,n1285);
    or g2244(n2699 ,n4[41] ,n2695);
    nand g2245(n1955 ,n1097 ,n1707);
    nand g2246(n1290 ,n5[20] ,n916);
    nor g2247(n2536 ,n4[52] ,n4[51]);
    xor g2248(n2244 ,n7[7] ,n4[0]);
    nand g2249(n1284 ,n5[22] ,n916);
    nand g2250(n2740 ,n4[51] ,n2735);
    nor g2251(n803 ,n5[14] ,n621);
    nor g2252(n1810 ,n896 ,n1743);
    nor g2253(n171 ,n126 ,n170);
    nand g2254(n1439 ,n698 ,n1229);
    nand g2255(n2021 ,n1358 ,n1806);
    dff g2256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n291), .Q(n8[0]));
    nor g2257(n1667 ,n851 ,n1479);
    nand g2258(n1855 ,n1065 ,n1600);
    or g2259(n605 ,n3[59] ,n463);
    nor g2260(n1684 ,n990 ,n1497);
    nand g2261(n1409 ,n817 ,n1193);
    nand g2262(n1938 ,n1161 ,n1687);
    nor g2263(n1840 ,n1039 ,n1773);
    nand g2264(n1727 ,n1537 ,n860);
    or g2265(n473 ,n4[16] ,n468);
    nor g2266(n1715 ,n837 ,n1524);
    nor g2267(n1257 ,n7[63] ,n907);
    nand g2268(n2394 ,n2090 ,n2089);
    nand g2269(n369 ,n2257 ,n311);
    nand g2270(n2190 ,n2043 ,n3[4]);
    nand g2271(n2135 ,n2042 ,n3[28]);
    or g2272(n2613 ,n4[17] ,n2609);
    nand g2273(n2772 ,n2533 ,n2771);
    nand g2274(n1169 ,n2[13] ,n557);
    nand g2275(n1121 ,n2[4] ,n657);
    nand g2276(n370 ,n2315 ,n275);
    or g2277(n480 ,n4[17] ,n468);
    nand g2278(n2109 ,n2[106] ,n6[1]);
    nand g2279(n2376 ,n2190 ,n2189);
    nor g2280(n1620 ,n933 ,n1430);
    nand g2281(n1240 ,n5[32] ,n922);
    nand g2282(n1443 ,n701 ,n1232);
    nand g2283(n1991 ,n1386 ,n1834);
    nand g2284(n425 ,n2311 ,n275);
    nand g2285(n957 ,n407 ,n599);
    nor g2286(n1679 ,n781 ,n1491);
    nand g2287(n2688 ,n2550 ,n2684);
    xnor g2288(n2323 ,n120 ,n164);
    nand g2289(n1128 ,n2[37] ,n559);
    nand g2290(n1320 ,n5[7] ,n910);
    dff g2291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1984), .Q(n4[53]));
    nand g2292(n877 ,n4[14] ,n558);
    nor g2293(n245 ,n132 ,n244);
    nor g2294(n2604 ,n2516 ,n2601);
    nand g2295(n1511 ,n665 ,n1203);
    nand g2296(n1221 ,n3[58] ,n924);
    nor g2297(n1624 ,n692 ,n1435);
    nor g2298(n2797 ,n2782 ,n1);
    dff g2299(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1934), .Q(n3[19]));
    nor g2300(n1793 ,n859 ,n1726);
    xor g2301(n2262 ,n2618 ,n4[18]);
    dff g2302(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1888), .Q(n5[33]));
    nand g2303(n2197 ,n2[70] ,n6[1]);
    nand g2304(n2194 ,n2043 ,n3[46]);
    nand g2305(n2117 ,n2043 ,n3[59]);
    nand g2306(n1856 ,n1066 ,n1601);
    dff g2307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2808), .Q(n7[15]));
    nand g2308(n1223 ,n5[39] ,n922);
    nor g2309(n2598 ,n2560 ,n2596);
    or g2310(n599 ,n4[42] ,n464);
    nor g2311(n46 ,n2455 ,n2391);
    or g2312(n687 ,n2348 ,n622);
    or g2313(n805 ,n2[15] ,n633);
    nand g2314(n1547 ,n2[76] ,n1254);
    dff g2315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2006), .Q(n4[31]));
    nand g2316(n1729 ,n1539 ,n863);
    or g2317(n2530 ,n4[12] ,n4[11]);
    nand g2318(n436 ,n2278 ,n273);
    nand g2319(n999 ,n403 ,n610);
    nor g2320(n1802 ,n878 ,n1735);
    nand g2321(n1275 ,n3[35] ,n918);
    nand g2322(n2048 ,n2[79] ,n6[1]);
    nand g2323(n1479 ,n757 ,n1281);
    or g2324(n592 ,n4[51] ,n470);
    nand g2325(n2158 ,n2[31] ,n6[1]);
    nor g2326(n1672 ,n765 ,n1484);
    or g2327(n598 ,n4[43] ,n464);
    nand g2328(n1442 ,n705 ,n1230);
    nand g2329(n2012 ,n1368 ,n1815);
    nor g2330(n1811 ,n898 ,n1744);
    nand g2331(n1926 ,n1104 ,n1637);
    nand g2332(n1544 ,n2[79] ,n1254);
    nand g2333(n1915 ,n1137 ,n1666);
    nand g2334(n2004 ,n1401 ,n1847);
    nor g2335(n1701 ,n1010 ,n1512);
    nand g2336(n2079 ,n2[95] ,n6[1]);
    nand g2337(n2015 ,n1365 ,n1812);
    nor g2338(n198 ,n67 ,n197);
    nor g2339(n746 ,n5[26] ,n638);
    or g2340(n701 ,n2[52] ,n642);
    or g2341(n585 ,n3[41] ,n464);
    dff g2342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2800), .Q(n9[2]));
    nand g2343(n1774 ,n1583 ,n1040);
    nand g2344(n1091 ,n2348 ,n651);
    nor g2345(n851 ,n5[23] ,n636);
    nand g2346(n946 ,n352 ,n515);
    nand g2347(n2013 ,n1367 ,n1814);
    xnor g2348(n2289 ,n2712 ,n4[45]);
    nand g2349(n1514 ,n800 ,n1318);
    nand g2350(n1010 ,n440 ,n478);
    nand g2351(n2164 ,n2[127] ,n6[1]);
    nand g2352(n2570 ,n4[2] ,n2568);
    or g2353(n753 ,n2332 ,n625);
    nand g2354(n2403 ,n2162 ,n2158);
    nand g2355(n1098 ,n2[54] ,n561);
    or g2356(n572 ,n4[38] ,n465);
    or g2357(n564 ,n457 ,n380);
    nor g2358(n1657 ,n969 ,n1596);
    nand g2359(n944 ,n4[49] ,n658);
    xnor g2360(n2249 ,n4[5] ,n2574);
    nand g2361(n415 ,n2368 ,n311);
    or g2362(n720 ,n2[46] ,n640);
    not g2363(n282 ,n2502);
    xor g2364(n2806 ,n2[3] ,n9[3]);
    nor g2365(n13 ,n2459 ,n2395);
    xnor g2366(n2248 ,n4[4] ,n2572);
    nand g2367(n1489 ,n772 ,n1292);
    nand g2368(n2161 ,n2[126] ,n6[1]);
    xnor g2369(n86 ,n2461 ,n2397);
    nand g2370(n1946 ,n1170 ,n1698);
    nand g2371(n2089 ,n2[22] ,n6[1]);
    nand g2372(n1318 ,n3[8] ,n915);
    nand g2373(n1055 ,n4[54] ,n658);
    nand g2374(n2209 ,n2[27] ,n6[1]);
    nand g2375(n1836 ,n1098 ,n1629);
    dff g2376(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1856), .Q(n5[56]));
    nand g2377(n1469 ,n2[91] ,n1252);
    nand g2378(n971 ,n431 ,n531);
    nand g2379(n1082 ,n2351 ,n651);
    nand g2380(n2440 ,n2140 ,n2213);
    nor g2381(n1638 ,n709 ,n1447);
    nand g2382(n1152 ,n2[23] ,n628);
    nand g2383(n1251 ,n7[39] ,n908);
    dff g2384(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1896), .Q(n3[43]));
    dff g2385(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1886), .Q(n3[49]));
    or g2386(n1367 ,n2[66] ,n1265);
    nor g2387(n53 ,n2457 ,n2393);
    nand g2388(n935 ,n410 ,n605);
    nor g2389(n228 ,n55 ,n227);
    nand g2390(n2129 ,n2[62] ,n6[1]);
    nand g2391(n2401 ,n2148 ,n2241);
    nor g2392(n814 ,n5[9] ,n621);
    nand g2393(n1250 ,n5[29] ,n919);
    nand g2394(n1285 ,n3[29] ,n917);
    nand g2395(n1035 ,n417 ,n600);
    nand g2396(n2052 ,n2043 ,n3[61]);
    nand g2397(n2134 ,n2[28] ,n6[1]);
    dff g2398(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1944), .Q(n3[13]));
    nor g2399(n142 ,n66 ,n141);
    nor g2400(n60 ,n2450 ,n2386);
    dff g2401(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1883), .Q(n5[38]));
    xnor g2402(n80 ,n2483 ,n2419);
    nand g2403(n1226 ,n5[38] ,n922);
    nand g2404(n1540 ,n2[83] ,n1253);
    not g2405(n2512 ,n4[26]);
    nand g2406(n1474 ,n703 ,n1277);
    nand g2407(n2603 ,n2562 ,n2598);
    nand g2408(n1572 ,n2[115] ,n1258);
    or g2409(n2588 ,n4[9] ,n2584);
    nand g2410(n2591 ,n2589 ,n2588);
    nand g2411(n1071 ,n2360 ,n654);
    or g2412(n589 ,n4[49] ,n470);
    nand g2413(n2618 ,n2614 ,n2613);
    nand g2414(n1578 ,n2[108] ,n1259);
    nand g2415(n2095 ,n2042 ,n3[18]);
    nor g2416(n201 ,n96 ,n200);
    nor g2417(n1717 ,n1045 ,n1526);
    nand g2418(n2147 ,n2[119] ,n6[1]);
    xnor g2419(n83 ,n2480 ,n2416);
    not g2420(n2578 ,n2577);
    nand g2421(n893 ,n423 ,n574);
    xnor g2422(n2301 ,n2761 ,n4[57]);
    nand g2423(n2149 ,n2[120] ,n6[1]);
    nand g2424(n1436 ,n773 ,n1225);
    xnor g2425(n89 ,n2498 ,n2434);
    nand g2426(n2061 ,n2[58] ,n6[1]);
    nand g2427(n1916 ,n1139 ,n1668);
    nor g2428(n1828 ,n1024 ,n1761);
    nand g2429(n1466 ,n778 ,n1269);
    dff g2430(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2801), .Q(n9[10]));
    dff g2431(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1869), .Q(n5[42]));
    or g2432(n540 ,n3[31] ,n466);
    xnor g2433(n2311 ,n98 ,n140);
    nand g2434(n422 ,n2301 ,n311);
    nor g2435(n2629 ,n2520 ,n2626);
    or g2436(n520 ,n3[46] ,n464);
    nor g2437(n685 ,n5[41] ,n635);
    nand g2438(n1448 ,n710 ,n1237);
    dff g2439(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1890), .Q(n5[32]));
    or g2440(n924 ,n457 ,n620);
    or g2441(n596 ,n4[54] ,n470);
    nor g2442(n1628 ,n694 ,n1437);
    nand g2443(n2212 ,n2[8] ,n6[1]);
    nand g2444(n1331 ,n5[2] ,n910);
    nand g2445(n1754 ,n1564 ,n994);
    nand g2446(n2006 ,n1403 ,n1849);
    nand g2447(n2007 ,n1404 ,n1850);
    nand g2448(n1763 ,n1573 ,n1053);
    dff g2449(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1959), .Q(n3[4]));
    nor g2450(n2767 ,n2523 ,n2763);
    nand g2451(n1426 ,n681 ,n1214);
    nand g2452(n1326 ,n3[0] ,n911);
    xnor g2453(n2275 ,n2656 ,n4[31]);
    xnor g2454(n94 ,n2476 ,n2412);
    nand g2455(n1537 ,n2[86] ,n1253);
    nand g2456(n394 ,n2333 ,n274);
    or g2457(n496 ,n4[0] ,n469);
    dff g2458(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1910), .Q(n5[25]));
    nor g2459(n1682 ,n987 ,n1493);
    nor g2460(n1801 ,n876 ,n1734);
    nand g2461(n981 ,n445 ,n482);
    xnor g2462(n79 ,n2466 ,n2402);
    nand g2463(n2142 ,n7[23] ,n2042);
    nor g2464(n1819 ,n1017 ,n1752);
    or g2465(n529 ,n3[38] ,n465);
    nand g2466(n270 ,n8[5] ,n268);
    dff g2467(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1992), .Q(n4[45]));
    or g2468(n789 ,n2[21] ,n634);
    or g2469(n525 ,n3[42] ,n464);
    nand g2470(n925 ,n4[47] ,n639);
    nor g2471(n1697 ,n834 ,n1517);
    nand g2472(n1225 ,n3[56] ,n924);
    or g2473(n2788 ,n9[4] ,n1);
    nand g2474(n2397 ,n2113 ,n2110);
    nand g2475(n1097 ,n2[6] ,n657);
    or g2476(n778 ,n2[39] ,n643);
    nand g2477(n983 ,n394 ,n548);
    nor g2478(n1704 ,n1019 ,n1514);
    nand g2479(n1307 ,n3[16] ,n909);
    nand g2480(n2198 ,n2043 ,n3[5]);
    nand g2481(n632 ,n7[7] ,n471);
    nand g2482(n2409 ,n2224 ,n2221);
    nand g2483(n2419 ,n2155 ,n2150);
    nand g2484(n895 ,n4[23] ,n565);
    dff g2485(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2819), .Q(n9[19]));
    nand g2486(n367 ,n2342 ,n275);
    nor g2487(n586 ,n7[47] ,n451);
    nand g2488(n2498 ,n2242 ,n2161);
    nand g2489(n1017 ,n382 ,n539);
    nor g2490(n559 ,n7[39] ,n472);
    xnor g2491(n2340 ,n87 ,n198);
    nor g2492(n1706 ,n821 ,n1463);
    nor g2493(n175 ,n129 ,n174);
    nand g2494(n2377 ,n2198 ,n2196);
    nand g2495(n1220 ,n5[40] ,n912);
    nand g2496(n1986 ,n1382 ,n1829);
    nand g2497(n1473 ,n748 ,n1276);
    or g2498(n601 ,n3[0] ,n469);
    not g2499(n471 ,n472);
    nand g2500(n1782 ,n1590 ,n960);
    dff g2501(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1908), .Q(n3[36]));
    nand g2502(n2131 ,n2[46] ,n6[1]);
    nand g2503(n1747 ,n1557 ,n903);
    nor g2504(n2641 ,n4[26] ,n2638);
    nand g2505(n1414 ,n790 ,n1197);
    nand g2506(n413 ,n2287 ,n311);
    nand g2507(n2469 ,n2139 ,n2087);
    nand g2508(n1321 ,n5[55] ,n920);
    nor g2509(n690 ,n5[40] ,n635);
    nand g2510(n2165 ,n2[64] ,n6[1]);
    xnor g2511(n118 ,n2450 ,n2386);
    not g2512(n461 ,n462);
    or g2513(n1392 ,n2[104] ,n1263);
    nand g2514(n1319 ,n3[11] ,n915);
    xor g2515(n2302 ,n2766 ,n4[58]);
    nand g2516(n1457 ,n725 ,n1244);
    xnor g2517(n124 ,n2444 ,n2380);
    nand g2518(n421 ,n2290 ,n312);
    nand g2519(n1230 ,n3[53] ,n923);
    nor g2520(n2652 ,n2650 ,n2648);
    nor g2521(n652 ,n7[31] ,n462);
    nand g2522(n320 ,n2370 ,n274);
    nor g2523(n66 ,n2439 ,n2375);
    nand g2524(n1045 ,n443 ,n601);
    xor g2525(n2309 ,n90 ,n72);
    nand g2526(n2203 ,n2043 ,n3[35]);
    or g2527(n597 ,n4[55] ,n470);
    dff g2528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1965), .Q(n3[0]));
    or g2529(n733 ,n2337 ,n625);
    nor g2530(n486 ,n7[55] ,n451);
    nand g2531(n2572 ,n4[3] ,n2571);
    dff g2532(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1897), .Q(n5[30]));
    or g2533(n594 ,n4[52] ,n470);
    nand g2534(n297 ,n2040 ,n277);
    nand g2535(n1231 ,n5[36] ,n922);
    nand g2536(n1150 ,n2[24] ,n556);
    nand g2537(n1498 ,n793 ,n1302);
    nand g2538(n2735 ,n4[50] ,n2732);
    or g2539(n917 ,n458 ,n620);
    xnor g2540(n2271 ,n2645 ,n4[27]);
    or g2541(n476 ,n4[28] ,n466);
    or g2542(n658 ,n456 ,n380);
    xnor g2543(n2327 ,n128 ,n172);
    nand g2544(n2204 ,n2[114] ,n6[1]);
    nor g2545(n1702 ,n814 ,n1407);
    nand g2546(n1992 ,n1387 ,n1835);
    nand g2547(n2238 ,n2[69] ,n6[1]);
    nand g2548(n1328 ,n3[3] ,n911);
    nor g2549(n232 ,n16 ,n231);
    nand g2550(n2373 ,n2177 ,n2174);
    nand g2551(n319 ,n2312 ,n273);
    nand g2552(n1910 ,n1132 ,n1661);
    dff g2553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2036), .Q(n4[25]));
    nand g2554(n865 ,n4[58] ,n564);
    or g2555(n680 ,n5[1] ,n631);
    or g2556(n783 ,n2316 ,n624);
    nand g2557(n1068 ,n2362 ,n654);
    nand g2558(n1219 ,n3[59] ,n924);
    xor g2559(n2814 ,n9[7] ,n9[0]);
    nand g2560(n2181 ,n2[2] ,n6[1]);
    or g2561(n794 ,n2324 ,n623);
    nor g2562(n749 ,n5[25] ,n638);
    nand g2563(n1066 ,n2364 ,n655);
    nand g2564(n1559 ,n2[64] ,n1255);
    nor g2565(n62 ,n2463 ,n2399);
    nand g2566(n2229 ,n2[38] ,n6[1]);
    nand g2567(n1306 ,n5[14] ,n913);
    nand g2568(n1911 ,n1133 ,n1662);
    nor g2569(n16 ,n2484 ,n2420);
    nand g2570(n2451 ,n2143 ,n2048);
    xnor g2571(n2319 ,n113 ,n156);
    or g2572(n770 ,n2[25] ,n637);
    or g2573(n1371 ,n2[116] ,n1264);
    nand g2574(n2196 ,n2[5] ,n6[1]);
    xnor g2575(n2298 ,n2748 ,n4[54]);
    xnor g2576(n133 ,n2458 ,n2394);
    dff g2577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2018), .Q(n4[7]));
    dff g2578(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2804), .Q(n9[18]));
    nand g2579(n1197 ,n5[53] ,n920);
    nand g2580(n1201 ,n5[50] ,n920);
    nand g2581(n377 ,n2334 ,n274);
    nor g2582(n24 ,n2444 ,n2380);
    dff g2583(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1924), .Q(n3[26]));
    nand g2584(n1425 ,n668 ,n1213);
    nand g2585(n1571 ,n2[116] ,n1258);
    or g2586(n493 ,n4[47] ,n464);
    nand g2587(n2496 ,n2242 ,n2172);
    nand g2588(n465 ,n7[39] ,n379);
    nand g2589(n960 ,n4[32] ,n656);
    nand g2590(n1298 ,n5[17] ,n916);
    nand g2591(n1142 ,n2330 ,n650);
    dff g2592(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1955), .Q(n3[6]));
    dff g2593(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1881), .Q(n5[39]));
    nor g2594(n804 ,n5[46] ,n635);
    xnor g2595(n2356 ,n105 ,n230);
    nor g2596(n1677 ,n774 ,n1489);
    not g2597(n2753 ,n2752);
    or g2598(n1366 ,n2[67] ,n1265);
    or g2599(n844 ,n2371 ,n646);
    dff g2600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1922), .Q(n5[21]));
    nand g2601(n2611 ,n2606 ,n2607);
    nor g2602(n454 ,n7[7] ,n378);
    not g2603(n2542 ,n2541);
    dff g2604(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1867), .Q(n5[45]));
    nand g2605(n1090 ,n2[58] ,n562);
    nand g2606(n338 ,n2249 ,n312);
    xnor g2607(n2351 ,n134 ,n220);
    dff g2608(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2812), .Q(n7[47]));
    nand g2609(n1507 ,n813 ,n1311);
    or g2610(n548 ,n3[25] ,n466);
    nand g2611(n2067 ,n2[53] ,n6[1]);
    nand g2612(n1913 ,n1136 ,n1665);
    nand g2613(n1332 ,n5[63] ,n914);
    nor g2614(n1792 ,n857 ,n1725);
    nand g2615(n435 ,n2266 ,n273);
    nand g2616(n1723 ,n1533 ,n1046);
    nand g2617(n1555 ,n2[68] ,n1255);
    or g2618(n843 ,n2367 ,n646);
    nor g2619(n2684 ,n4[39] ,n2682);
    nor g2620(n2804 ,n2786 ,n1);
    or g2621(n514 ,n4[62] ,n463);
    nand g2622(n1338 ,n5[11] ,n913);
    xnor g2623(n76 ,n2464 ,n2400);
    dff g2624(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1913), .Q(n3[32]));
    xnor g2625(n97 ,n2485 ,n2421);
    or g2626(n757 ,n2331 ,n623);
    nand g2627(n1735 ,n1545 ,n877);
    nor g2628(n654 ,n7[55] ,n462);
    nand g2629(n1873 ,n1086 ,n1618);
    nor g2630(n1850 ,n1057 ,n1784);
    nor g2631(n1795 ,n862 ,n1728);
    nand g2632(n1146 ,n2[26] ,n556);
    nor g2633(n1656 ,n743 ,n1341);
    nand g2634(n1021 ,n4[42] ,n639);
    nand g2635(n1954 ,n1119 ,n1705);
    nor g2636(n1608 ,n666 ,n1418);
    nor g2637(n620 ,n1 ,n449);
    nor g2638(n207 ,n107 ,n206);
    nand g2639(n1058 ,n4[43] ,n639);
    nor g2640(n674 ,n5[45] ,n635);
    or g2641(n779 ,n2326 ,n623);
    nand g2642(n1983 ,n1378 ,n1826);
    dff g2643(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1860), .Q(n5[52]));
    nor g2644(n285 ,n280 ,n1);
    or g2645(n639 ,n460 ,n380);
    nand g2646(n984 ,n368 ,n549);
    nand g2647(n2202 ,n2043 ,n3[6]);
    nand g2648(n1417 ,n660 ,n1201);
    nand g2649(n1337 ,n5[61] ,n914);
    nand g2650(n1568 ,n2[119] ,n1258);
    nand g2651(n1144 ,n2329 ,n650);
    nor g2652(n258 ,n36 ,n257);
    xnor g2653(n2369 ,n112 ,n256);
    xnor g2654(n2306 ,n2775 ,n4[62]);
    nor g2655(n1808 ,n892 ,n1741);
    nand g2656(n1030 ,n416 ,n572);
    nand g2657(n1446 ,n708 ,n1235);
    nand g2658(n1440 ,n750 ,n1228);
    nor g2659(n2690 ,n2687 ,n2684);
    nand g2660(n1242 ,n3[46] ,n921);
    or g2661(n1375 ,n2[121] ,n1266);
    nand g2662(n1918 ,n1141 ,n1669);
    nand g2663(n1330 ,n5[3] ,n910);
    or g2664(n914 ,n452 ,n526);
    xnor g2665(n2324 ,n102 ,n166);
    xnor g2666(n92 ,n2492 ,n2428);
    nand g2667(n1340 ,n3[18] ,n909);
    nand g2668(n1093 ,n2347 ,n653);
    or g2669(n1391 ,n2[105] ,n1263);
    nand g2670(n882 ,n4[12] ,n558);
    nand g2671(n2547 ,n4[61] ,n7[63]);
    nor g2672(n1671 ,n979 ,n1483);
    xnor g2673(n2314 ,n135 ,n146);
    nor g2674(n1843 ,n1005 ,n1776);
    xnor g2675(n2279 ,n2671 ,n4[35]);
    nand g2676(n2491 ,n2243 ,n2147);
    dff g2677(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1956), .Q(n5[8]));
    or g2678(n731 ,n2338 ,n625);
    nand g2679(n441 ,n2369 ,n273);
    nand g2680(n1872 ,n1084 ,n1616);
    nor g2681(n1693 ,n998 ,n1504);
    xnor g2682(n2257 ,n2596 ,n4[13]);
    nand g2683(n2479 ,n2138 ,n2112);
    nor g2684(n1661 ,n749 ,n1473);
    or g2685(n792 ,n2[20] ,n634);
    dff g2686(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1974), .Q(n5[18]));
    not g2687(n2781 ,n9[11]);
    nand g2688(n427 ,n2270 ,n273);
    or g2689(n723 ,n2[45] ,n640);
    dff g2690(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1862), .Q(n5[50]));
    nand g2691(n2558 ,n2557 ,n2542);
    nand g2692(n1113 ,n2[45] ,n560);
    nand g2693(n1246 ,n5[31] ,n919);
    nand g2694(n1583 ,n2[103] ,n1256);
    nand g2695(n2758 ,n2539 ,n2757);
    nor g2696(n707 ,n5[35] ,n641);
    nand g2697(n1584 ,n2[102] ,n1256);
    nand g2698(n1109 ,n2341 ,n653);
    nand g2699(n317 ,n2325 ,n275);
    nor g2700(n291 ,n8[0] ,n1);
    xnor g2701(n2503 ,n8[4] ,n267);
    nand g2702(n2423 ,n2237 ,n2227);
    nor g2703(n2565 ,n2553 ,n2536);
    not g2704(n284 ,n2505);
    nand g2705(n2391 ,n2065 ,n2062);
    nand g2706(n2589 ,n4[9] ,n2585);
    nand g2707(n2640 ,n4[25] ,n2635);
    nand g2708(n1984 ,n1379 ,n1827);
    nand g2709(n977 ,n372 ,n502);
    nand g2710(n1101 ,n2344 ,n653);
    nand g2711(n1087 ,n2349 ,n651);
    nand g2712(n1935 ,n1159 ,n1681);
    dff g2713(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1925), .Q(n3[25]));
    nor g2714(n1674 ,n982 ,n1486);
    nor g2715(n1800 ,n871 ,n1733);
    nor g2716(n181 ,n136 ,n180);
    nand g2717(n1235 ,n3[50] ,n923);
    nand g2718(n1742 ,n1552 ,n988);
    or g2719(n574 ,n4[7] ,n469);
    nand g2720(n969 ,n361 ,n530);
    nand g2721(n2412 ,n2130 ,n2075);
    nor g2722(n224 ,n52 ,n223);
    nand g2723(n1871 ,n1083 ,n1615);
    nor g2724(n1630 ,n699 ,n1439);
    nor g2725(n29 ,n2473 ,n2409);
    nor g2726(n1688 ,n992 ,n1499);
    nand g2727(n1202 ,n5[49] ,n920);
    nand g2728(n1866 ,n1078 ,n1610);
    xor g2729(n2300 ,n2564 ,n2756);
    nand g2730(n1437 ,n695 ,n1226);
    nand g2731(n1162 ,n2[17] ,n628);
    nand g2732(n390 ,n2276 ,n274);
    nand g2733(n1510 ,n816 ,n1319);
    nor g2734(n1615 ,n928 ,n1425);
    dff g2735(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1981), .Q(n4[56]));
    nand g2736(n1975 ,n1380 ,n1818);
    nand g2737(n937 ,n346 ,n503);
    or g2738(n530 ,n3[37] ,n465);
    nand g2739(n2717 ,n4[46] ,n2715);
    nand g2740(n936 ,n341 ,n484);
    nand g2741(n986 ,n4[35] ,n656);
    nand g2742(n2457 ,n2142 ,n2064);
    or g2743(n704 ,n2[51] ,n642);
    nand g2744(n2155 ,n2042 ,n3[47]);
    nand g2745(n442 ,n2271 ,n312);
    nor g2746(n380 ,n314 ,n312);
    nand g2747(n359 ,n2363 ,n275);
    dff g2748(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2023), .Q(n4[12]));
    xnor g2749(n2259 ,n2603 ,n4[15]);
    nor g2750(n2667 ,n4[34] ,n2664);
    or g2751(n500 ,n4[2] ,n469);
    or g2752(n494 ,n4[1] ,n469);
    xnor g2753(n2348 ,n94 ,n214);
    or g2754(n698 ,n2345 ,n627);
    dff g2755(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1947), .Q(n3[11]));
    nor g2756(n780 ,n5[28] ,n638);
    xnor g2757(n2255 ,n4[11] ,n2593);
    nand g2758(n1279 ,n5[24] ,n919);
    nand g2759(n1070 ,n2318 ,n649);
    nand g2760(n1941 ,n1165 ,n1693);
    nand g2761(n1140 ,n2[8] ,n557);
    or g2762(n784 ,n2336 ,n625);
    nand g2763(n1108 ,n2[48] ,n561);
    nand g2764(n1932 ,n1155 ,n1683);
    nor g2765(n241 ,n127 ,n240);
    nor g2766(n1623 ,n936 ,n1432);
    xnor g2767(n2276 ,n2563 ,n2660);
    not g2768(n2668 ,n2667);
    not g2769(n2525 ,n4[36]);
    nand g2770(n1304 ,n5[15] ,n913);
    nor g2771(n205 ,n88 ,n204);
    nor g2772(n63 ,n2447 ,n2383);
    nand g2773(n1083 ,n2[63] ,n562);
    nand g2774(n1971 ,n1102 ,n1632);
    nor g2775(n17 ,n2451 ,n2387);
    nor g2776(n457 ,n7[63] ,n378);
    nor g2777(n1643 ,n954 ,n1452);
    nor g2778(n1640 ,n716 ,n1449);
    nand g2779(n2177 ,n2043 ,n3[1]);
    nand g2780(n1292 ,n5[19] ,n916);
    nand g2781(n2243 ,n7[55] ,n2042);
    nor g2782(n208 ,n34 ,n207);
    nor g2783(n1651 ,n735 ,n1462);
    nand g2784(n1879 ,n1091 ,n1621);
    nand g2785(n2206 ,n2[7] ,n6[1]);
    nand g2786(n1079 ,n2354 ,n651);
    dff g2787(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1870), .Q(n5[43]));
    nand g2788(n1569 ,n2[118] ,n1258);
    xor g2789(n2280 ,n2676 ,n4[36]);
    nand g2790(n2032 ,n1347 ,n1795);
    or g2791(n787 ,n2[10] ,n633);
    or g2792(n839 ,n5[3] ,n631);
    nor g2793(n21 ,n2441 ,n2377);
    nor g2794(n143 ,n100 ,n142);
    nor g2795(n199 ,n87 ,n198);
    nand g2796(n1459 ,n731 ,n1247);
    or g2797(n1398 ,n2[99] ,n1251);
    nand g2798(n382 ,n2305 ,n312);
    nor g2799(n179 ,n133 ,n178);
    nand g2800(n353 ,n2307 ,n275);
    nand g2801(n403 ,n2322 ,n273);
    nand g2802(n329 ,n2357 ,n275);
    not g2803(n2507 ,n7[47]);
    nand g2804(n1554 ,n2[69] ,n1255);
    nand g2805(n1088 ,n2[60] ,n562);
    nand g2806(n1424 ,n677 ,n1212);
    nand g2807(n1100 ,n2[53] ,n561);
    nor g2808(n1839 ,n1036 ,n1772);
    nand g2809(n1779 ,n1588 ,n1050);
    or g2810(n527 ,n3[39] ,n465);
    or g2811(n715 ,n2341 ,n627);
    nand g2812(n468 ,n7[23] ,n379);
    nand g2813(n463 ,n7[63] ,n379);
    not g2814(n2515 ,n4[44]);
    nand g2815(n2068 ,n2[42] ,n6[1]);
    nand g2816(n2816 ,n2814 ,n2815);
    nand g2817(n1745 ,n1555 ,n929);
    nand g2818(n1023 ,n4[52] ,n658);
    nor g2819(n236 ,n27 ,n235);
    nand g2820(n2283 ,n2689 ,n2688);
    nor g2821(n1610 ,n689 ,n1420);
    xnor g2822(n2359 ,n116 ,n236);
    nand g2823(n2110 ,n2[25] ,n6[1]);
    or g2824(n510 ,n3[54] ,n470);
    nand g2825(n1743 ,n1553 ,n894);
    nand g2826(n947 ,n335 ,n591);
    nor g2827(n149 ,n106 ,n148);
    nor g2828(n1842 ,n1030 ,n1775);
    nand g2829(n2454 ,n2142 ,n2146);
    nand g2830(n2382 ,n2223 ,n2222);
    nand g2831(n1465 ,n784 ,n1267);
    nand g2832(n386 ,n2347 ,n274);
    xnor g2833(n2347 ,n119 ,n212);
    xnor g2834(n114 ,n2448 ,n2384);
    nor g2835(n147 ,n135 ,n146);
    or g2836(n1345 ,n2[87] ,n1261);
    nand g2837(n2054 ,n2042 ,n3[52]);
    nor g2838(n1796 ,n864 ,n1729);
    or g2839(n662 ,n2354 ,n622);
    xnor g2840(n2315 ,n106 ,n148);
    nand g2841(n2466 ,n2141 ,n2074);
    dff g2842(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1894), .Q(n3[45]));
    nand g2843(n1724 ,n1534 ,n854);
    xnor g2844(n132 ,n2491 ,n2427);
    dff g2845(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1854), .Q(n5[58]));
    nand g2846(n2752 ,n2751 ,n2749);
    dff g2847(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1988), .Q(n4[49]));
    nor g2848(n64 ,n2496 ,n2432);
    nor g2849(n834 ,n5[11] ,n621);
    nor g2850(n57 ,n2489 ,n2425);
    nand g2851(n1027 ,n325 ,n528);
    nand g2852(n1533 ,n2[90] ,n1252);
    nor g2853(n229 ,n80 ,n228);
    or g2854(n532 ,n3[7] ,n469);
    or g2855(n1359 ,n2[73] ,n1262);
    nand g2856(n2092 ,n2[99] ,n6[1]);
    not g2857(n280 ,n2504);
    dff g2858(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2031), .Q(n4[20]));
    dff g2859(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1903), .Q(n5[27]));
    nor g2860(n257 ,n112 ,n256);
    nand g2861(n2026 ,n1353 ,n1801);
    dff g2862(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2802), .Q(n9[1]));
    nand g2863(n1429 ,n848 ,n1215);
    nor g2864(n1827 ,n1022 ,n1760);
    nand g2865(n644 ,n7[55] ,n450);
    nand g2866(n1149 ,n2327 ,n650);
    nand g2867(n1042 ,n4[38] ,n656);
    nor g2868(n2612 ,n2610 ,n2608);
    or g2869(n714 ,n2[48] ,n642);
    nand g2870(n2407 ,n2203 ,n2199);
    nor g2871(n788 ,n5[17] ,n636);
    nand g2872(n640 ,n7[47] ,n471);
    or g2873(n848 ,n2349 ,n622);
    nand g2874(n420 ,n2320 ,n273);
    nand g2875(n905 ,n447 ,n500);
    dff g2876(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1917), .Q(n5[23]));
    nand g2877(n1460 ,n730 ,n1248);
    nand g2878(n2137 ,n2[71] ,n6[1]);
    xnor g2879(n2273 ,n2652 ,n4[29]);
    nand g2880(n1749 ,n1559 ,n926);
    or g2881(n578 ,n4[63] ,n463);
    nor g2882(n722 ,n5[62] ,n645);
    nand g2883(n2495 ,n2242 ,n2175);
    nand g2884(n2097 ,n2[23] ,n6[1]);
    or g2885(n593 ,n4[50] ,n470);
    nor g2886(n1714 ,n1038 ,n1525);
    xnor g2887(n2329 ,n131 ,n176);
    nand g2888(n1126 ,n2335 ,n652);
    nand g2889(n1471 ,n744 ,n1274);
    dff g2890(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1976), .Q(n4[61]));
    dff g2891(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2013), .Q(n4[2]));
    nor g2892(n1676 ,n983 ,n1488);
    nand g2893(n1247 ,n5[30] ,n919);
    nand g2894(n1011 ,n402 ,n521);
    nand g2895(n1178 ,n2314 ,n648);
    or g2896(n488 ,n4[5] ,n469);
    nand g2897(n1785 ,n1330 ,n1400);
    or g2898(n1389 ,n2[107] ,n1263);
    nor g2899(n735 ,n5[29] ,n638);
    nand g2900(n1553 ,n2[70] ,n1255);
    nand g2901(n987 ,n388 ,n552);
    or g2902(n750 ,n2[54] ,n642);
    nand g2903(n1757 ,n1567 ,n1014);
    nand g2904(n1998 ,n1393 ,n1841);
    nand g2905(n1196 ,n5[54] ,n920);
    nand g2906(n630 ,n7[63] ,n471);
    nor g2907(n2818 ,n1 ,n2817);
    dff g2908(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1927), .Q(n3[24]));
    or g2909(n705 ,n2[53] ,n642);
    nand g2910(n2232 ,n2[67] ,n6[1]);
    not g2911(n2526 ,n4[21]);
    nor g2912(n220 ,n26 ,n219);
    nor g2913(n23 ,n2485 ,n2421);
    nand g2914(n2221 ,n2[37] ,n6[1]);
    nor g2915(n2802 ,n2778 ,n1);
    nor g2916(n1616 ,n930 ,n1427);
    nand g2917(n2548 ,n4[38] ,n2508);
    nand g2918(n930 ,n320 ,n553);
    nand g2919(n1778 ,n1587 ,n986);
    nand g2920(n2459 ,n2142 ,n2060);
    nand g2921(n263 ,n8[1] ,n8[0]);
    or g2922(n760 ,n2330 ,n623);
    or g2923(n571 ,n4[20] ,n468);
    or g2924(n752 ,n2362 ,n626);
    nand g2925(n1170 ,n2[12] ,n557);
    nand g2926(n1211 ,n5[44] ,n912);
    nand g2927(n1966 ,n1186 ,n1720);
    dff g2928(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2795), .Q(n9[0]));
    nand g2929(n2056 ,n2[83] ,n6[1]);
    nand g2930(n1928 ,n1149 ,n1677);
    nor g2931(n1805 ,n886 ,n1738);
    nor g2932(n2698 ,n2697 ,n2696);
    nand g2933(n368 ,n2332 ,n273);
    nand g2934(n2441 ,n2140 ,n2238);
    nand g2935(n1512 ,n787 ,n1314);
    xnor g2936(n2256 ,n2595 ,n4[12]);
    dff g2937(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1958), .Q(n5[7]));
    nand g2938(n952 ,n336 ,n510);
    nand g2939(n1412 ,n775 ,n1321);
    or g2940(n850 ,n5[60] ,n645);
    or g2941(n588 ,n4[46] ,n464);
    nand g2942(n1020 ,n4[53] ,n658);
    nor g2943(n1607 ,n776 ,n1417);
    xnor g2944(n98 ,n2439 ,n2375);
    nand g2945(n2680 ,n4[37] ,n2677);
    nand g2946(n2075 ,n2[40] ,n6[1]);
    xnor g2947(n2296 ,n2747 ,n4[52]);
    nand g2948(n366 ,n2277 ,n275);
    dff g2949(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1957), .Q(n3[5]));
    not g2950(n2649 ,n2648);
    nand g2951(n2444 ,n2143 ,n2180);
    dff g2952(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1995), .Q(n4[42]));
    xnor g2953(n113 ,n2447 ,n2383);
    or g2954(n777 ,n2[24] ,n637);
    nand g2955(n1523 ,n815 ,n1315);
    nand g2956(n1576 ,n2[110] ,n1259);
    nand g2957(n2700 ,n4[41] ,n2697);
    dff g2958(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1901), .Q(n3[40]));
    or g2959(n2749 ,n4[54] ,n2743);
    nand g2960(n1411 ,n808 ,n1195);
    nand g2961(n1480 ,n759 ,n1283);
    nand g2962(n2151 ,n2[121] ,n6[1]);
    dff g2963(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2809), .Q(n7[7]));
    nor g2964(n1614 ,n679 ,n1424);
    nor g2965(n1696 ,n1000 ,n1508);
    or g2966(n732 ,n2[41] ,n640);
    nor g2967(n653 ,n7[39] ,n462);
    xnor g2968(n82 ,n2467 ,n2403);
    xnor g2969(n104 ,n2493 ,n2429);
    not g2970(n450 ,n451);
    dff g2971(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2796), .Q(n9[6]));
    nand g2972(n2720 ,n7[47] ,n2717);
    nand g2973(n324 ,n2299 ,n273);
    not g2974(n2616 ,n2615);
    nor g2975(n2774 ,n2534 ,n2772);
    dff g2976(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n288), .Q(n8[5]));
    nand g2977(n927 ,n409 ,n496);
    dff g2978(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1882), .Q(n3[55]));
    nand g2979(n1445 ,n704 ,n1233);
    nand g2980(n2427 ,n2136 ,n2125);
    or g2981(n607 ,n3[11] ,n467);
    nand g2982(n1538 ,n2[85] ,n1253);
    nand g2983(n1012 ,n422 ,n567);
    dff g2984(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2811), .Q(n7[63]));
    xnor g2985(n2318 ,n111 ,n154);
    nand g2986(n1115 ,n2339 ,n652);
    dff g2987(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1972), .Q(n5[37]));
    nand g2988(n1517 ,n737 ,n1338);
    nor g2989(n145 ,n103 ,n144);
    nand g2990(n982 ,n377 ,n479);
    or g2991(n728 ,n2[6] ,n632);
    nand g2992(n1423 ,n675 ,n1211);
    xnor g2993(n2252 ,n2516 ,n2586);
    nand g2994(n1904 ,n1125 ,n1653);
    or g2995(n1348 ,n2[84] ,n1261);
    or g2996(n796 ,n2323 ,n624);
    or g2997(n675 ,n2352 ,n622);
    nand g2998(n1420 ,n697 ,n1207);
    nand g2999(n1893 ,n1115 ,n1642);
    or g3000(n573 ,n4[37] ,n465);
    dff g3001(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1951), .Q(n5[10]));
    nand g3002(n2145 ,n2042 ,n3[16]);
    nand g3003(n2174 ,n2[1] ,n6[1]);
    nor g3004(n1849 ,n948 ,n1783);
    nor g3005(n1794 ,n874 ,n1727);
    nand g3006(n2775 ,n2567 ,n2773);
    xnor g3007(n2343 ,n88 ,n204);
    nor g3008(n151 ,n124 ,n150);
    nor g3009(n1804 ,n883 ,n1737);
    nand g3010(n2396 ,n2235 ,n2104);
    nand g3011(n2499 ,n2242 ,n2164);
    nand g3012(n1037 ,n4[40] ,n639);
    nand g3013(n1089 ,n2[59] ,n562);
    nor g3014(n2719 ,n2529 ,n2716);
    dff g3015(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1874), .Q(n3[60]));
    nand g3016(n339 ,n2341 ,n312);
    or g3017(n673 ,n2353 ,n622);
    or g3018(n920 ,n452 ,n486);
    or g3019(n758 ,n2[31] ,n637);
    nand g3020(n2434 ,n2205 ,n2129);
    or g3021(n849 ,n2368 ,n646);
    dff g3022(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n381), .Q(n6[0]));
    nor g3023(n215 ,n94 ,n214);
    nor g3024(n195 ,n79 ,n194);
    nand g3025(n1171 ,n2319 ,n649);
    xnor g3026(n2330 ,n133 ,n178);
    nor g3027(n1633 ,n702 ,n1441);
    or g3028(n582 ,n3[15] ,n467);
    not g3029(n2782 ,n9[18]);
    dff g3030(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2020), .Q(n4[9]));
    dff g3031(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1971), .Q(n3[52]));
    nand g3032(n1127 ,n2[38] ,n559);
    nand g3033(n1133 ,n2[34] ,n559);
    nand g3034(n318 ,n2265 ,n275);
    nand g3035(n396 ,n2326 ,n275);
    nand g3036(n1165 ,n2[15] ,n557);
    dff g3037(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1891), .Q(n3[47]));
    nand g3038(n71 ,n2438 ,n2374);
    nor g3039(n222 ,n58 ,n221);
    nor g3040(n1825 ,n993 ,n1758);
endmodule
