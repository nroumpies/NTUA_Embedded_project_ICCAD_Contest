module top (n0, n1, n2, n3, n4);
    input n0, n1;
    input [31:0] n2;
    input [3:0] n3;
    output [15:0] n4;
    wire n0, n1;
    wire [31:0] n2;
    wire [3:0] n3;
    wire [15:0] n4;
    wire [7:0] n5;
    wire [15:0] n6;
    wire [7:0] n7;
    wire [15:0] n8;
    wire [15:0] n9;
    wire [3:0] n10;
    wire [2:0] n11;
    wire [63:0] n12;
    wire [63:0] n13;
    wire [15:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335;
    nor g0(n117 ,n100 ,n75);
    nor g1(n163 ,n90 ,n125);
    dff g2(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n272), .Q(n11[2]));
    not g3(n73 ,n72);
    or g4(n224 ,n13[9] ,n211);
    nand g5(n166 ,n3[0] ,n129);
    nand g6(n26 ,n18 ,n25);
    dff g7(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[13]), .Q(n14[14]));
    not g8(n48 ,n9[8]);
    dff g9(.RN(n335), .SN(1'b1), .CK(n0), .D(n330), .Q(n13[10]));
    dff g10(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n204), .Q(n7[1]));
    not g11(n85 ,n303);
    dff g12(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n252), .Q(n6[14]));
    nand g13(n190 ,n308 ,n175);
    nand g14(n306 ,n34 ,n32);
    nor g15(n198 ,n11[2] ,n181);
    dff g16(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n118), .Q(n10[3]));
    xnor g17(n4[9] ,n285 ,n6[9]);
    or g18(n215 ,n13[3] ,n211);
    nand g19(n37 ,n7[1] ,n7[0]);
    xor g20(n12[40] ,n2[8] ,n3[0]);
    xor g21(n12[44] ,n2[12] ,n3[0]);
    nor g22(n113 ,n76 ,n8[1]);
    or g23(n314 ,n19 ,n28);
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n134), .Q(n8[0]));
    not g25(n209 ,n208);
    nor g26(n119 ,n109 ,n75);
    nand g27(n233 ,n13[14] ,n212);
    nor g28(n122 ,n99 ,n75);
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n133), .Q(n8[1]));
    xnor g30(n300 ,n9[10] ,n65);
    nand g31(n269 ,n11[1] ,n257);
    or g32(n222 ,n13[11] ,n211);
    dff g33(.RN(n335), .SN(1'b1), .CK(n0), .D(n14[7]), .Q(n14[8]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n271), .Q(n11[1]));
    xor g35(n327 ,n12[39] ,n14[7]);
    xnor g36(n4[7] ,n285 ,n6[7]);
    nand g37(n44 ,n7[5] ,n42);
    nand g38(n60 ,n9[6] ,n59);
    not g39(n124 ,n125);
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n202), .Q(n7[5]));
    nor g41(n139 ,n98 ,n75);
    not g42(n78 ,n292);
    or g43(n221 ,n13[12] ,n211);
    nand g44(n246 ,n11[0] ,n214);
    xor g45(n319 ,n12[46] ,n14[14]);
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n200), .Q(n7[7]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n258), .Q(n6[9]));
    nor g48(n160 ,n88 ,n125);
    nand g49(n240 ,n13[7] ,n212);
    xnor g50(n307 ,n7[7] ,n46);
    xor g51(n331 ,n12[45] ,n14[13]);
    nand g52(n177 ,n112 ,n173);
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n163), .Q(n9[7]));
    or g54(n220 ,n13[13] ,n211);
    nand g55(n283 ,n5[1] ,n281);
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n201), .Q(n7[0]));
    nor g57(n16 ,n9[13] ,n9[12]);
    not g58(n59 ,n58);
    xnor g59(n298 ,n9[8] ,n62);
    nor g60(n154 ,n89 ,n125);
    xnor g61(n310 ,n7[4] ,n41);
    nand g62(n202 ,n180 ,n196);
    nor g63(n134 ,n75 ,n87);
    nand g64(n250 ,n216 ,n231);
    nand g65(n211 ,n1 ,n207);
    nand g66(n266 ,n128 ,n246);
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n264), .Q(n6[4]));
    xnor g68(n305 ,n74 ,n9[15]);
    nand g69(n165 ,n113 ,n115);
    nor g70(n210 ,n126 ,n207);
    dff g71(.RN(n335), .SN(1'b1), .CK(n0), .D(n331), .Q(n13[13]));
    not g72(n247 ,n246);
    nor g73(n281 ,n277 ,n280);
    not g74(n66 ,n65);
    nand g75(n188 ,n7[0] ,n176);
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n255), .Q(n6[0]));
    xor g77(n12[41] ,n2[9] ,n3[1]);
    nor g78(n147 ,n9[0] ,n125);
    dff g79(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[4]), .Q(n14[5]));
    xor g80(n322 ,n12[43] ,n14[11]);
    xor g81(n284 ,n282 ,n315);
    nand g82(n121 ,n11[0] ,n94);
    xor g83(n330 ,n12[42] ,n14[10]);
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n142), .Q(n5[4]));
    or g85(n223 ,n13[10] ,n211);
    nand g86(n189 ,n313 ,n175);
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n120), .Q(n8[6]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n116), .Q(n5[3]));
    not g89(n167 ,n164);
    dff g90(.RN(n335), .SN(1'b1), .CK(n0), .D(n332), .Q(n13[12]));
    nor g91(n132 ,n108 ,n75);
    or g92(n146 ,n315 ,n121);
    xnor g93(n311 ,n7[3] ,n39);
    nand g94(n200 ,n182 ,n192);
    dff g95(.RN(n335), .SN(1'b1), .CK(n0), .D(n316), .Q(n13[0]));
    xor g96(n12[35] ,n2[3] ,n3[3]);
    nor g97(n276 ,n289 ,n5[0]);
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n160), .Q(n9[14]));
    nor g99(n291 ,n52 ,n50);
    nand g100(n179 ,n7[1] ,n176);
    nor g101(n42 ,n35 ,n41);
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n119), .Q(n10[2]));
    dff g103(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[2]), .Q(n14[3]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n248), .Q(n6[11]));
    nand g105(n69 ,n9[11] ,n68);
    nand g106(n242 ,n13[5] ,n212);
    xnor g107(n4[8] ,n285 ,n6[8]);
    not g108(n95 ,n11[0]);
    xor g109(n12[32] ,n2[0] ,n3[0]);
    nor g110(n175 ,n75 ,n168);
    not g111(n335 ,n1);
    xnor g112(n301 ,n9[11] ,n67);
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n136), .Q(n5[6]));
    not g114(n108 ,n8[1]);
    nor g115(n71 ,n9[13] ,n70);
    not g116(n76 ,n8[2]);
    xnor g117(n4[5] ,n285 ,n6[5]);
    nand g118(n253 ,n220 ,n234);
    nor g119(n131 ,n76 ,n75);
    nand g120(n74 ,n9[14] ,n73);
    nor g121(n181 ,n174 ,n170);
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n130), .Q(n8[4]));
    nand g123(n237 ,n13[10] ,n212);
    dff g124(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[10]), .Q(n14[11]));
    nor g125(n153 ,n91 ,n125);
    xor g126(n334 ,n325 ,n326);
    xor g127(n12[36] ,n2[4] ,n3[0]);
    nor g128(n141 ,n77 ,n75);
    nor g129(n149 ,n92 ,n125);
    xnor g130(n4[6] ,n285 ,n6[6]);
    dff g131(.RN(n335), .SN(1'b1), .CK(n0), .D(n14[0]), .Q(n14[1]));
    dff g132(.RN(n335), .SN(1'b1), .CK(n0), .D(n320), .Q(n13[3]));
    dff g133(.RN(n335), .SN(1'b1), .CK(n0), .D(n328), .Q(n13[6]));
    xor g134(n12[46] ,n2[14] ,n3[2]);
    not g135(n102 ,n8[4]);
    xnor g136(n293 ,n9[3] ,n53);
    xnor g137(n296 ,n9[6] ,n58);
    xnor g138(n294 ,n9[4] ,n55);
    nor g139(n133 ,n97 ,n75);
    dff g140(.RN(n335), .SN(1'b1), .CK(n0), .D(n327), .Q(n13[7]));
    xnor g141(n278 ,n10[0] ,n11[0]);
    nor g142(n155 ,n83 ,n125);
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n141), .Q(n5[2]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n199), .Q(n7[6]));
    nand g145(n199 ,n185 ,n190);
    nor g146(n17 ,n9[10] ,n9[9]);
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n127), .Q(n5[0]));
    nand g148(n245 ,n13[2] ,n212);
    or g149(n123 ,n8[7] ,n11[1]);
    xor g150(n318 ,n12[47] ,n14[15]);
    nand g151(n41 ,n7[3] ,n40);
    nand g152(n272 ,n191 ,n269);
    xor g153(n317 ,n12[36] ,n14[4]);
    nand g154(n280 ,n276 ,n275);
    nor g155(n197 ,n123 ,n177);
    nor g156(n309 ,n43 ,n45);
    nor g157(n208 ,n183 ,n197);
    nor g158(n267 ,n213 ,n266);
    xor g159(n320 ,n12[35] ,n14[3]);
    nand g160(n235 ,n13[12] ,n212);
    nor g161(n270 ,n94 ,n266);
    xnor g162(n302 ,n9[12] ,n69);
    nor g163(n213 ,n11[0] ,n209);
    nand g164(n248 ,n222 ,n236);
    nand g165(n194 ,n311 ,n175);
    not g166(n127 ,n126);
    nor g167(n150 ,n80 ,n125);
    xor g168(n324 ,n12[37] ,n14[5]);
    nor g169(n118 ,n107 ,n75);
    xor g170(n12[42] ,n2[10] ,n3[2]);
    xor g171(n12[38] ,n2[6] ,n3[2]);
    nor g172(n50 ,n9[1] ,n9[0]);
    or g173(n226 ,n13[7] ,n211);
    nand g174(n58 ,n9[5] ,n56);
    nand g175(n39 ,n7[2] ,n38);
    dff g176(.RN(n335), .SN(1'b1), .CK(n0), .D(n324), .Q(n13[5]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n259), .Q(n6[8]));
    xor g178(n316 ,n12[32] ,n14[0]);
    not g179(n54 ,n53);
    nand g180(n234 ,n13[13] ,n212);
    dff g181(.RN(n335), .SN(1'b1), .CK(n0), .D(n318), .Q(n13[15]));
    nand g182(n204 ,n179 ,n189);
    not g183(n81 ,n300);
    nand g184(n137 ,n11[1] ,n314);
    or g185(n229 ,n13[4] ,n211);
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n251), .Q(n6[15]));
    nand g187(n164 ,n145 ,n114);
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n203), .Q(n7[4]));
    nor g189(n143 ,n111 ,n75);
    nand g190(n72 ,n9[13] ,n70);
    or g191(n227 ,n13[6] ,n211);
    nand g192(n249 ,n230 ,n245);
    not g193(n286 ,n5[2]);
    nand g194(n191 ,n315 ,n175);
    nand g195(n55 ,n9[3] ,n54);
    not g196(n84 ,n293);
    not g197(n83 ,n294);
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n265), .Q(n6[10]));
    not g199(n91 ,n298);
    or g200(n148 ,n290 ,n135);
    nor g201(n159 ,n82 ,n125);
    nor g202(n275 ,n288 ,n5[4]);
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n155), .Q(n9[4]));
    nand g204(n214 ,n137 ,n208);
    nand g205(n34 ,n7[3] ,n33);
    not g206(n98 ,n10[0]);
    not g207(n35 ,n7[4]);
    nand g208(n192 ,n307 ,n175);
    xnor g209(n4[3] ,n285 ,n6[3]);
    dff g210(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[14]), .Q(n14[15]));
    not g211(n99 ,n8[6]);
    nor g212(n136 ,n110 ,n75);
    nor g213(n217 ,n13[0] ,n211);
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n263), .Q(n6[5]));
    or g215(n172 ,n138 ,n148);
    not g216(n86 ,n291);
    nand g217(n232 ,n13[15] ,n212);
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n152), .Q(n9[10]));
    xor g219(n12[47] ,n2[15] ,n3[3]);
    dff g220(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n267), .Q(n11[0]));
    nor g221(n313 ,n38 ,n36);
    nor g222(n162 ,n85 ,n125);
    nand g223(n62 ,n9[7] ,n61);
    not g224(n80 ,n302);
    nand g225(n67 ,n9[10] ,n66);
    dff g226(.RN(1'b1), .SN(n335), .CK(n0), .D(n334), .Q(n14[0]));
    nor g227(n120 ,n106 ,n75);
    xnor g228(n4[2] ,n285 ,n6[2]);
    nand g229(n203 ,n184 ,n193);
    nor g230(n56 ,n47 ,n55);
    nand g231(n201 ,n188 ,n178);
    xor g232(n12[37] ,n2[5] ,n3[1]);
    nand g233(n65 ,n9[9] ,n63);
    nand g234(n21 ,n17 ,n15);
    not g235(n89 ,n295);
    not g236(n52 ,n51);
    nand g237(n238 ,n13[9] ,n212);
    nand g238(n24 ,n20 ,n23);
    nor g239(n57 ,n9[5] ,n56);
    not g240(n104 ,n8[3]);
    not g241(n47 ,n9[4]);
    nor g242(n174 ,n94 ,n167);
    nor g243(n115 ,n102 ,n8[3]);
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n131), .Q(n8[3]));
    nand g245(n259 ,n225 ,n239);
    not g246(n68 ,n67);
    nor g247(n158 ,n86 ,n125);
    nand g248(n261 ,n227 ,n241);
    nand g249(n125 ,n1 ,n3[0]);
    dff g250(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[11]), .Q(n14[12]));
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n158), .Q(n9[1]));
    nand g252(n170 ,n146 ,n166);
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n122), .Q(n8[7]));
    not g254(n92 ,n305);
    nand g255(n186 ,n7[2] ,n176);
    nand g256(n290 ,n10[0] ,n273);
    not g257(n287 ,n5[6]);
    nand g258(n252 ,n219 ,n233);
    nor g259(n36 ,n7[1] ,n7[0]);
    xnor g260(n308 ,n7[6] ,n44);
    nor g261(n212 ,n75 ,n207);
    xnor g262(n304 ,n9[14] ,n72);
    or g263(n225 ,n13[8] ,n211);
    nand g264(n231 ,n13[1] ,n212);
    dff g265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n205), .Q(n7[2]));
    dff g266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n162), .Q(n9[13]));
    xor g267(n332 ,n12[44] ,n14[12]);
    not g268(n77 ,n5[1]);
    dff g269(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[6]), .Q(n14[7]));
    nor g270(n25 ,n9[0] ,n24);
    not g271(n45 ,n44);
    or g272(n228 ,n13[5] ,n211);
    xnor g273(n4[10] ,n285 ,n6[10]);
    dff g274(.RN(n335), .SN(1'b1), .CK(n0), .D(n319), .Q(n13[14]));
    not g275(n103 ,n5[2]);
    xnor g276(n4[11] ,n285 ,n6[11]);
    xnor g277(n282 ,n278 ,n7[0]);
    or g278(n33 ,n7[0] ,n30);
    not g279(n109 ,n10[1]);
    dff g280(.RN(n335), .SN(1'b1), .CK(n0), .D(n321), .Q(n13[2]));
    nor g281(n129 ,n11[0] ,n11[1]);
    or g282(n230 ,n13[2] ,n211);
    xnor g283(n292 ,n9[2] ,n51);
    not g284(n111 ,n5[6]);
    nor g285(n128 ,n75 ,n11[2]);
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n124), .Q(n10[0]));
    dff g287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n149), .Q(n9[15]));
    nand g288(n187 ,n7[3] ,n176);
    dff g289(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[1]), .Q(n14[2]));
    not g290(n38 ,n37);
    nor g291(n151 ,n79 ,n125);
    nand g292(n243 ,n13[4] ,n212);
    nor g293(n176 ,n75 ,n169);
    not g294(n100 ,n5[0]);
    nand g295(n135 ,n10[1] ,n10[2]);
    xnor g296(n4[1] ,n285 ,n6[1]);
    dff g297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n250), .Q(n6[1]));
    nor g298(n152 ,n81 ,n125);
    or g299(n30 ,n7[2] ,n7[1]);
    xnor g300(n4[4] ,n285 ,n6[4]);
    xnor g301(n312 ,n7[2] ,n37);
    or g302(n315 ,n274 ,n283);
    nand g303(n265 ,n223 ,n237);
    dff g304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n261), .Q(n6[6]));
    not g305(n273 ,n11[0]);
    dff g306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n260), .Q(n6[7]));
    dff g307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n117), .Q(n5[1]));
    nand g308(n264 ,n229 ,n243);
    dff g309(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n253), .Q(n6[13]));
    nor g310(n112 ,n99 ,n8[5]);
    not g311(n40 ,n39);
    dff g312(.RN(n335), .SN(1'b1), .CK(n0), .D(n329), .Q(n13[8]));
    dff g313(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n153), .Q(n9[8]));
    xor g314(n12[43] ,n2[11] ,n3[3]);
    or g315(n19 ,n9[15] ,n9[14]);
    not g316(n93 ,n296);
    dff g317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n150), .Q(n9[12]));
    nand g318(n27 ,n9[11] ,n26);
    not g319(n96 ,n7[0]);
    not g320(n87 ,n2[0]);
    xnor g321(n4[13] ,n285 ,n6[13]);
    nand g322(n193 ,n310 ,n175);
    not g323(n90 ,n297);
    xnor g324(n297 ,n9[7] ,n60);
    nor g325(n299 ,n64 ,n66);
    not g326(n257 ,n256);
    nand g327(n126 ,n1 ,n13[0]);
    or g328(n218 ,n13[15] ,n211);
    dff g329(.RN(n335), .SN(1'b1), .CK(n0), .D(n14[3]), .Q(n14[4]));
    nand g330(n262 ,n215 ,n244);
    not g331(n97 ,n8[0]);
    not g332(n107 ,n10[2]);
    dff g333(.RN(n335), .SN(1'b1), .CK(n0), .D(n14[12]), .Q(n14[13]));
    dff g334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n132), .Q(n8[2]));
    dff g335(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n154), .Q(n9[5]));
    dff g336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n156), .Q(n9[3]));
    not g337(n79 ,n301);
    not g338(n169 ,n168);
    nand g339(n53 ,n9[2] ,n52);
    xnor g340(n279 ,n8[0] ,n9[0]);
    xnor g341(n326 ,n14[10] ,n14[12]);
    nand g342(n236 ,n13[11] ,n212);
    nor g343(n171 ,n98 ,n168);
    dff g344(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n144), .Q(n8[5]));
    nand g345(n256 ,n128 ,n247);
    xor g346(n12[39] ,n2[7] ,n3[3]);
    dff g347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n262), .Q(n6[3]));
    nand g348(n178 ,n96 ,n175);
    nor g349(n43 ,n7[5] ,n42);
    nor g350(n64 ,n9[9] ,n63);
    dff g351(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n143), .Q(n5[7]));
    xor g352(n328 ,n12[38] ,n14[6]);
    dff g353(.RN(n335), .SN(1'b1), .CK(n0), .D(n317), .Q(n13[4]));
    nand g354(n182 ,n7[7] ,n176);
    nand g355(n277 ,n5[7] ,n287);
    nand g356(n185 ,n7[6] ,n176);
    xor g357(n323 ,n12[33] ,n14[1]);
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n157), .Q(n9[2]));
    nor g359(n23 ,n9[5] ,n22);
    or g360(n255 ,n210 ,n217);
    nand g361(n251 ,n218 ,n232);
    nor g362(n116 ,n103 ,n75);
    nor g363(n303 ,n71 ,n73);
    not g364(n94 ,n11[1]);
    nor g365(n140 ,n101 ,n75);
    dff g366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n206), .Q(n7[3]));
    not g367(n49 ,n9[12]);
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n249), .Q(n6[2]));
    nand g369(n183 ,n166 ,n172);
    dff g370(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n147), .Q(n9[0]));
    nor g371(n63 ,n48 ,n62);
    dff g372(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n254), .Q(n6[12]));
    dff g373(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n140), .Q(n5[5]));
    dff g374(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n161), .Q(n9[6]));
    or g375(n207 ,n171 ,n198);
    not g376(n288 ,n5[5]);
    xnor g377(n4[15] ,n285 ,n6[15]);
    nor g378(n157 ,n78 ,n125);
    nor g379(n268 ,n11[1] ,n256);
    xor g380(n12[45] ,n2[13] ,n3[1]);
    xor g381(n329 ,n12[40] ,n14[8]);
    nand g382(n254 ,n221 ,n235);
    xnor g383(n4[14] ,n285 ,n6[14]);
    not g384(n105 ,n5[3]);
    or g385(n22 ,n9[4] ,n21);
    nor g386(n70 ,n49 ,n69);
    nor g387(n18 ,n9[2] ,n9[1]);
    nand g388(n274 ,n5[3] ,n286);
    dff g389(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[9]), .Q(n14[10]));
    nand g390(n195 ,n312 ,n175);
    dff g391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n151), .Q(n9[11]));
    nor g392(n295 ,n57 ,n59);
    or g393(n219 ,n13[14] ,n211);
    nor g394(n15 ,n9[8] ,n9[7]);
    xor g395(n12[34] ,n2[2] ,n3[2]);
    nor g396(n142 ,n105 ,n75);
    not g397(n106 ,n8[5]);
    xor g398(n321 ,n12[34] ,n14[2]);
    or g399(n271 ,n270 ,n268);
    nand g400(n263 ,n228 ,n242);
    nor g401(n32 ,n31 ,n29);
    nor g402(n161 ,n93 ,n125);
    nor g403(n173 ,n145 ,n165);
    not g404(n61 ,n60);
    nor g405(n130 ,n104 ,n75);
    nand g406(n260 ,n226 ,n240);
    nand g407(n145 ,n8[0] ,n11[0]);
    nor g408(n144 ,n102 ,n75);
    or g409(n29 ,n7[5] ,n7[4]);
    or g410(n31 ,n7[7] ,n7[6]);
    nand g411(n196 ,n309 ,n175);
    nand g412(n51 ,n9[1] ,n9[0]);
    nand g413(n205 ,n186 ,n195);
    nand g414(n138 ,n10[3] ,n11[1]);
    not g415(n88 ,n304);
    xnor g416(n285 ,n279 ,n284);
    not g417(n101 ,n5[4]);
    nand g418(n114 ,n9[0] ,n95);
    or g419(n216 ,n13[1] ,n211);
    xnor g420(n325 ,n14[13] ,n14[15]);
    nand g421(n206 ,n187 ,n194);
    not g422(n289 ,n306);
    nand g423(n180 ,n7[5] ,n176);
    nand g424(n244 ,n13[3] ,n212);
    xnor g425(n4[0] ,n285 ,n6[0]);
    xnor g426(n4[12] ,n285 ,n6[12]);
    not g427(n75 ,n1);
    nand g428(n28 ,n16 ,n27);
    dff g429(.RN(n335), .SN(1'b1), .CK(n0), .D(n14[5]), .Q(n14[6]));
    nand g430(n184 ,n7[4] ,n176);
    nor g431(n156 ,n84 ,n125);
    dff g432(.RN(n335), .SN(1'b1), .CK(n0), .D(n322), .Q(n13[11]));
    dff g433(.RN(n335), .SN(1'b1), .CK(n0), .D(n323), .Q(n13[1]));
    nand g434(n239 ,n13[8] ,n212);
    nand g435(n46 ,n7[6] ,n45);
    dff g436(.RN(1'b1), .SN(n335), .CK(n0), .D(n14[8]), .Q(n14[9]));
    xor g437(n12[33] ,n2[1] ,n3[1]);
    nor g438(n20 ,n9[6] ,n9[3]);
    dff g439(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n139), .Q(n10[1]));
    not g440(n110 ,n5[5]);
    nand g441(n258 ,n224 ,n238);
    nand g442(n168 ,n11[2] ,n129);
    dff g443(.RN(n335), .SN(1'b1), .CK(n0), .D(n333), .Q(n13[9]));
    dff g444(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n159), .Q(n9[9]));
    xor g445(n333 ,n12[41] ,n14[9]);
    nand g446(n241 ,n13[6] ,n212);
    not g447(n82 ,n299);
endmodule
