module top (n0, n1, n4, n6, n5, n2, n11, n12, n13, n14, n17, n15, n16, n3, n7, n8, n9, n10);
    input n0, n1, n2, n3;
    input [7:0] n4;
    input [3:0] n5;
    output [7:0] n6, n7, n8, n9, n10;
    output n11, n12, n13, n14, n15, n16;
    output [3:0] n17;
    wire n0, n1, n2, n3;
    wire [7:0] n4;
    wire [3:0] n5;
    wire [7:0] n6, n7, n8, n9, n10;
    wire n11, n12, n13, n14, n15, n16;
    wire [3:0] n17;
    wire [3:0] n18;
    wire [3:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [7:0] n23;
    wire [7:0] n24;
    wire [7:0] n25;
    wire [7:0] n26;
    wire [7:0] n27;
    wire [7:0] n28;
    wire [7:0] n29;
    wire [7:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [4:0] n36;
    wire [3:0] n37;
    wire [3:0] n38;
    wire [7:0] n39;
    wire [2:0] n40;
    wire [7:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [7:0] n44;
    wire [7:0] n45;
    wire [7:0] n46;
    wire [7:0] n47;
    wire [7:0] n48;
    wire [7:0] n49;
    wire [7:0] n50;
    wire [7:0] n51;
    wire [7:0] n52;
    wire [7:0] n53;
    wire [7:0] n54;
    wire [7:0] n55;
    wire [7:0] n56;
    wire [4:0] n57;
    wire [3:0] n58;
    wire [3:0] n59;
    wire [7:0] n60;
    wire n61, n62, n63, n64, n65, n66, n67, n68;
    wire n69, n70, n71, n72, n73, n74, n75, n76;
    wire n77, n78, n79, n80, n81, n82, n83, n84;
    wire n85, n86, n87, n88, n89, n90, n91, n92;
    wire n93, n94, n95, n96, n97, n98, n99, n100;
    wire n101, n102, n103, n104, n105, n106, n107, n108;
    wire n109, n110, n111, n112, n113, n114, n115, n116;
    wire n117, n118, n119, n120, n121, n122, n123, n124;
    wire n125, n126, n127, n128, n129, n130, n131, n132;
    wire n133, n134, n135, n136, n137, n138, n139, n140;
    wire n141, n142, n143, n144, n145, n146, n147, n148;
    wire n149, n150, n151, n152, n153, n154, n155, n156;
    wire n157, n158, n159, n160, n161, n162, n163, n164;
    wire n165, n166, n167, n168, n169, n170, n171, n172;
    wire n173, n174, n175, n176, n177, n178, n179, n180;
    wire n181, n182, n183, n184, n185, n186, n187, n188;
    wire n189, n190, n191, n192, n193, n194, n195, n196;
    wire n197, n198, n199, n200, n201, n202, n203, n204;
    wire n205, n206, n207, n208, n209, n210, n211, n212;
    wire n213, n214, n215, n216, n217, n218, n219, n220;
    wire n221, n222, n223, n224, n225, n226, n227, n228;
    wire n229, n230, n231, n232, n233, n234, n235, n236;
    wire n237, n238, n239, n240, n241, n242, n243, n244;
    wire n245, n246, n247, n248, n249, n250, n251, n252;
    wire n253, n254, n255, n256, n257, n258, n259, n260;
    wire n261, n262, n263, n264, n265, n266, n267, n268;
    wire n269, n270, n271, n272, n273, n274, n275, n276;
    wire n277, n278, n279, n280, n281, n282, n283, n284;
    wire n285, n286, n287, n288, n289, n290, n291, n292;
    wire n293, n294, n295, n296, n297, n298, n299, n300;
    wire n301, n302, n303, n304, n305, n306, n307, n308;
    wire n309, n310, n311, n312, n313, n314, n315, n316;
    wire n317, n318, n319, n320, n321, n322, n323, n324;
    wire n325, n326, n327, n328, n329, n330, n331, n332;
    wire n333, n334, n335, n336, n337, n338, n339, n340;
    wire n341, n342, n343, n344, n345, n346, n347, n348;
    wire n349, n350, n351, n352, n353, n354, n355, n356;
    wire n357, n358, n359, n360, n361, n362, n363, n364;
    wire n365, n366, n367, n368, n369, n370, n371, n372;
    wire n373, n374, n375, n376, n377, n378, n379, n380;
    wire n381, n382, n383, n384, n385, n386, n387, n388;
    wire n389, n390, n391, n392, n393, n394, n395, n396;
    wire n397, n398, n399, n400, n401, n402, n403, n404;
    wire n405, n406, n407, n408, n409, n410, n411, n412;
    wire n413, n414, n415, n416, n417, n418, n419, n420;
    wire n421, n422, n423, n424, n425, n426, n427, n428;
    wire n429, n430, n431, n432, n433, n434, n435, n436;
    wire n437, n438, n439, n440, n441, n442, n443, n444;
    wire n445, n446, n447, n448, n449, n450, n451, n452;
    wire n453, n454, n455, n456, n457, n458, n459, n460;
    wire n461, n462, n463, n464, n465, n466, n467, n468;
    wire n469, n470, n471, n472, n473, n474, n475, n476;
    wire n477, n478, n479, n480, n481, n482, n483, n484;
    wire n485, n486, n487, n488, n489, n490, n491, n492;
    wire n493, n494, n495, n496, n497, n498, n499, n500;
    wire n501, n502, n503, n504, n505, n506, n507, n508;
    wire n509, n510, n511, n512, n513, n514, n515, n516;
    wire n517, n518, n519, n520, n521, n522, n523, n524;
    wire n525, n526, n527, n528, n529, n530, n531, n532;
    wire n533, n534, n535, n536, n537, n538, n539, n540;
    wire n541, n542, n543, n544, n545, n546, n547, n548;
    wire n549, n550, n551, n552, n553, n554, n555, n556;
    wire n557, n558, n559, n560, n561, n562, n563, n564;
    wire n565, n566, n567, n568, n569, n570, n571, n572;
    wire n573, n574, n575, n576, n577, n578, n579, n580;
    wire n581, n582, n583, n584, n585, n586, n587, n588;
    wire n589, n590, n591, n592, n593, n594, n595, n596;
    wire n597, n598, n599, n600, n601, n602, n603, n604;
    wire n605, n606, n607, n608, n609, n610, n611, n612;
    wire n613, n614, n615, n616, n617, n618, n619, n620;
    wire n621, n622, n623, n624, n625, n626, n627, n628;
    wire n629, n630, n631, n632, n633, n634, n635, n636;
    wire n637, n638, n639, n640, n641, n642, n643, n644;
    wire n645, n646, n647, n648, n649, n650, n651, n652;
    wire n653, n654, n655, n656, n657, n658, n659, n660;
    wire n661, n662, n663, n664, n665, n666, n667, n668;
    wire n669, n670, n671, n672, n673, n674, n675, n676;
    wire n677, n678, n679, n680, n681, n682, n683, n684;
    wire n685, n686, n687, n688, n689, n690, n691, n692;
    wire n693, n694, n695, n696, n697, n698, n699, n700;
    wire n701, n702, n703, n704, n705, n706, n707, n708;
    wire n709, n710, n711, n712, n713, n714, n715, n716;
    wire n717, n718, n719, n720, n721, n722, n723, n724;
    wire n725, n726, n727, n728, n729, n730, n731, n732;
    wire n733, n734, n735, n736, n737, n738, n739, n740;
    wire n741, n742, n743, n744, n745, n746, n747, n748;
    wire n749, n750, n751, n752, n753, n754, n755, n756;
    wire n757, n758, n759, n760, n761, n762, n763, n764;
    wire n765, n766, n767, n768, n769, n770, n771, n772;
    wire n773, n774, n775, n776, n777, n778, n779, n780;
    wire n781, n782, n783, n784, n785, n786, n787, n788;
    wire n789, n790, n791, n792, n793, n794, n795, n796;
    wire n797, n798, n799, n800, n801, n802, n803, n804;
    wire n805, n806, n807, n808, n809, n810, n811, n812;
    wire n813, n814, n815, n816, n817, n818, n819, n820;
    wire n821, n822, n823, n824, n825, n826, n827, n828;
    wire n829, n830, n831, n832, n833, n834, n835, n836;
    wire n837, n838, n839, n840, n841, n842, n843, n844;
    wire n845, n846, n847, n848, n849, n850, n851, n852;
    wire n853, n854, n855, n856, n857, n858, n859, n860;
    wire n861, n862, n863, n864, n865, n866, n867, n868;
    wire n869, n870, n871, n872, n873, n874, n875, n876;
    wire n877, n878, n879, n880, n881, n882, n883, n884;
    wire n885, n886, n887, n888, n889, n890, n891, n892;
    wire n893, n894, n895, n896, n897, n898, n899, n900;
    wire n901, n902, n903, n904, n905, n906, n907, n908;
    wire n909, n910, n911, n912, n913, n914, n915, n916;
    wire n917, n918, n919, n920, n921, n922, n923, n924;
    wire n925, n926, n927, n928, n929, n930, n931, n932;
    wire n933, n934, n935, n936, n937, n938, n939, n940;
    wire n941, n942, n943, n944, n945, n946, n947, n948;
    wire n949, n950, n951, n952, n953, n954, n955, n956;
    wire n957, n958, n959, n960, n961, n962, n963, n964;
    wire n965, n966, n967, n968, n969, n970, n971, n972;
    wire n973, n974, n975, n976, n977, n978, n979, n980;
    wire n981, n982, n983, n984, n985, n986, n987, n988;
    wire n989, n990, n991, n992, n993, n994, n995, n996;
    wire n997, n998, n999, n1000, n1001, n1002, n1003, n1004;
    wire n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012;
    wire n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
    wire n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
    wire n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
    wire n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044;
    wire n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
    wire n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060;
    wire n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068;
    wire n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076;
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084;
    wire n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092;
    wire n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100;
    wire n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108;
    wire n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116;
    wire n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124;
    wire n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132;
    wire n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140;
    wire n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148;
    wire n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156;
    wire n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164;
    wire n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172;
    wire n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180;
    wire n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188;
    wire n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196;
    wire n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204;
    wire n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
    wire n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220;
    wire n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228;
    wire n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236;
    wire n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244;
    wire n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252;
    wire n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260;
    wire n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268;
    wire n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276;
    wire n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284;
    wire n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292;
    wire n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300;
    wire n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308;
    wire n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;
    wire n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;
    wire n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332;
    wire n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340;
    wire n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348;
    wire n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356;
    wire n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364;
    wire n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372;
    wire n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380;
    wire n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388;
    wire n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;
    wire n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404;
    wire n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412;
    wire n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;
    wire n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428;
    wire n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436;
    wire n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444;
    wire n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452;
    wire n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;
    wire n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468;
    wire n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476;
    wire n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
    wire n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492;
    wire n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500;
    wire n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508;
    wire n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516;
    wire n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524;
    wire n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532;
    wire n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540;
    wire n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548;
    wire n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556;
    wire n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564;
    wire n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572;
    wire n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580;
    wire n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588;
    wire n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596;
    wire n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604;
    wire n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612;
    wire n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620;
    wire n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628;
    wire n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636;
    wire n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644;
    wire n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652;
    wire n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660;
    wire n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668;
    wire n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676;
    wire n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684;
    wire n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692;
    wire n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700;
    wire n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708;
    wire n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716;
    wire n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724;
    wire n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732;
    wire n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740;
    wire n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748;
    wire n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756;
    wire n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764;
    wire n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772;
    wire n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780;
    wire n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788;
    wire n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796;
    wire n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804;
    wire n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812;
    wire n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820;
    wire n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828;
    wire n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836;
    wire n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844;
    wire n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852;
    wire n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860;
    wire n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868;
    wire n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876;
    wire n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884;
    wire n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892;
    wire n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900;
    wire n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908;
    wire n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916;
    wire n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924;
    wire n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932;
    wire n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940;
    wire n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948;
    wire n1949, n1950, n1951, n1952, n1953, n1954, n1955;
    dff g0(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1917), .Q(n6[0]));
    dff g1(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1737), .Q(n26[5]));
    nand g2(n761 ,n46[5] ,n485);
    nor g3(n1939 ,n87 ,n85);
    nand g4(n461 ,n6[6] ,n310);
    buf g5(n8[5], 1'b0);
    nand g6(n1501 ,n35[0] ,n1087);
    nor g7(n154 ,n111 ,n4[0]);
    nand g8(n1679 ,n436 ,n1083);
    or g9(n279 ,n38[3] ,n223);
    nand g10(n265 ,n15 ,n216);
    dff g11(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1883), .Q(n60[4]));
    not g12(n948 ,n826);
    nand g13(n1778 ,n1505 ,n1381);
    nand g14(n1732 ,n1450 ,n1361);
    nor g15(n1900 ,n1191 ,n1889);
    or g16(n1101 ,n425 ,n722);
    not g17(n127 ,n5[2]);
    nand g18(n1056 ,n4[4] ,n708);
    dff g19(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1629), .Q(n45[6]));
    nand g20(n1820 ,n1557 ,n1278);
    nand g21(n609 ,n24[0] ,n410);
    or g22(n1714 ,n1206 ,n1335);
    or g23(n1346 ,n1125 ,n1234);
    or g24(n258 ,n111 ,n206);
    nand g25(n554 ,n45[0] ,n397);
    nand g26(n1017 ,n4[2] ,n720);
    nand g27(n682 ,n51[2] ,n401);
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1663), .Q(n41[7]));
    nand g29(n1384 ,n176 ,n1090);
    nand g30(n90 ,n57[3] ,n89);
    nand g31(n849 ,n47[1] ,n417);
    nand g32(n837 ,n42[2] ,n475);
    nand g33(n1051 ,n4[2] ,n713);
    nand g34(n355 ,n38[1] ,n263);
    nand g35(n1013 ,n4[7] ,n720);
    nor g36(n486 ,n231 ,n347);
    nand g37(n166 ,n40[0] ,n1);
    nand g38(n191 ,n19[1] ,n38[0]);
    nand g39(n1249 ,n735 ,n909);
    nand g40(n1137 ,n615 ,n612);
    nand g41(n1604 ,n1057 ,n589);
    nand g42(n861 ,n22[1] ,n409);
    not g43(n120 ,n18[0]);
    nand g44(n1648 ,n990 ,n635);
    nand g45(n1822 ,n1561 ,n1267);
    nand g46(n1239 ,n934 ,n947);
    nand g47(n581 ,n50[2] ,n380);
    nor g48(n394 ,n237 ,n344);
    nand g49(n1005 ,n4[7] ,n718);
    nand g50(n1495 ,n35[6] ,n1087);
    nand g51(n1597 ,n1086 ,n532);
    nand g52(n1138 ,n894 ,n817);
    nor g53(n1906 ,n1241 ,n1881);
    nand g54(n1190 ,n869 ,n677);
    nand g55(n733 ,n22[5] ,n409);
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1817), .Q(n29[5]));
    nand g57(n1692 ,n447 ,n1082);
    nand g58(n1831 ,n1649 ,n1300);
    nand g59(n744 ,n44[7] ,n478);
    nand g60(n1039 ,n4[1] ,n711);
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1803), .Q(n31[3]));
    nand g62(n735 ,n29[5] ,n407);
    nor g63(n325 ,n119 ,n254);
    nand g64(n700 ,n56[7] ,n378);
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1771), .Q(n22[3]));
    nand g66(n1796 ,n1523 ,n1415);
    nand g67(n1455 ,n26[4] ,n1103);
    nand g68(n1063 ,n4[4] ,n707);
    buf g69(n9[7], 1'b0);
    nand g70(n1023 ,n4[2] ,n719);
    nand g71(n1767 ,n1486 ,n1428);
    nand g72(n546 ,n54[4] ,n392);
    nand g73(n1887 ,n878 ,n1860);
    nand g74(n1672 ,n1004 ,n657);
    nand g75(n929 ,n29[1] ,n407);
    nand g76(n1197 ,n895 ,n623);
    buf g77(n7[0], 1'b0);
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1600), .Q(n49[7]));
    nand g79(n1624 ,n966 ,n793);
    nor g80(n1327 ,n1160 ,n1190);
    nand g81(n881 ,n42[4] ,n475);
    nand g82(n94 ,n59[2] ,n93);
    nor g83(n402 ,n233 ,n351);
    nand g84(n522 ,n153 ,n383);
    nand g85(n886 ,n48[6] ,n395);
    nand g86(n1439 ,n30[4] ,n1094);
    or g87(n1315 ,n173 ,n1105);
    not g88(n87 ,n86);
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1909), .Q(n6[4]));
    nand g90(n775 ,n48[3] ,n483);
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n287), .Q(n7[5]));
    nand g92(n1382 ,n170 ,n1090);
    nand g93(n1240 ,n461 ,n699);
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1535), .Q(n56[7]));
    nor g95(n274 ,n125 ,n230);
    nor g96(n419 ,n220 ,n311);
    nand g97(n1602 ,n1055 ,n680);
    nand g98(n221 ,n129 ,n163);
    nand g99(n469 ,n334 ,n330);
    nand g100(n903 ,n53[5] ,n408);
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1828), .Q(n28[2]));
    nand g102(n1947 ,n62 ,n61);
    nor g103(n1286 ,n1245 ,n1251);
    nand g104(n1456 ,n26[3] ,n1103);
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1626), .Q(n46[2]));
    nand g106(n323 ,n59[2] ,n252);
    nand g107(n1707 ,n1297 ,n1323);
    nand g108(n781 ,n46[4] ,n485);
    nand g109(n639 ,n43[7] ,n376);
    or g110(n953 ,n508 ,n507);
    nand g111(n1155 ,n201 ,n524);
    nand g112(n1521 ,n32[4] ,n1101);
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1800), .Q(n31[6]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1646), .Q(n43[3]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1799), .Q(n31[7]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n440), .Q(n17[2]));
    nand g117(n1361 ,n180 ,n1092);
    nand g118(n1201 ,n618 ,n785);
    nand g119(n455 ,n60[7] ,n348);
    nand g120(n459 ,n3 ,n321);
    nand g121(n829 ,n42[7] ,n475);
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1589), .Q(n51[4]));
    nand g123(n946 ,n55[7] ,n416);
    or g124(n362 ,n298 ,n291);
    nand g125(n1909 ,n1293 ,n1896);
    nand g126(n892 ,n49[4] ,n418);
    not g127(n131 ,n58[2]);
    nand g128(n513 ,n153 ,n369);
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1692), .Q(n58[3]));
    nor g130(n348 ,n130 ,n265);
    not g131(n189 ,n188);
    nand g132(n630 ,n20[2] ,n405);
    nand g133(n975 ,n4[2] ,n715);
    nor g134(n410 ,n213 ,n346);
    nand g135(n1545 ,n29[7] ,n1097);
    nand g136(n1560 ,n1016 ,n620);
    not g137(n387 ,n388);
    nand g138(n1647 ,n989 ,n634);
    nand g139(n1159 ,n870 ,n871);
    nand g140(n1779 ,n1506 ,n1402);
    nor g141(n151 ,n111 ,n56[0]);
    nand g142(n1514 ,n33[3] ,n1109);
    nand g143(n376 ,n255 ,n314);
    or g144(n510 ,n146 ,n375);
    nand g145(n1734 ,n1451 ,n1265);
    nand g146(n1085 ,n277 ,n703);
    nor g147(n417 ,n238 ,n311);
    or g148(n73 ,n57[4] ,n57[1]);
    nand g149(n1445 ,n27[6] ,n1091);
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1558), .Q(n54[4]));
    nor g151(n313 ,n111 ,n254);
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1756), .Q(n24[2]));
    nand g153(n1827 ,n1573 ,n1285);
    nand g154(n1550 ,n29[5] ,n1097);
    nand g155(n1683 ,n36[3] ,n1110);
    nand g156(n1662 ,n21[1] ,n1095);
    buf g157(n10[0], 1'b0);
    not g158(n128 ,n40[0]);
    nand g159(n999 ,n4[6] ,n709);
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1805), .Q(n31[1]));
    nand g161(n1889 ,n883 ,n1867);
    nand g162(n797 ,n46[1] ,n480);
    or g163(n1102 ,n425 ,n721);
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1619), .Q(n47[2]));
    nand g165(n183 ,n39[6] ,n1);
    xnor g166(n1924 ,n59[3] ,n94);
    nand g167(n742 ,n31[0] ,n402);
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1581), .Q(n52[4]));
    nor g169(n1898 ,n1120 ,n1890);
    xnor g170(n1940 ,n57[2] ,n86);
    nand g171(n1630 ,n972 ,n619);
    nand g172(n1183 ,n599 ,n645);
    buf g173(n8[0], 1'b0);
    nand g174(n664 ,n45[6] ,n397);
    nand g175(n992 ,n4[6] ,n710);
    not g176(n1103 ,n1104);
    nand g177(n556 ,n53[1] ,n370);
    nand g178(n632 ,n43[5] ,n376);
    nand g179(n460 ,n37[2] ,n310);
    nand g180(n1476 ,n23[7] ,n1089);
    nand g181(n1916 ,n1340 ,n1903);
    nand g182(n1505 ,n34[4] ,n1102);
    nor g183(n103 ,n38[1] ,n38[0]);
    nand g184(n831 ,n42[6] ,n475);
    nor g185(n487 ,n214 ,n350);
    nand g186(n1814 ,n1501 ,n1260);
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1632), .Q(n45[3]));
    not g188(n320 ,n319);
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1837), .Q(n21[1]));
    nor g190(n420 ,n111 ,n349);
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1840), .Q(n59[1]));
    nand g192(n1635 ,n977 ,n744);
    nor g193(n356 ,n228 ,n304);
    nor g194(n208 ,n185 ,n190);
    nand g195(n1655 ,n994 ,n881);
    nand g196(n1855 ,n1676 ,n1314);
    nand g197(n1690 ,n1923 ,n1111);
    nand g198(n1594 ,n1006 ,n577);
    nand g199(n1370 ,n178 ,n1107);
    nand g200(n1492 ,n22[0] ,n1108);
    nor g201(n429 ,n111 ,n338);
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1079), .Q(n55[0]));
    nand g203(n1791 ,n1518 ,n1432);
    nand g204(n896 ,n49[3] ,n418);
    nor g205(n263 ,n40[0] ,n212);
    nand g206(n991 ,n4[7] ,n710);
    nand g207(n1253 ,n1928 ,n726);
    nand g208(n374 ,n257 ,n318);
    xnor g209(n1936 ,n36[3] ,n82);
    nand g210(n1913 ,n1344 ,n1906);
    nand g211(n1701 ,n1286 ,n1280);
    nand g212(n650 ,n41[6] ,n372);
    nor g213(n499 ,n154 ,n483);
    not g214(n149 ,n55[0]);
    nand g215(n1169 ,n929 ,n861);
    nand g216(n1817 ,n1550 ,n1275);
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1543), .Q(n55[6]));
    or g218(n512 ,n142 ,n371);
    nand g219(n1176 ,n848 ,n597);
    nand g220(n1775 ,n1502 ,n1430);
    nand g221(n1829 ,n1577 ,n1289);
    nor g222(n1862 ,n1123 ,n1702);
    nand g223(n652 ,n41[5] ,n372);
    not g224(n70 ,n69);
    not g225(n167 ,n166);
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1538), .Q(n56[4]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n271), .Q(n13));
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1667), .Q(n41[4]));
    nand g229(n1425 ,n182 ,n1107);
    nand g230(n1875 ,n756 ,n1718);
    or g231(n1699 ,n1012 ,n1436);
    not g232(n245 ,n246);
    not g233(n270 ,n229);
    nand g234(n1449 ,n27[1] ,n1091);
    not g235(n1921 ,n1938);
    nand g236(n597 ,n41[6] ,n400);
    nand g237(n1187 ,n887 ,n923);
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1823), .Q(n28[7]));
    or g239(n1313 ,n175 ,n1105);
    nand g240(n1571 ,n28[4] ,n1096);
    or g241(n1420 ,n175 ,n1098);
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n727), .Q(n57[3]));
    nand g243(n562 ,n52[5] ,n384);
    nor g244(n206 ,n190 ,n157);
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1727), .Q(n27[7]));
    nor g246(n1337 ,n1250 ,n1208);
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1580), .Q(n52[5]));
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1747), .Q(n25[3]));
    nand g249(n1014 ,n4[6] ,n720);
    or g250(n1260 ,n156 ,n1087);
    nand g251(n1182 ,n525 ,n569);
    nor g252(n291 ,n177 ,n244);
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1653), .Q(n42[6]));
    nor g254(n1092 ,n422 ,n721);
    nand g255(n895 ,n42[4] ,n403);
    nand g256(n344 ,n58[0] ,n248);
    nand g257(n805 ,n50[4] ,n412);
    nand g258(n879 ,n31[1] ,n402);
    nand g259(n1461 ,n25[6] ,n1106);
    nand g260(n1266 ,n23[0] ,n1089);
    nand g261(n184 ,n19[0] ,n19[1]);
    nand g262(n555 ,n27[5] ,n486);
    dff g263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1719), .Q(n30[7]));
    nor g264(n422 ,n111 ,n332);
    nand g265(n106 ,n38[2] ,n105);
    nand g266(n1473 ,n24[2] ,n1099);
    not g267(n251 ,n252);
    nand g268(n1792 ,n1519 ,n1411);
    nand g269(n1763 ,n1480 ,n1385);
    dff g270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1816), .Q(n29[6]));
    dff g271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1910), .Q(n6[3]));
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1833), .Q(n21[5]));
    nand g273(n762 ,n42[3] ,n403);
    nand g274(n1019 ,n4[7] ,n719);
    nand g275(n1001 ,n4[4] ,n709);
    nor g276(n95 ,n37[1] ,n37[0]);
    nand g277(n1077 ,n517 ,n513);
    nand g278(n1458 ,n26[1] ,n1103);
    nand g279(n1470 ,n24[5] ,n1099);
    nand g280(n1500 ,n35[1] ,n1087);
    dff g281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1746), .Q(n25[4]));
    nand g282(n229 ,n166 ,n188);
    dff g283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n960), .Q(n50[0]));
    nor g284(n409 ,n233 ,n346);
    nand g285(n877 ,n44[2] ,n398);
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1569), .Q(n53[5]));
    nand g287(n214 ,n116 ,n164);
    nand g288(n588 ,n43[3] ,n419);
    nor g289(n1088 ,n423 ,n721);
    nand g290(n622 ,n45[3] ,n382);
    nand g291(n1049 ,n4[4] ,n713);
    nand g292(n1480 ,n23[3] ,n1089);
    nor g293(n400 ,n221 ,n311);
    nand g294(n433 ,n37[0] ,n310);
    dff g295(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1633), .Q(n45[2]));
    nand g296(n955 ,n510 ,n506);
    nand g297(n1120 ,n462 ,n573);
    nand g298(n434 ,n58[1] ,n313);
    nand g299(n983 ,n4[1] ,n717);
    nand g300(n779 ,n35[3] ,n481);
    nor g301(n1110 ,n309 ,n704);
    nor g302(n1318 ,n1159 ,n1173);
    nor g303(n365 ,n203 ,n355);
    nor g304(n360 ,n203 ,n353);
    nand g305(n1114 ,n835 ,n555);
    or g306(n1415 ,n181 ,n1101);
    nand g307(n1657 ,n995 ,n836);
    nor g308(n1292 ,n1203 ,n1126);
    nor g309(n440 ,n273 ,n305);
    nand g310(n1812 ,n1499 ,n1401);
    nand g311(n1069 ,n4[6] ,n706);
    not g312(n174 ,n175);
    nand g313(n1661 ,n997 ,n838);
    nand g314(n905 ,n60[7] ,n396);
    nor g315(n416 ,n239 ,n311);
    buf g316(n9[4], 1'b0);
    not g317(n1091 ,n1092);
    nand g318(n596 ,n45[3] ,n397);
    or g319(n366 ,n300 ,n286);
    nand g320(n1559 ,n29[1] ,n1097);
    or g321(n1403 ,n181 ,n1102);
    nand g322(n1516 ,n33[1] ,n1109);
    dff g323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1913), .Q(n60[6]));
    not g324(n474 ,n475);
    nand g325(n1616 ,n1070 ,n602);
    nor g326(n306 ,n17[3] ,n253);
    or g327(n504 ,n137 ,n381);
    not g328(n379 ,n380);
    nand g329(n1457 ,n26[2] ,n1103);
    nand g330(n978 ,n4[6] ,n717);
    nand g331(n678 ,n45[7] ,n397);
    nor g332(n714 ,n186 ,n488);
    or g333(n160 ,n111 ,n36[0]);
    nand g334(n1615 ,n1069 ,n601);
    dff g335(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n956), .Q(n42[0]));
    nand g336(n392 ,n256 ,n317);
    or g337(n317 ,n111 ,n269);
    nand g338(n1830 ,n1582 ,n1268);
    nand g339(n924 ,n30[1] ,n399);
    nand g340(n1784 ,n1511 ,n1405);
    nor g341(n272 ,n126 ,n230);
    nand g342(n1687 ,n36[1] ,n1110);
    nand g343(n933 ,n56[0] ,n476);
    nand g344(n987 ,n4[4] ,n712);
    nand g345(n1172 ,n670 ,n607);
    nand g346(n1374 ,n172 ,n1107);
    nand g347(n687 ,n27[0] ,n486);
    or g348(n517 ,n138 ,n369);
    nand g349(n919 ,n33[6] ,n404);
    nand g350(n561 ,n20[0] ,n405);
    nand g351(n1525 ,n32[0] ,n1101);
    nor g352(n722 ,n111 ,n360);
    or g353(n346 ,n37[3] ,n262);
    nand g354(n1070 ,n4[5] ,n706);
    not g355(n176 ,n177);
    nand g356(n1364 ,n178 ,n1104);
    nand g357(n945 ,n55[2] ,n416);
    nand g358(n674 ,n26[1] ,n393);
    nand g359(n657 ,n41[1] ,n372);
    nand g360(n574 ,n51[3] ,n386);
    nand g361(n1617 ,n1071 ,n604);
    or g362(n1324 ,n160 ,n1110);
    xor g363(n1946 ,n57[4] ,n72);
    nor g364(n294 ,n196 ,n282);
    nand g365(n729 ,n20[5] ,n405);
    nand g366(n1910 ,n1298 ,n1902);
    or g367(n1302 ,n179 ,n1095);
    nand g368(n1748 ,n1465 ,n1373);
    nor g369(n721 ,n111 ,n365);
    nor g370(n1320 ,n1200 ,n1118);
    dff g371(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1537), .Q(n56[5]));
    nand g372(n465 ,n6[4] ,n310);
    nand g373(n1468 ,n24[7] ,n1099);
    nand g374(n882 ,n47[7] ,n417);
    nor g375(n1319 ,n1167 ,n1166);
    or g376(n367 ,n194 ,n353);
    nand g377(n803 ,n46[1] ,n485);
    nand g378(n92 ,n59[1] ,n59[0]);
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1842), .Q(n59[3]));
    nand g380(n86 ,n57[1] ,n57[0]);
    nand g381(n1133 ,n778 ,n598);
    nand g382(n1593 ,n1005 ,n543);
    dff g383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n442), .Q(n17[3]));
    nand g384(n1160 ,n667 ,n873);
    nor g385(n193 ,n130 ,n15);
    nand g386(n1735 ,n1452 ,n1424);
    nor g387(n710 ,n157 ,n427);
    nor g388(n716 ,n186 ,n427);
    nand g389(n1080 ,n38[0] ,n703);
    nand g390(n673 ,n53[6] ,n370);
    or g391(n1392 ,n181 ,n1108);
    nand g392(n296 ,n172 ,n244);
    nand g393(n656 ,n27[3] ,n486);
    not g394(n426 ,n425);
    or g395(n1270 ,n156 ,n1105);
    not g396(n1697 ,n1684);
    nand g397(n752 ,n44[3] ,n398);
    buf g398(n10[5], n7[7]);
    nand g399(n1250 ,n907 ,n734);
    nor g400(n280 ,n118 ,n234);
    nand g401(n1908 ,n1327 ,n1905);
    nand g402(n550 ,n54[1] ,n392);
    nand g403(n445 ,n1953 ,n315);
    nand g404(n898 ,n50[3] ,n412);
    nor g405(n168 ,n123 ,n40[1]);
    dff g406(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1729), .Q(n27[5]));
    nand g407(n1717 ,n1343 ,n1339);
    nor g408(n248 ,n184 ,n230);
    nand g409(n1703 ,n1296 ,n1294);
    or g410(n1706 ,n1174 ,n1321);
    dff g411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1809), .Q(n35[5]));
    nor g412(n1340 ,n1162 ,n1216);
    nand g413(n867 ,n50[7] ,n412);
    nand g414(n1747 ,n1464 ,n1372);
    nand g415(n100 ,n58[1] ,n58[0]);
    dff g416(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1732), .Q(n27[2]));
    or g417(n1331 ,n1195 ,n1138);
    nor g418(n1303 ,n1140 ,n1132);
    dff g419(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1849), .Q(n36[3]));
    dff g420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1604), .Q(n49[3]));
    nand g421(n1715 ,n1348 ,n1337);
    buf g422(n9[0], 1'b0);
    nand g423(n567 ,n55[2] ,n374);
    nand g424(n538 ,n55[5] ,n374);
    nand g425(n959 ,n497 ,n519);
    nand g426(n326 ,n59[3] ,n252);
    nand g427(n1223 ,n628 ,n545);
    nand g428(n1737 ,n1454 ,n1364);
    nand g429(n566 ,n60[2] ,n420);
    nand g430(n1164 ,n860 ,n859);
    nand g431(n921 ,n28[1] ,n487);
    nand g432(n757 ,n22[4] ,n409);
    not g433(n125 ,n5[1]);
    nand g434(n1367 ,n180 ,n1104);
    nand g435(n1774 ,n1492 ,n1259);
    nand g436(n1835 ,n1658 ,n1305);
    nand g437(n1444 ,n27[7] ,n1091);
    nand g438(n1028 ,n4[5] ,n705);
    nand g439(n731 ,n464 ,n492);
    nand g440(n698 ,n24[6] ,n410);
    nor g441(n442 ,n272 ,n306);
    nand g442(n1075 ,n4[4] ,n714);
    nand g443(n268 ,n40[1] ,n225);
    nand g444(n1793 ,n1520 ,n1412);
    dff g445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1149), .Q(n16));
    dff g446(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n740), .Q(n18[1]));
    nand g447(n957 ,n512 ,n509);
    nand g448(n1368 ,n172 ,n1104);
    or g449(n1886 ,n1223 ,n1870);
    nand g450(n1537 ,n1028 ,n690);
    nand g451(n971 ,n4[6] ,n715);
    nor g452(n408 ,n237 ,n311);
    dff g453(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1623), .Q(n46[5]));
    nand g454(n1366 ,n174 ,n1104);
    nand g455(n212 ,n132 ,n198);
    nand g456(n1258 ,n155 ,n1090);
    nand g457(n1848 ,n1685 ,n1697);
    or g458(n231 ,n116 ,n200);
    nand g459(n591 ,n51[7] ,n401);
    nand g460(n1020 ,n4[6] ,n719);
    nand g461(n534 ,n27[1] ,n486);
    dff g462(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1830), .Q(n28[0]));
    nand g463(n972 ,n4[5] ,n715);
    nand g464(n573 ,n21[1] ,n406);
    nor g465(n1341 ,n1218 ,n1217);
    nand g466(n785 ,n30[7] ,n399);
    nand g467(n654 ,n53[4] ,n370);
    dff g468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n668), .Q(n39[0]));
    or g469(n1407 ,n177 ,n1109);
    nand g470(n1200 ,n866 ,n591);
    nand g471(n1095 ,n421 ,n723);
    not g472(n172 ,n173);
    or g473(n1428 ,n183 ,n1108);
    nand g474(n1811 ,n1498 ,n1397);
    nor g475(n199 ,n114 ,n58[3]);
    nand g476(n962 ,n493 ,n521);
    nand g477(n1536 ,n1027 ,n697);
    nand g478(n1175 ,n741 ,n874);
    nand g479(n1257 ,n155 ,n1100);
    nand g480(n343 ,n276 ,n241);
    nand g481(n1219 ,n834 ,n852);
    or g482(n1395 ,n179 ,n1087);
    nor g483(n425 ,n111 ,n294);
    nand g484(n386 ,n255 ,n318);
    nand g485(n587 ,n49[4] ,n388);
    nand g486(n1045 ,n4[1] ,n714);
    nand g487(n1664 ,n999 ,n650);
    nand g488(n1213 ,n858 ,n877);
    or g489(n293 ,n254 ,n215);
    nand g490(n1807 ,n1494 ,n1429);
    nand g491(n1759 ,n1476 ,n1427);
    nand g492(n449 ,n16 ,n349);
    dff g493(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1884), .Q(n60[3]));
    not g494(n373 ,n374);
    nand g495(n844 ,n23[2] ,n413);
    nor g496(n136 ,n111 ,n48[0]);
    dff g497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1780), .Q(n34[2]));
    nand g498(n1709 ,n1329 ,n1317);
    nand g499(n1494 ,n35[7] ,n1087);
    nand g500(n1801 ,n1528 ,n1418);
    nand g501(n1645 ,n987 ,n694);
    dff g502(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1776), .Q(n34[6]));
    nand g503(n537 ,n55[7] ,n374);
    dff g504(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1578), .Q(n52[7]));
    nor g505(n169 ,n121 ,n111);
    nand g506(n1671 ,n20[6] ,n1105);
    not g507(n81 ,n80);
    or g508(n496 ,n145 ,n383);
    dff g509(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1761), .Q(n23[5]));
    nor g510(n396 ,n312 ,n348);
    nand g511(n319 ,n112 ,n249);
    not g512(n312 ,n313);
    or g513(n1399 ,n171 ,n1102);
    dff g514(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n951), .Q(n46[0]));
    nand g515(n1497 ,n35[4] ,n1087);
    nand g516(n771 ,n48[5] ,n483);
    dff g517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1648), .Q(n43[1]));
    nand g518(n1022 ,n4[4] ,n719);
    or g519(n1401 ,n181 ,n1087);
    nand g520(n1191 ,n463 ,n676);
    nand g521(n1948 ,n65 ,n64);
    dff g522(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1605), .Q(n49[2]));
    nand g523(n1556 ,n1026 ,n666);
    dff g524(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1812), .Q(n35[2]));
    nand g525(n1055 ,n4[5] ,n708);
    nand g526(n1533 ,n31[0] ,n1098);
    nand g527(n71 ,n57[2] ,n67);
    dff g528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1536), .Q(n56[6]));
    nand g529(n1116 ,n578 ,n749);
    nand g530(n631 ,n43[6] ,n376);
    nand g531(n1719 ,n1534 ,n1434);
    dff g532(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1801), .Q(n31[5]));
    nand g533(n636 ,n21[2] ,n406);
    nand g534(n1771 ,n1489 ,n1391);
    nand g535(n1033 ,n4[7] ,n705);
    nand g536(n613 ,n60[0] ,n420);
    nand g537(n1504 ,n34[5] ,n1102);
    nand g538(n557 ,n51[0] ,n401);
    nand g539(n1512 ,n33[5] ,n1109);
    or g540(n1881 ,n1179 ,n1866);
    not g541(n89 ,n88);
    nand g542(n1580 ,n1021 ,n562);
    dff g543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1741), .Q(n26[1]));
    or g544(n1404 ,n173 ,n1102);
    nand g545(n681 ,n55[6] ,n374);
    xnor g546(n1941 ,n57[3] ,n88);
    nand g547(n1787 ,n1514 ,n1408);
    dff g548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1859), .Q(n20[6]));
    nand g549(n832 ,n42[5] ,n475);
    not g550(n1087 ,n1088);
    nand g551(n187 ,n59[1] ,n115);
    nand g552(n1736 ,n1453 ,n1363);
    nand g553(n1040 ,n4[7] ,n714);
    nand g554(n1574 ,n1044 ,n644);
    dff g555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1647), .Q(n43[2]));
    nand g556(n1205 ,n566 ,n596);
    nand g557(n559 ,n52[7] ,n384);
    dff g558(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1634), .Q(n45[1]));
    nor g559(n266 ,n19[0] ,n228);
    nand g560(n1508 ,n34[1] ,n1102);
    dff g561(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1594), .Q(n50[6]));
    nor g562(n107 ,n18[1] ,n18[0]);
    nand g563(n204 ,n18[0] ,n18[2]);
    nand g564(n977 ,n4[7] ,n717);
    nand g565(n1745 ,n1462 ,n1370);
    nand g566(n1823 ,n1564 ,n1281);
    nand g567(n691 ,n56[2] ,n378);
    nand g568(n1084 ,n1926 ,n725);
    nor g569(n156 ,n111 ,n3);
    nand g570(n963 ,n4[7] ,n716);
    nand g571(n1890 ,n899 ,n1865);
    nand g572(n853 ,n53[3] ,n408);
    dff g573(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1759), .Q(n23[7]));
    nand g574(n887 ,n33[1] ,n404);
    not g575(n101 ,n100);
    nand g576(n1479 ,n23[4] ,n1089);
    nand g577(n1749 ,n1466 ,n1374);
    not g578(n477 ,n478);
    dff g579(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1822), .Q(n29[0]));
    nand g580(n489 ,n59[3] ,n354);
    nand g581(n960 ,n494 ,n520);
    nand g582(n470 ,n337 ,n329);
    nand g583(n1245 ,n743 ,n687);
    nor g584(n413 ,n233 ,n347);
    nand g585(n1546 ,n1036 ,n582);
    or g586(n1418 ,n179 ,n1098);
    dff g587(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1857), .Q(n20[4]));
    nor g588(n290 ,n17[1] ,n253);
    dff g589(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1664), .Q(n41[6]));
    dff g590(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1643), .Q(n43[6]));
    xor g591(n1949 ,n36[3] ,n63);
    not g592(n479 ,n480);
    nand g593(n427 ,n113 ,n354);
    nand g594(n271 ,n226 ,n230);
    nand g595(n1469 ,n24[6] ,n1099);
    nor g596(n164 ,n37[2] ,n40[0]);
    nand g597(n815 ,n44[3] ,n478);
    nand g598(n451 ,n57[0] ,n316);
    not g599(n178 ,n179);
    nor g600(n1288 ,n1114 ,n1113);
    nand g601(n868 ,n42[7] ,n403);
    nor g602(n1925 ,n97 ,n95);
    nor g603(n1904 ,n1237 ,n1879);
    dff g604(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1739), .Q(n26[3]));
    nand g605(n1643 ,n985 ,n631);
    nand g606(n1618 ,n1072 ,n605);
    not g607(n105 ,n104);
    nor g608(n1861 ,n1112 ,n1701);
    nand g609(n1768 ,n1695 ,n1388);
    buf g610(n10[1], 1'b0);
    or g611(n358 ,n295 ,n308);
    nand g612(n1147 ,n822 ,n830);
    nand g613(n1583 ,n1025 ,n614);
    or g614(n505 ,n151 ,n377);
    nand g615(n1450 ,n27[2] ,n1091);
    nand g616(n612 ,n20[3] ,n405);
    nor g617(n152 ,n111 ,n54[0]);
    not g618(n421 ,n422);
    dff g619(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n356), .Q(n15));
    dff g620(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1085), .Q(n12));
    nand g621(n1529 ,n31[4] ,n1098);
    nand g622(n840 ,n53[4] ,n408);
    nand g623(n826 ,n449 ,n455);
    dff g624(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n958), .Q(n48[0]));
    nand g625(n1653 ,n992 ,n831);
    nand g626(n388 ,n258 ,n318);
    or g627(n1878 ,n1212 ,n1715);
    nand g628(n330 ,n1941 ,n249);
    nand g629(n1073 ,n4[2] ,n706);
    dff g630(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1788), .Q(n33[2]));
    nand g631(n1606 ,n1059 ,n592);
    dff g632(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1493), .Q(n36[4]));
    nand g633(n532 ,n50[3] ,n380);
    nand g634(n1441 ,n30[2] ,n1094);
    nand g635(n615 ,n24[3] ,n410);
    or g636(n61 ,n36[1] ,n36[0]);
    or g637(n1393 ,n173 ,n1108);
    nand g638(n390 ,n257 ,n314);
    or g639(n1432 ,n183 ,n1101);
    dff g640(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1829), .Q(n28[1]));
    nand g641(n1000 ,n4[5] ,n709);
    nand g642(n454 ,n341 ,n333);
    nand g643(n777 ,n48[1] ,n483);
    nand g644(n765 ,n34[5] ,n411);
    nand g645(n1554 ,n29[3] ,n1097);
    nand g646(n1483 ,n155 ,n1093);
    nand g647(n540 ,n50[5] ,n380);
    nand g648(n444 ,n18[3] ,n345);
    nand g649(n804 ,n44[1] ,n398);
    nand g650(n585 ,n49[6] ,n388);
    or g651(n257 ,n111 ,n208);
    dff g652(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1856), .Q(n20[3]));
    nand g653(n1743 ,n1460 ,n1425);
    nand g654(n1086 ,n4[3] ,n718);
    nand g655(n838 ,n42[1] ,n475);
    nand g656(n1836 ,n1660 ,n1306);
    dff g657(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1876), .Q(n38[3]));
    nand g658(n1451 ,n27[0] ,n1091);
    nand g659(n108 ,n18[1] ,n18[0]);
    or g660(n1421 ,n181 ,n1098);
    dff g661(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1779), .Q(n34[3]));
    nand g662(n1841 ,n323 ,n1690);
    or g663(n1389 ,n179 ,n1108);
    or g664(n1321 ,n1142 ,n1171);
    nand g665(n697 ,n56[6] ,n378);
    dff g666(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n343), .Q(n11));
    nand g667(n774 ,n48[4] ,n483);
    nand g668(n617 ,n45[6] ,n382);
    nand g669(n994 ,n4[4] ,n710);
    nand g670(n437 ,n327 ,n319);
    nand g671(n238 ,n58[2] ,n199);
    nand g672(n1770 ,n1488 ,n1390);
    nand g673(n98 ,n37[2] ,n97);
    nand g674(n530 ,n26[5] ,n393);
    nor g675(n137 ,n111 ,n45[0]);
    nand g676(n1481 ,n23[2] ,n1089);
    nand g677(n680 ,n49[5] ,n388);
    nand g678(n551 ,n53[7] ,n370);
    nand g679(n1072 ,n4[3] ,n706);
    nand g680(n1507 ,n34[2] ,n1102);
    dff g681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1811), .Q(n35[3]));
    nand g682(n1520 ,n32[5] ,n1101);
    nand g683(n488 ,n59[3] ,n320);
    nand g684(n1596 ,n1008 ,n579);
    or g685(n359 ,n297 ,n285);
    nor g686(n713 ,n187 ,n488);
    or g687(n1419 ,n177 ,n1098);
    or g688(n501 ,n149 ,n373);
    dff g689(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1802), .Q(n31[4]));
    nand g690(n916 ,n44[6] ,n398);
    not g691(n383 ,n384);
    nand g692(n589 ,n49[3] ,n388);
    or g693(n232 ,n128 ,n184);
    nand g694(n672 ,n25[1] ,n415);
    dff g695(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1612), .Q(n48[2]));
    nand g696(n1555 ,n1014 ,n542);
    nand g697(n1044 ,n4[2] ,n714);
    or g698(n1269 ,n156 ,n1095);
    nor g699(n144 ,n111 ,n44[0]);
    or g700(n1268 ,n156 ,n1096);
    dff g701(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1826), .Q(n28[4]));
    nand g702(n1695 ,n22[6] ,n1108);
    or g703(n241 ,n188 ,n232);
    nand g704(n982 ,n4[2] ,n717);
    dff g705(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1770), .Q(n22[4]));
    nand g706(n739 ,n35[5] ,n481);
    nand g707(n1726 ,n1443 ,n1483);
    or g708(n314 ,n111 ,n242);
    nand g709(n1764 ,n1481 ,n1386);
    nand g710(n611 ,n25[3] ,n415);
    nand g711(n1452 ,n26[7] ,n1103);
    nand g712(n1666 ,n1000 ,n652);
    or g713(n1414 ,n175 ,n1101);
    nand g714(n1601 ,n1054 ,n585);
    nand g715(n1252 ,n530 ,n733);
    nor g716(n1336 ,n1122 ,n1207);
    nand g717(n1621 ,n963 ,n789);
    nor g718(n324 ,n119 ,n259);
    nand g719(n336 ,n1947 ,n246);
    nand g720(n770 ,n29[4] ,n407);
    nand g721(n1818 ,n1552 ,n1276);
    or g722(n1400 ,n179 ,n1102);
    nand g723(n670 ,n26[7] ,n393);
    dff g724(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1763), .Q(n23[3]));
    nand g725(n872 ,n28[5] ,n487);
    nand g726(n927 ,n60[5] ,n396);
    nand g727(n1676 ,n20[2] ,n1105);
    nand g728(n302 ,n253 ,n247);
    nand g729(n984 ,n4[7] ,n712);
    nand g730(n1113 ,n552 ,n872);
    nor g731(n418 ,n236 ,n311);
    nand g732(n1665 ,n21[0] ,n1095);
    nand g733(n1551 ,n1039 ,n536);
    nand g734(n1502 ,n34[7] ,n1102);
    nand g735(n1605 ,n1058 ,n590);
    dff g736(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1843), .Q(n36[0]));
    or g737(n1287 ,n181 ,n1096);
    nand g738(n788 ,n31[3] ,n402);
    nand g739(n746 ,n47[6] ,n417);
    nand g740(n179 ,n39[4] ,n1);
    xor g741(n1938 ,n19[1] ,n19[0]);
    dff g742(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1806), .Q(n31[0]));
    dff g743(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1838), .Q(n21[0]));
    nand g744(n1236 ,n931 ,n930);
    nor g745(n139 ,n111 ,n47[0]);
    nand g746(n1161 ,n857 ,n674);
    or g747(n311 ,n58[0] ,n247);
    nand g748(n935 ,n34[0] ,n411);
    nand g749(n1487 ,n22[5] ,n1108);
    nand g750(n1377 ,n176 ,n1100);
    nand g751(n65 ,n36[2] ,n61);
    nand g752(n1154 ,n851 ,n854);
    nand g753(n1725 ,n1442 ,n1356);
    nand g754(n1752 ,n1469 ,n1375);
    nand g755(n942 ,n21[6] ,n406);
    dff g756(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1791), .Q(n32[7]));
    nand g757(n334 ,n1945 ,n248);
    nor g758(n1907 ,n1225 ,n1886);
    nor g759(n1343 ,n1229 ,n1220);
    not g760(n1698 ,n1686);
    or g761(n255 ,n111 ,n211);
    nand g762(n1834 ,n1656 ,n1304);
    dff g763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n331), .Q(n19[1]));
    nor g764(n242 ,n59[0] ,n217);
    dff g765(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1744), .Q(n25[6]));
    nor g766(n288 ,n184 ,n268);
    nand g767(n584 ,n49[7] ,n388);
    dff g768(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1858), .Q(n20[5]));
    nand g769(n793 ,n46[4] ,n480);
    nand g770(n662 ,n25[0] ,n415);
    nor g771(n397 ,n219 ,n311);
    buf g772(n8[6], 1'b0);
    nand g773(n845 ,n35[2] ,n481);
    nand g774(n1037 ,n4[3] ,n711);
    nand g775(n545 ,n41[1] ,n400);
    dff g776(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1787), .Q(n33[3]));
    nand g777(n541 ,n41[7] ,n400);
    nand g778(n1608 ,n1061 ,n760);
    dff g779(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1789), .Q(n33[1]));
    dff g780(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1728), .Q(n27[6]));
    dff g781(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n731), .Q(n57[1]));
    nand g782(n1234 ,n763 ,n594);
    nor g783(n142 ,n111 ,n41[0]);
    nand g784(n1585 ,n1024 ,n570);
    dff g785(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n962), .Q(n51[0]));
    nand g786(n647 ,n45[2] ,n382);
    nand g787(n506 ,n153 ,n375);
    buf g788(n9[6], 1'b0);
    nand g789(n1729 ,n1446 ,n1358);
    nand g790(n653 ,n41[4] ,n372);
    nand g791(n624 ,n45[1] ,n382);
    nand g792(n883 ,n32[7] ,n414);
    nand g793(n1575 ,n1045 ,n556);
    nand g794(n217 ,n113 ,n159);
    nand g795(n854 ,n30[2] ,n399);
    not g796(n129 ,n58[3]);
    nand g797(n979 ,n4[5] ,n717);
    nand g798(n1917 ,n1303 ,n1897);
    or g799(n303 ,n37[0] ,n245);
    nand g800(n1145 ,n637 ,n892);
    nand g801(n642 ,n43[1] ,n419);
    nand g802(n926 ,n23[5] ,n413);
    nand g803(n1387 ,n172 ,n1090);
    nor g804(n1865 ,n1187 ,n1709);
    nand g805(n808 ,n22[3] ,n409);
    nand g806(n1386 ,n180 ,n1090);
    nand g807(n1678 ,n20[0] ,n1105);
    nand g808(n544 ,n26[4] ,n393);
    nand g809(n533 ,n56[4] ,n378);
    nand g810(n1042 ,n4[5] ,n714);
    or g811(n1429 ,n183 ,n1087);
    nand g812(n813 ,n35[7] ,n481);
    nor g813(n706 ,n185 ,n428);
    nand g814(n1115 ,n696 ,n560);
    nand g815(n968 ,n4[2] ,n716);
    or g816(n1390 ,n177 ,n1108);
    nand g817(n577 ,n50[6] ,n380);
    nor g818(n1931 ,n105 ,n103);
    nand g819(n1373 ,n180 ,n1107);
    nand g820(n1668 ,n20[7] ,n1105);
    nand g821(n1165 ,n1936 ,n704);
    nand g822(n1076 ,n496 ,n522);
    nand g823(n940 ,n444 ,n445);
    nand g824(n1720 ,n1437 ,n1351);
    dff g825(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n324), .Q(n7[3]));
    nand g826(n1786 ,n1513 ,n1407);
    dff g827(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1657), .Q(n42[3]));
    nand g828(n1911 ,n1316 ,n1899);
    nand g829(n1199 ,n813 ,n846);
    nand g830(n1140 ,n806 ,n802);
    nand g831(n1506 ,n34[3] ,n1102);
    nand g832(n1206 ,n745 ,n640);
    nor g833(n1901 ,n1240 ,n1891);
    nand g834(n1059 ,n4[1] ,n708);
    dff g835(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n728), .Q(n57[0]));
    nand g836(n852 ,n42[1] ,n403);
    nand g837(n1380 ,n172 ,n1100);
    or g838(n1388 ,n171 ,n1108);
    nand g839(n1853 ,n1933 ,n1485);
    dff g840(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1620), .Q(n47[1]));
    dff g841(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1631), .Q(n45[4]));
    nand g842(n875 ,n31[7] ,n402);
    dff g843(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1736), .Q(n26[6]));
    or g844(n1411 ,n171 ,n1101);
    nand g845(n219 ,n129 ,n192);
    nand g846(n993 ,n4[5] ,n710);
    not g847(n119 ,n57[4]);
    nand g848(n1142 ,n684 ,n867);
    nand g849(n1826 ,n1571 ,n1284);
    nor g850(n216 ,n40[0] ,n184);
    nor g851(n393 ,n231 ,n346);
    nand g852(n620 ,n54[3] ,n392);
    nand g853(n1547 ,n1037 ,n539);
    nand g854(n278 ,n1942 ,n215);
    or g855(n1335 ,n1205 ,n1204);
    nor g856(n403 ,n221 ,n344);
    nand g857(n986 ,n4[5] ,n712);
    buf g858(n9[3], 1'b0);
    dff g859(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1078), .Q(n54[0]));
    not g860(n111 ,n1);
    nand g861(n864 ,n34[7] ,n411);
    nand g862(n1682 ,n335 ,n1165);
    nand g863(n768 ,n48[7] ,n483);
    nand g864(n435 ,n37[1] ,n310);
    nand g865(n1568 ,n28[5] ,n1096);
    or g866(n1274 ,n171 ,n1097);
    nand g867(n614 ,n52[3] ,n384);
    nand g868(n1799 ,n1526 ,n1433);
    nor g869(n299 ,n177 ,n243);
    nand g870(n203 ,n19[0] ,n38[2]);
    dff g871(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1769), .Q(n20[7]));
    nand g872(n1539 ,n1029 ,n686);
    nor g873(n246 ,n40[0] ,n234);
    nor g874(n1107 ,n422 ,n722);
    nand g875(n1079 ,n501 ,n702);
    nand g876(n835 ,n31[5] ,n402);
    or g877(n1879 ,n1236 ,n1875);
    nand g878(n1765 ,n1482 ,n1387);
    nand g879(n954 ,n500 ,n516);
    nand g880(n676 ,n24[7] ,n410);
    nand g881(n236 ,n58[3] ,n163);
    nand g882(n483 ,n257 ,n352);
    nand g883(n569 ,n43[6] ,n419);
    nand g884(n1212 ,n917 ,n626);
    nand g885(n1221 ,n825 ,n819);
    nand g886(n1385 ,n174 ,n1090);
    nand g887(n1592 ,n1052 ,n576);
    nor g888(n1860 ,n1247 ,n1700);
    nand g889(n80 ,n36[1] ,n36[0]);
    nand g890(n542 ,n54[6] ,n392);
    dff g891(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1635), .Q(n44[7]));
    dff g892(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1565), .Q(n53[7]));
    nand g893(n1680 ,n460 ,n1084);
    nand g894(n1509 ,n34[0] ,n1102);
    nand g895(n863 ,n340 ,n438);
    nand g896(n740 ,n473 ,n448);
    or g897(n1354 ,n175 ,n1094);
    nand g898(n661 ,n26[0] ,n393);
    dff g899(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n730), .Q(n57[2]));
    nand g900(n889 ,n46[7] ,n485);
    nand g901(n1809 ,n1496 ,n1395);
    nand g902(n1144 ,n918 ,n927);
    nand g903(n980 ,n4[4] ,n717);
    nand g904(n1639 ,n981 ,n815);
    nand g905(n1534 ,n30[7] ,n1094);
    nand g906(n693 ,n43[3] ,n376);
    nand g907(n1892 ,n845 ,n1864);
    nand g908(n1637 ,n979 ,n812);
    nand g909(n1869 ,n1844 ,n1851);
    nor g910(n414 ,n213 ,n350);
    or g911(n1314 ,n181 ,n1105);
    nand g912(n811 ,n44[6] ,n478);
    not g913(n1937 ,n84);
    dff g914(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1599), .Q(n50[1]));
    or g915(n1309 ,n183 ,n1105);
    dff g916(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1773), .Q(n22[1]));
    nand g917(n623 ,n41[4] ,n400);
    nand g918(n747 ,n49[2] ,n418);
    or g919(n1285 ,n175 ,n1096);
    nand g920(n1884 ,n1336 ,n1874);
    dff g921(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1762), .Q(n23[4]));
    nand g922(n1466 ,n25[1] ,n1106);
    nand g923(n734 ,n53[2] ,n408);
    dff g924(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1547), .Q(n55[3]));
    not g925(n377 ,n378);
    nand g926(n859 ,n28[7] ,n487);
    nand g927(n1204 ,n900 ,n762);
    dff g928(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1815), .Q(n29[7]));
    nand g929(n1150 ,n828 ,n833);
    nand g930(n828 ,n34[2] ,n411);
    not g931(n138 ,n53[0]);
    nor g932(n1329 ,n1180 ,n1169);
    nand g933(n738 ,n52[3] ,n484);
    or g934(n1259 ,n156 ,n1108);
    nand g935(n1423 ,n182 ,n1092);
    nand g936(n728 ,n357 ,n451);
    nand g937(n885 ,n56[6] ,n476);
    nand g938(n917 ,n48[2] ,n395);
    or g939(n1108 ,n429 ,n724);
    buf g940(n8[3], 1'b0);
    dff g941(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1764), .Q(n23[2]));
    nand g942(n1824 ,n1566 ,n1282);
    nand g943(n925 ,n53[0] ,n408);
    nor g944(n1334 ,n1201 ,n1199);
    nand g945(n1808 ,n1495 ,n1394);
    nor g946(n1298 ,n1143 ,n1141);
    nand g947(n1528 ,n31[5] ,n1098);
    nand g948(n1192 ,n840 ,n888);
    or g949(n361 ,n299 ,n283);
    nand g950(n671 ,n60[3] ,n420);
    nand g951(n1046 ,n4[7] ,n713);
    dff g952(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1755), .Q(n24[3]));
    nand g953(n1578 ,n1019 ,n559);
    nand g954(n237 ,n58[3] ,n192);
    nor g955(n1342 ,n1147 ,n1219);
    xnor g956(n1933 ,n38[3] ,n106);
    nand g957(n1591 ,n1051 ,n563);
    not g958(n424 ,n423);
    nand g959(n568 ,n52[2] ,n384);
    nand g960(n549 ,n54[2] ,n392);
    nand g961(n1163 ,n1937 ,n704);
    nand g962(n619 ,n45[5] ,n382);
    dff g963(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1804), .Q(n31[2]));
    nand g964(n578 ,n25[4] ,n415);
    dff g965(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1850), .Q(n20[0]));
    nor g966(n407 ,n214 ,n351);
    nand g967(n1124 ,n466 ,n755);
    nand g968(n1821 ,n1559 ,n1279);
    nand g969(n1629 ,n971 ,n617);
    not g970(n492 ,n470);
    buf g971(n726 ,n248);
    or g972(n1381 ,n177 ,n1102);
    nor g973(n165 ,n111 ,n40[1]);
    nand g974(n606 ,n47[2] ,n390);
    nand g975(n1788 ,n1515 ,n1409);
    nor g976(n146 ,n111 ,n43[0]);
    nand g977(n1478 ,n23[5] ,n1089);
    nand g978(n981 ,n4[3] ,n717);
    or g979(n1356 ,n173 ,n1094);
    not g980(n202 ,n201);
    nand g981(n1758 ,n1475 ,n1257);
    nand g982(n1705 ,n1320 ,n1319);
    nand g983(n976 ,n4[1] ,n715);
    dff g984(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1553), .Q(n54[7]));
    dff g985(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1778), .Q(n34[4]));
    or g986(n1261 ,n156 ,n1102);
    not g987(n117 ,n19[0]);
    nor g988(n297 ,n175 ,n243);
    not g989(n262 ,n261);
    nand g990(n985 ,n4[6] ,n712);
    nand g991(n1955 ,n74 ,n75);
    nand g992(n776 ,n48[2] ,n483);
    nand g993(n807 ,n54[4] ,n394);
    nand g994(n1220 ,n914 ,n913);
    dff g995(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1641), .Q(n44[1]));
    nand g996(n1849 ,n1683 ,n1696);
    nand g997(n1255 ,n155 ,n1104);
    nand g998(n1677 ,n20[1] ,n1105);
    nor g999(n406 ,n214 ,n347);
    nor g1000(n1899 ,n1156 ,n1892);
    nand g1001(n1816 ,n1548 ,n1274);
    nand g1002(n1209 ,n904 ,n942);
    dff g1003(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1603), .Q(n49[4]));
    nand g1004(n784 ,n28[0] ,n487);
    nand g1005(n1237 ,n557 ,n932);
    nor g1006(n1718 ,n1346 ,n1345);
    nand g1007(n1773 ,n1491 ,n1393);
    nor g1008(n711 ,n185 ,n488);
    nand g1009(n1243 ,n944 ,n893);
    dff g1010(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1638), .Q(n44[4]));
    nand g1011(n1649 ,n21[7] ,n1095);
    nand g1012(n1803 ,n1530 ,n1420);
    nand g1013(n727 ,n456 ,n491);
    dff g1014(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1808), .Q(n35[6]));
    nand g1015(n1194 ,n773 ,n901);
    not g1016(n133 ,n59[1]);
    dff g1017(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1754), .Q(n24[4]));
    nand g1018(n1054 ,n4[6] ,n708);
    not g1019(n482 ,n483);
    dff g1020(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1819), .Q(n29[3]));
    not g1021(n112 ,n59[0]);
    nand g1022(n1859 ,n1671 ,n1310);
    nand g1023(n1031 ,n4[1] ,n705);
    dff g1024(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1556), .Q(n54[5]));
    nand g1025(n1383 ,n178 ,n1090);
    nand g1026(n357 ,n161 ,n293);
    nand g1027(n996 ,n4[2] ,n710);
    nor g1028(n717 ,n187 ,n427);
    nor g1029(n1871 ,n1233 ,n1717);
    or g1030(n1430 ,n183 ,n1102);
    nand g1031(n1424 ,n182 ,n1104);
    buf g1032(n8[7], 1'b0);
    nand g1033(n1008 ,n4[4] ,n718);
    nand g1034(n855 ,n42[6] ,n403);
    nand g1035(n823 ,n22[2] ,n409);
    dff g1036(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1666), .Q(n41[5]));
    nand g1037(n1673 ,n20[5] ,n1105);
    dff g1038(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1749), .Q(n25[1]));
    dff g1039(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1810), .Q(n35[4]));
    nand g1040(n458 ,n6[2] ,n310);
    nand g1041(n529 ,n446 ,n368);
    nor g1042(n395 ,n238 ,n344);
    nor g1043(n1874 ,n1714 ,n1713);
    nand g1044(n1378 ,n174 ,n1100);
    dff g1045(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1551), .Q(n55[1]));
    dff g1046(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n362), .Q(n39[4]));
    nand g1047(n754 ,n48[7] ,n395);
    nand g1048(n850 ,n31[2] ,n402);
    nand g1049(n601 ,n47[6] ,n390);
    nand g1050(n448 ,n1951 ,n315);
    nor g1051(n287 ,n57[4] ,n259);
    nand g1052(n1628 ,n970 ,n616);
    nand g1053(n1129 ,n897 ,n764);
    nand g1054(n973 ,n4[4] ,n715);
    nand g1055(n1482 ,n23[1] ,n1089);
    nand g1056(n339 ,n1948 ,n246);
    dff g1057(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1588), .Q(n51[5]));
    dff g1058(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n953), .Q(n44[0]));
    nand g1059(n227 ,n1955 ,n168);
    dff g1060(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1659), .Q(n42[2]));
    nand g1061(n1198 ,n781 ,n610);
    nor g1062(n1317 ,n1161 ,n1158);
    nor g1063(n411 ,n231 ,n350);
    or g1064(n1281 ,n183 ,n1096);
    dff g1065(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1751), .Q(n24[7]));
    nand g1066(n906 ,n56[2] ,n476);
    not g1067(n490 ,n454);
    nand g1068(n897 ,n56[3] ,n476);
    or g1069(n1109 ,n423 ,n722);
    dff g1070(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1591), .Q(n51[2]));
    nand g1071(n473 ,n18[1] ,n345);
    nand g1072(n732 ,n24[5] ,n410);
    nand g1073(n1741 ,n1458 ,n1368);
    nand g1074(n1806 ,n1533 ,n1264);
    nor g1075(n308 ,n179 ,n244);
    dff g1076(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1795), .Q(n32[3]));
    nand g1077(n1526 ,n31[7] ,n1098);
    dff g1078(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1636), .Q(n44[6]));
    dff g1079(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1616), .Q(n47[5]));
    nand g1080(n1586 ,n1046 ,n571);
    nand g1081(n1711 ,n1330 ,n1328);
    nor g1082(n338 ,n196 ,n279);
    dff g1083(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1608), .Q(n48[6]));
    or g1084(n493 ,n135 ,n385);
    nand g1085(n438 ,n36[4] ,n310);
    dff g1086(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n955), .Q(n43[0]));
    not g1087(n391 ,n392);
    nand g1088(n1135 ,n788 ,n783);
    nor g1089(n1905 ,n1189 ,n1882);
    nand g1090(n531 ,n55[6] ,n416);
    nand g1091(n745 ,n54[3] ,n394);
    or g1092(n1416 ,n173 ,n1101);
    nand g1093(n1858 ,n1673 ,n1311);
    nand g1094(n1139 ,n467 ,n656);
    not g1095(n381 ,n382);
    nand g1096(n1134 ,n779 ,n782);
    nand g1097(n1222 ,n1950 ,n704);
    nand g1098(n1015 ,n4[4] ,n720);
    nand g1099(n1228 ,n613 ,n803);
    or g1100(n1885 ,n1213 ,n1878);
    nand g1101(n1658 ,n21[3] ,n1095);
    nand g1102(n847 ,n53[7] ,n408);
    not g1103(n126 ,n5[3]);
    dff g1104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1672), .Q(n41[1]));
    nand g1105(n1893 ,n801 ,n1863);
    dff g1106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1765), .Q(n23[1]));
    nand g1107(n1833 ,n1652 ,n1302);
    nand g1108(n352 ,n1 ,n267);
    dff g1109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1585), .Q(n52[1]));
    nor g1110(n415 ,n213 ,n347);
    nand g1111(n1486 ,n22[7] ,n1108);
    or g1112(n1870 ,n1221 ,n1716);
    nand g1113(n102 ,n58[2] ,n101);
    nand g1114(n1006 ,n4[6] ,n718);
    nand g1115(n1027 ,n4[6] ,n705);
    nand g1116(n322 ,n59[1] ,n252);
    nand g1117(n1078 ,n518 ,n523);
    dff g1118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1916), .Q(n60[2]));
    nor g1119(n498 ,n136 ,n482);
    nor g1120(n705 ,n185 ,n489);
    dff g1121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n940), .Q(n18[3]));
    nand g1122(n1563 ,n1018 ,n550);
    nand g1123(n457 ,n58[0] ,n313);
    or g1124(n1413 ,n177 ,n1101);
    nand g1125(n1590 ,n1050 ,n574);
    nand g1126(n197 ,n18[1] ,n122);
    nand g1127(n1247 ,n739 ,n926);
    nand g1128(n799 ,n31[6] ,n402);
    nand g1129(n1577 ,n28[1] ,n1096);
    nand g1130(n1208 ,n796 ,n824);
    nand g1131(n824 ,n60[2] ,n396);
    nand g1132(n1538 ,n1032 ,n533);
    not g1133(n135 ,n51[0]);
    nand g1134(n1488 ,n22[4] ,n1108);
    nand g1135(n1216 ,n682 ,n747);
    or g1136(n1284 ,n177 ,n1096);
    or g1137(n500 ,n139 ,n389);
    not g1138(n243 ,n244);
    dff g1139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1758), .Q(n24[0]));
    nand g1140(n524 ,n36[4] ,n432);
    nand g1141(n818 ,n44[1] ,n478);
    nand g1142(n1011 ,n4[2] ,n718);
    not g1143(n349 ,n348);
    dff g1144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1775), .Q(n34[7]));
    nor g1145(n69 ,n57[2] ,n67);
    nand g1146(n755 ,n32[0] ,n414);
    nand g1147(n570 ,n52[1] ,n384);
    nand g1148(n890 ,n49[5] ,n418);
    dff g1149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n328), .Q(n7[2]));
    nand g1150(n663 ,n24[2] ,n410);
    nand g1151(n282 ,n38[3] ,n224);
    xnor g1152(n1932 ,n38[2] ,n104);
    buf g1153(n10[4], n7[7]);
    nand g1154(n190 ,n2 ,n128);
    nand g1155(n1518 ,n32[7] ,n1101);
    nor g1156(n161 ,n111 ,n57[0]);
    not g1157(n310 ,n309);
    nand g1158(n822 ,n48[1] ,n395);
    dff g1159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1820), .Q(n29[2]));
    nand g1160(n456 ,n57[3] ,n316);
    dff g1161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1880), .Q(n60[7]));
    dff g1162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1743), .Q(n25[7]));
    nand g1163(n860 ,n23[7] ,n413);
    nand g1164(n1226 ,n935 ,n939);
    nor g1165(n284 ,n36[4] ,n260);
    nand g1166(n1251 ,n742 ,n688);
    nand g1167(n1730 ,n1447 ,n1359);
    nor g1168(n1436 ,n111 ,n1080);
    nor g1169(n1864 ,n1153 ,n1704);
    nand g1170(n923 ,n34[1] ,n411);
    nor g1171(n209 ,n57[3] ,n162);
    nand g1172(n1894 ,n750 ,n1861);
    or g1173(n1431 ,n183 ,n1109);
    nor g1174(n275 ,n124 ,n230);
    nand g1175(n1186 ,n603 ,n903);
    dff g1176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n266), .Q(n19[0]));
    nand g1177(n743 ,n33[0] ,n404);
    dff g1178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1655), .Q(n42[4]));
    nand g1179(n1064 ,n4[3] ,n707);
    or g1180(n1311 ,n179 ,n1105);
    nand g1181(n802 ,n23[0] ,n413);
    nand g1182(n787 ,n49[0] ,n418);
    nand g1183(n1825 ,n1568 ,n1283);
    nand g1184(n1131 ,n588 ,n896);
    nor g1185(n1485 ,n703 ,n1088);
    nand g1186(n820 ,n48[4] ,n395);
    nand g1187(n741 ,n54[6] ,n394);
    nand g1188(n1527 ,n31[6] ,n1098);
    nand g1189(n1188 ,n683 ,n890);
    dff g1190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1575), .Q(n53[1]));
    nand g1191(n1224 ,n916 ,n664);
    dff g1192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n952), .Q(n56[0]));
    nand g1193(n1235 ,n661 ,n561);
    dff g1194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1155), .Q(n8[1]));
    nand g1195(n839 ,n29[2] ,n407);
    dff g1196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1855), .Q(n20[2]));
    nand g1197(n1007 ,n4[5] ,n718);
    nand g1198(n1600 ,n1053 ,n584);
    nand g1199(n1030 ,n4[2] ,n705);
    nand g1200(n1794 ,n1521 ,n1413);
    nand g1201(n1800 ,n1527 ,n1417);
    or g1202(n1278 ,n181 ,n1097);
    nand g1203(n1565 ,n1040 ,n551);
    nor g1204(n300 ,n181 ,n243);
    nand g1205(n1625 ,n967 ,n794);
    nor g1206(n192 ,n131 ,n58[1]);
    buf g1207(n9[2], 1'b0);
    nand g1208(n730 ,n452 ,n490);
    nand g1209(n660 ,n27[2] ,n486);
    dff g1210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1679), .Q(n37[3]));
    not g1211(n141 ,n49[0]);
    nand g1212(n1462 ,n25[5] ,n1106);
    not g1213(n264 ,n263);
    nand g1214(n1847 ,n1687 ,n1698);
    nand g1215(n1177 ,n876 ,n875);
    nand g1216(n644 ,n53[2] ,n370);
    or g1217(n1098 ,n423 ,n724);
    buf g1218(n725 ,n246);
    nand g1219(n830 ,n53[1] ,n408);
    nand g1220(n1241 ,n880 ,n531);
    nand g1221(n851 ,n33[2] ,n404);
    or g1222(n1262 ,n156 ,n1109);
    not g1223(n182 ,n183);
    nand g1224(n1702 ,n1291 ,n1290);
    nand g1225(n1127 ,n465 ,n922);
    nor g1226(n75 ,n57[3] ,n73);
    nand g1227(n580 ,n51[3] ,n401);
    nand g1228(n911 ,n47[2] ,n417);
    not g1229(n93 ,n92);
    nand g1230(n880 ,n52[6] ,n484);
    nand g1231(n1242 ,n695 ,n701);
    or g1232(n1406 ,n179 ,n1109);
    nand g1233(n1136 ,n792 ,n611);
    nand g1234(n463 ,n6[7] ,n310);
    nand g1235(n1465 ,n25[2] ,n1106);
    nand g1236(n1612 ,n1065 ,n776);
    nand g1237(n1609 ,n1062 ,n771);
    nand g1238(n220 ,n131 ,n199);
    dff g1239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n961), .Q(n57[4]));
    dff g1240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1615), .Q(n47[6]));
    nand g1241(n629 ,n52[6] ,n384);
    nand g1242(n1669 ,n1002 ,n595);
    nand g1243(n1689 ,n1924 ,n1111);
    or g1244(n497 ,n141 ,n387);
    nor g1245(n712 ,n187 ,n428);
    nand g1246(n748 ,n48[0] ,n395);
    nand g1247(n1214 ,n912 ,n737);
    dff g1248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1772), .Q(n22[2]));
    nor g1249(n484 ,n222 ,n344);
    dff g1250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1611), .Q(n48[3]));
    nand g1251(n970 ,n4[7] ,n715);
    nand g1252(n1035 ,n4[5] ,n711);
    nor g1253(n1873 ,n1712 ,n1711);
    or g1254(n1391 ,n175 ,n1108);
    or g1255(n1866 ,n1178 ,n1707);
    nand g1256(n96 ,n37[1] ,n37[0]);
    dff g1257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1584), .Q(n52[2]));
    nand g1258(n88 ,n57[2] ,n87);
    nand g1259(n858 ,n54[2] ,n394);
    dff g1260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n441), .Q(n17[1]));
    nand g1261(n1493 ,n949 ,n1163);
    dff g1262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1661), .Q(n42[1]));
    nand g1263(n1511 ,n33[6] ,n1109);
    xnor g1264(n1930 ,n58[3] ,n102);
    dff g1265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1768), .Q(n22[6]));
    nand g1266(n998 ,n4[7] ,n709);
    nand g1267(n798 ,n56[5] ,n476);
    nand g1268(n1845 ,n38[2] ,n1484);
    nor g1269(n441 ,n274 ,n290);
    nand g1270(n563 ,n51[2] ,n386);
    nand g1271(n665 ,n45[4] ,n397);
    nand g1272(n865 ,n56[7] ,n476);
    nand g1273(n668 ,n296 ,n459);
    nor g1274(n1863 ,n1137 ,n1703);
    nand g1275(n974 ,n4[3] ,n715);
    nand g1276(n767 ,n23[4] ,n413);
    dff g1277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n809), .Q(n18[2]));
    or g1278(n1398 ,n173 ,n1087);
    dff g1279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1563), .Q(n54[1]));
    nand g1280(n1943 ,n68 ,n67);
    buf g1281(n7[6], n7[7]);
    dff g1282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1841), .Q(n59[2]));
    or g1283(n1422 ,n173 ,n1098);
    nand g1284(n1918 ,n1295 ,n1907);
    nor g1285(n85 ,n57[1] ,n57[0]);
    nand g1286(n684 ,n60[6] ,n420);
    nor g1287(n345 ,n228 ,n243);
    nor g1288(n143 ,n111 ,n50[0]);
    dff g1289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1726), .Q(n30[0]));
    nand g1290(n1517 ,n33[0] ,n1109);
    nand g1291(n564 ,n52[4] ,n384);
    nand g1292(n1844 ,n38[1] ,n1484);
    nor g1293(n1104 ,n429 ,n721);
    nand g1294(n812 ,n44[5] ,n478);
    nand g1295(n1062 ,n4[5] ,n707);
    nand g1296(n1153 ,n844 ,n841);
    nand g1297(n1713 ,n1292 ,n1333);
    nand g1298(n750 ,n22[0] ,n409);
    nand g1299(n1566 ,n28[6] ,n1096);
    nand g1300(n230 ,n40[0] ,n165);
    dff g1301(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1076), .Q(n52[0]));
    nand g1302(n1573 ,n28[3] ,n1096);
    nand g1303(n950 ,n504 ,n515);
    dff g1304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1839), .Q(n22[5]));
    not g1305(n1089 ,n1090);
    nand g1306(n337 ,n1943 ,n248);
    nand g1307(n1180 ,n879 ,n534);
    dff g1308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1825), .Q(n28[5]));
    nand g1309(n904 ,n32[6] ,n414);
    nand g1310(n1047 ,n4[6] ,n713);
    not g1311(n249 ,n250);
    nand g1312(n110 ,n18[2] ,n109);
    not g1313(n281 ,n280);
    nand g1314(n1651 ,n991 ,n829);
    nand g1315(n466 ,n6[0] ,n310);
    nand g1316(n969 ,n4[1] ,n716);
    nand g1317(n1010 ,n4[1] ,n718);
    nand g1318(n1034 ,n4[7] ,n711);
    nand g1319(n1052 ,n4[1] ,n713);
    nand g1320(n1162 ,n675 ,n937);
    nand g1321(n1083 ,n1927 ,n725);
    nand g1322(n1474 ,n24[1] ,n1099);
    nand g1323(n1496 ,n35[5] ,n1087);
    nor g1324(n273 ,n127 ,n230);
    nand g1325(n1888 ,n759 ,n1862);
    nand g1326(n1167 ,n882 ,n827);
    nand g1327(n1003 ,n4[2] ,n709);
    nand g1328(n1620 ,n1074 ,n608);
    nand g1329(n1694 ,n434 ,n1253);
    dff g1330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1793), .Q(n32[5]));
    dff g1331(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1627), .Q(n46[1]));
    nand g1332(n1170 ,n1935 ,n704);
    nand g1333(n666 ,n54[5] ,n392);
    dff g1334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1595), .Q(n50[5]));
    nand g1335(n989 ,n4[2] ,n712);
    nand g1336(n446 ,n18[0] ,n345);
    not g1337(n118 ,n37[0]);
    nand g1338(n967 ,n4[3] ,n716);
    dff g1339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n169), .Q(n7[7]));
    nor g1340(n305 ,n17[2] ,n253);
    nand g1341(n1572 ,n1043 ,n651);
    dff g1342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1567), .Q(n53[6]));
    nand g1343(n509 ,n153 ,n371);
    dff g1344(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n529), .Q(n18[0]));
    nand g1345(n1562 ,n1017 ,n549);
    nor g1346(n74 ,n57[2] ,n57[0]);
    dff g1347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1077), .Q(n53[0]));
    nand g1348(n1626 ,n968 ,n795);
    nand g1349(n351 ,n37[3] ,n280);
    nand g1350(n891 ,n52[4] ,n484);
    nand g1351(n234 ,n1954 ,n165);
    nand g1352(n1146 ,n633 ,n630);
    buf g1353(n8[2], 1'b0);
    nand g1354(n635 ,n43[1] ,n376);
    nor g1355(n707 ,n185 ,n427);
    nand g1356(n899 ,n35[1] ,n481);
    dff g1357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1748), .Q(n25[2]));
    dff g1358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1669), .Q(n41[3]));
    dff g1359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1911), .Q(n6[2]));
    not g1360(n170 ,n171);
    nand g1361(n1854 ,n1677 ,n1315);
    nand g1362(n1619 ,n1073 ,n606);
    not g1363(n115 ,n59[2]);
    nand g1364(n1181 ,n936 ,n855);
    nand g1365(n1644 ,n986 ,n632);
    nand g1366(n1519 ,n32[6] ,n1101);
    dff g1367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1624), .Q(n46[4]));
    nand g1368(n1684 ,n339 ,n1170);
    nand g1369(n260 ,n140 ,n210);
    nand g1370(n1189 ,n798 ,n884);
    nand g1371(n1058 ,n4[2] ,n708);
    or g1372(n1868 ,n1186 ,n1710);
    nand g1373(n628 ,n51[1] ,n401);
    nand g1374(n1920 ,n1349 ,n1901);
    nand g1375(n1081 ,n232 ,n527);
    nand g1376(n801 ,n33[3] ,n404);
    nand g1377(n786 ,n50[0] ,n412);
    nand g1378(n901 ,n50[5] ,n412);
    nand g1379(n267 ,n59[0] ,n218);
    nand g1380(n1032 ,n4[4] ,n705);
    nand g1381(n937 ,n42[2] ,n403);
    nand g1382(n565 ,n51[4] ,n386);
    nand g1383(n350 ,n37[3] ,n261);
    dff g1384(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1544), .Q(n55[5]));
    nor g1385(n316 ,n254 ,n251);
    or g1386(n1283 ,n179 ,n1096);
    nand g1387(n1376 ,n178 ,n1100);
    not g1388(n122 ,n18[3]);
    nor g1389(n495 ,n147 ,n474);
    nand g1390(n1178 ,n885 ,n648);
    not g1391(n703 ,n704);
    nand g1392(n333 ,n1940 ,n249);
    nand g1393(n1634 ,n976 ,n624);
    nand g1394(n1755 ,n1472 ,n1378);
    nand g1395(n618 ,n27[7] ,n486);
    nor g1396(n1347 ,n1239 ,n1238);
    nand g1397(n641 ,n25[2] ,n415);
    nand g1398(n1944 ,n71 ,n70);
    or g1399(n1434 ,n183 ,n1094);
    nand g1400(n1691 ,n1922 ,n1111);
    nand g1401(n825 ,n50[1] ,n412);
    nand g1402(n84 ,n36[3] ,n83);
    nand g1403(n595 ,n41[3] ,n372);
    or g1404(n222 ,n58[2] ,n195);
    dff g1405(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1824), .Q(n28[6]));
    nand g1406(n1233 ,n799 ,n780);
    nor g1407(n1012 ,n38[0] ,n703);
    nand g1408(n789 ,n46[7] ,n480);
    nand g1409(n759 ,n28[4] ,n487);
    dff g1410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1834), .Q(n21[4]));
    nor g1411(n315 ,n228 ,n244);
    nand g1412(n196 ,n19[1] ,n134);
    nor g1413(n1296 ,n1136 ,n1135);
    nand g1414(n223 ,n205 ,n193);
    dff g1415(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1757), .Q(n24[1]));
    or g1416(n1289 ,n173 ,n1096);
    nand g1417(n68 ,n57[1] ,n57[0]);
    nand g1418(n941 ,n49[6] ,n418);
    nor g1419(n1332 ,n1198 ,n1197);
    nand g1420(n965 ,n4[5] ,n716);
    nand g1421(n766 ,n34[4] ,n411);
    nand g1422(n1954 ,n77 ,n78);
    nand g1423(n626 ,n43[2] ,n419);
    nand g1424(n723 ,n1 ,n367);
    nor g1425(n1293 ,n1130 ,n1128);
    or g1426(n1301 ,n171 ,n1095);
    nand g1427(n1358 ,n178 ,n1092);
    nand g1428(n688 ,n21[0] ,n406);
    dff g1429(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1597), .Q(n50[3]));
    nand g1430(n1738 ,n1455 ,n1365);
    nor g1431(n1291 ,n1121 ,n1116);
    nand g1432(n907 ,n52[2] ,n484);
    nor g1433(n709 ,n157 ,n428);
    nand g1434(n244 ,n193 ,n216);
    nand g1435(n637 ,n43[4] ,n419);
    nand g1436(n1215 ,n945 ,n911);
    dff g1437(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1579), .Q(n52[6]));
    nand g1438(n1068 ,n4[7] ,n706);
    nand g1439(n1727 ,n1444 ,n1423);
    or g1440(n1264 ,n156 ,n1098);
    not g1441(n1099 ,n1100);
    dff g1442(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1734), .Q(n27[0]));
    nor g1443(n704 ,n36[4] ,n431);
    nand g1444(n1375 ,n170 ,n1100);
    dff g1445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1617), .Q(n47[4]));
    nor g1446(n285 ,n181 ,n244);
    nand g1447(n1152 ,n891 ,n643);
    nand g1448(n1371 ,n176 ,n1107);
    nand g1449(n756 ,n54[0] ,n394);
    nand g1450(n1659 ,n996 ,n837);
    nand g1451(n814 ,n44[4] ,n478);
    nand g1452(n1442 ,n30[1] ,n1094);
    dff g1453(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1731), .Q(n27[3]));
    dff g1454(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1836), .Q(n21[2]));
    nand g1455(n1360 ,n174 ,n1092);
    not g1456(n124 ,n5[0]);
    dff g1457(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1699), .Q(n38[0]));
    nor g1458(n78 ,n36[3] ,n76);
    nand g1459(n579 ,n50[4] ,n380);
    nand g1460(n843 ,n60[1] ,n396);
    nand g1461(n1132 ,n784 ,n609);
    nand g1462(n1761 ,n1478 ,n1383);
    nor g1463(n207 ,n190 ,n186);
    nand g1464(n436 ,n37[3] ,n310);
    or g1465(n1276 ,n177 ,n1097);
    or g1466(n1397 ,n175 ,n1087);
    not g1467(n123 ,n2);
    nand g1468(n1700 ,n1273 ,n1272);
    nand g1469(n1513 ,n33[4] ,n1109);
    nand g1470(n841 ,n32[2] ,n414);
    nor g1471(n1902 ,n1139 ,n1893);
    nand g1472(n1544 ,n1035 ,n538);
    not g1473(n949 ,n863);
    dff g1474(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1592), .Q(n51[1]));
    nand g1475(n648 ,n51[6] ,n401);
    nand g1476(n1843 ,n1688 ,n1324);
    nand g1477(n1810 ,n1497 ,n1396);
    dff g1478(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1798), .Q(n32[0]));
    or g1479(n1394 ,n171 ,n1087);
    xnor g1480(n1952 ,n18[2] ,n108);
    nand g1481(n1231 ,n786 ,n925);
    nand g1482(n1082 ,n1930 ,n726);
    nand g1483(n1036 ,n4[4] ,n711);
    nand g1484(n608 ,n47[1] ,n390);
    nor g1485(n404 ,n213 ,n351);
    nand g1486(n1857 ,n1674 ,n1312);
    not g1487(n162 ,n161);
    nand g1488(n1060 ,n4[7] ,n707);
    nand g1489(n1217 ,n915 ,n843);
    nor g1490(n1950 ,n81 ,n79);
    dff g1491(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1832), .Q(n21[6]));
    or g1492(n1410 ,n173 ,n1109);
    dff g1493(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n361), .Q(n39[3]));
    dff g1494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1742), .Q(n26[0]));
    nor g1495(n508 ,n144 ,n477);
    nand g1496(n1846 ,n38[3] ,n1484);
    or g1497(n1351 ,n171 ,n1094);
    nand g1498(n796 ,n46[2] ,n485);
    nand g1499(n1798 ,n1525 ,n1263);
    nand g1500(n780 ,n22[6] ,n409);
    nand g1501(n1024 ,n4[1] ,n719);
    nand g1502(n1564 ,n28[7] ,n1096);
    buf g1503(n8[4], 1'b0);
    dff g1504(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1583), .Q(n52[3]));
    nand g1505(n1675 ,n20[3] ,n1105);
    nand g1506(n794 ,n46[3] ,n480);
    nor g1507(n1294 ,n1134 ,n1133);
    nand g1508(n1553 ,n1013 ,n689);
    nor g1509(n1100 ,n429 ,n722);
    nor g1510(n1272 ,n1252 ,n1244);
    dff g1511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1818), .Q(n29[4]));
    nand g1512(n1919 ,n1347 ,n1904);
    nand g1513(n1579 ,n1020 ,n629);
    dff g1514(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n358), .Q(n39[5]));
    nand g1515(n873 ,n44[5] ,n398);
    nor g1516(n66 ,n36[3] ,n64);
    dff g1517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1618), .Q(n47[3]));
    nand g1518(n1670 ,n1003 ,n655);
    nand g1519(n655 ,n41[2] ,n372);
    nand g1520(n478 ,n255 ,n352);
    nand g1521(n443 ,n1952 ,n315);
    nor g1522(n252 ,n111 ,n215);
    nor g1523(n145 ,n111 ,n52[0]);
    nand g1524(n1723 ,n1440 ,n1354);
    dff g1525(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1752), .Q(n24[6]));
    nand g1526(n1667 ,n1001 ,n653);
    nand g1527(n516 ,n153 ,n389);
    dff g1528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1539), .Q(n56[3]));
    nand g1529(n1640 ,n982 ,n856);
    nand g1530(n1522 ,n32[3] ,n1101);
    nor g1531(n1316 ,n1154 ,n1157);
    nand g1532(n645 ,n20[7] ,n405);
    nand g1533(n1218 ,n646 ,n642);
    not g1534(n224 ,n223);
    nor g1535(n1290 ,n1117 ,n1115);
    nor g1536(n1093 ,n425 ,n724);
    nand g1537(n1772 ,n1490 ,n1392);
    nor g1538(n211 ,n190 ,n187);
    nand g1539(n1740 ,n1457 ,n1367);
    nand g1540(n384 ,n255 ,n317);
    nand g1541(n1780 ,n1507 ,n1403);
    dff g1542(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1733), .Q(n27[1]));
    nand g1543(n1490 ,n22[2] ,n1108);
    nor g1544(n398 ,n220 ,n344);
    nor g1545(n1273 ,n1248 ,n1249);
    or g1546(n1307 ,n173 ,n1095);
    nand g1547(n605 ,n47[3] ,n390);
    nor g1548(n1903 ,n1215 ,n1885);
    nand g1549(n1561 ,n29[0] ,n1097);
    nand g1550(n1721 ,n1438 ,n1352);
    dff g1551(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1670), .Q(n41[2]));
    dff g1552(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1546), .Q(n55[4]));
    nand g1553(n1158 ,n672 ,n669);
    nand g1554(n1588 ,n1048 ,n572);
    nor g1555(n289 ,n171 ,n244);
    nand g1556(n1038 ,n4[2] ,n711);
    nand g1557(n1184 ,n908 ,n658);
    dff g1558(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n284), .Q(n7[4]));
    not g1559(n64 ,n63);
    nand g1560(n1498 ,n35[3] ,n1087);
    dff g1561(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1645), .Q(n43[4]));
    dff g1562(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1602), .Q(n49[5]));
    nand g1563(n1379 ,n180 ,n1100);
    nand g1564(n462 ,n6[1] ,n310);
    nand g1565(n737 ,n30[6] ,n399);
    nor g1566(n72 ,n57[3] ,n70);
    or g1567(n1282 ,n171 ,n1096);
    nor g1568(n719 ,n187 ,n489);
    nand g1569(n1173 ,n847 ,n905);
    nand g1570(n1632 ,n974 ,n622);
    nand g1571(n1002 ,n4[3] ,n709);
    nor g1572(n225 ,n204 ,n197);
    nand g1573(n995 ,n4[3] ,n710);
    nand g1574(n431 ,n225 ,n321);
    nand g1575(n1815 ,n1545 ,n1271);
    dff g1576(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1642), .Q(n43[7]));
    nand g1577(n593 ,n27[4] ,n486);
    nand g1578(n1638 ,n980 ,n814);
    nand g1579(n521 ,n153 ,n385);
    nor g1580(n1896 ,n1127 ,n1888);
    nor g1581(n261 ,n37[0] ,n234);
    nand g1582(n1832 ,n1650 ,n1301);
    nor g1583(n283 ,n175 ,n244);
    xnor g1584(n1929 ,n58[2] ,n100);
    not g1585(n1111 ,n250);
    nand g1586(n1227 ,n849 ,n692);
    nand g1587(n646 ,n55[1] ,n416);
    or g1588(n1312 ,n177 ,n1105);
    nand g1589(n1636 ,n978 ,n811);
    buf g1590(n9[5], 1'b0);
    nand g1591(n1611 ,n1064 ,n775);
    dff g1592(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1572), .Q(n53[3]));
    dff g1593(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1541), .Q(n56[1]));
    not g1594(n97 ,n96);
    nand g1595(n1914 ,n1288 ,n1895);
    nand g1596(n931 ,n47[0] ,n417);
    nand g1597(n1802 ,n1529 ,n1419);
    dff g1598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1777), .Q(n34[5]));
    or g1599(n1300 ,n183 ,n1095);
    nand g1600(n1733 ,n1449 ,n1362);
    dff g1601(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n189), .Q(n10[7]));
    nand g1602(n525 ,n60[5] ,n420);
    xnor g1603(n1953 ,n18[3] ,n110);
    not g1604(n198 ,n197);
    dff g1605(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1740), .Q(n26[2]));
    dff g1606(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n439), .Q(n17[0]));
    nand g1607(n952 ,n505 ,n514);
    or g1608(n1306 ,n181 ,n1095);
    nand g1609(n329 ,n1939 ,n249);
    nor g1610(n269 ,n112 ,n235);
    nand g1611(n1362 ,n172 ,n1092);
    nand g1612(n368 ,n120 ,n315);
    dff g1613(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1587), .Q(n51[6]));
    or g1614(n958 ,n498 ,n499);
    nor g1615(n1090 ,n422 ,n724);
    nand g1616(n1716 ,n1342 ,n1341);
    nand g1617(n1776 ,n1503 ,n1399);
    nand g1618(n870 ,n52[7] ,n484);
    nand g1619(n934 ,n52[0] ,n484);
    nand g1620(n447 ,n58[3] ,n313);
    nand g1621(n480 ,n256 ,n352);
    nand g1622(n1783 ,n1510 ,n1431);
    nand g1623(n1440 ,n30[3] ,n1094);
    nand g1624(n1459 ,n26[0] ,n1103);
    nand g1625(n1543 ,n1067 ,n681);
    not g1626(n153 ,n154);
    nand g1627(n990 ,n4[1] ,n712);
    dff g1628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1783), .Q(n33[7]));
    nand g1629(n453 ,n6[5] ,n310);
    dff g1630(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1721), .Q(n30[5]));
    nand g1631(n1453 ,n26[6] ,n1103);
    nand g1632(n604 ,n47[4] ,n390);
    dff g1633(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1854), .Q(n20[1]));
    nand g1634(n1728 ,n1445 ,n1357);
    nand g1635(n758 ,n35[0] ,n481);
    nand g1636(n1674 ,n20[4] ,n1105);
    nand g1637(n571 ,n51[7] ,n386);
    nor g1638(n1344 ,n1182 ,n1181);
    nand g1639(n836 ,n42[3] ,n475);
    nand g1640(n1850 ,n1678 ,n1270);
    nand g1641(n1880 ,n1318 ,n1872);
    nand g1642(n1207 ,n558 ,n902);
    dff g1643(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1693), .Q(n58[2]));
    nand g1644(n467 ,n6[3] ,n310);
    nand g1645(n1168 ,n864 ,n862);
    nand g1646(n842 ,n34[6] ,n411);
    dff g1647(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1797), .Q(n32[1]));
    nor g1648(n1339 ,n1214 ,n1209);
    nand g1649(n600 ,n47[7] ,n390);
    nand g1650(n1838 ,n1665 ,n1269);
    nand g1651(n1157 ,n850 ,n663);
    nand g1652(n1009 ,n1925 ,n725);
    nand g1653(n1685 ,n36[2] ,n1110);
    nand g1654(n1426 ,n182 ,n1100);
    dff g1655(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n359), .Q(n39[2]));
    nand g1656(n1557 ,n29[2] ,n1097);
    nand g1657(n592 ,n49[1] ,n388);
    dff g1658(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1606), .Q(n49[1]));
    nand g1659(n1130 ,n770 ,n767);
    nand g1660(n520 ,n153 ,n379);
    dff g1661(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1609), .Q(n48[5]));
    or g1662(n1412 ,n179 ,n1101);
    or g1663(n363 ,n301 ,n289);
    nor g1664(n399 ,n233 ,n350);
    nand g1665(n943 ,n457 ,n311);
    nor g1666(n79 ,n36[1] ,n36[0]);
    nand g1667(n695 ,n25[6] ,n415);
    nor g1668(n1328 ,n1152 ,n1192);
    nand g1669(n1569 ,n1042 ,n553);
    nand g1670(n1622 ,n964 ,n790);
    not g1671(n180 ,n181);
    nand g1672(n909 ,n32[5] ,n414);
    nor g1673(n140 ,n36[1] ,n36[2]);
    nand g1674(n1195 ,n807 ,n805);
    dff g1675(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1694), .Q(n58[1]));
    nor g1676(n412 ,n236 ,n344);
    nor g1677(n1435 ,n111 ,n1081);
    or g1678(n951 ,n503 ,n502);
    nand g1679(n1464 ,n25[3] ,n1106);
    nand g1680(n1731 ,n1448 ,n1360);
    nand g1681(n276 ,n11 ,n229);
    nand g1682(n1071 ,n4[4] ,n706);
    nand g1683(n1185 ,n761 ,n625);
    nand g1684(n649 ,n41[7] ,n372);
    nand g1685(n848 ,n53[6] ,n408);
    nand g1686(n1128 ,n766 ,n586);
    not g1687(n1942 ,n90);
    nand g1688(n1693 ,n471 ,n1254);
    not g1689(n83 ,n82);
    nand g1690(n327 ,n59[0] ,n252);
    nand g1691(n1174 ,n868 ,n678);
    nand g1692(n1117 ,n769 ,n593);
    nand g1693(n1066 ,n4[1] ,n707);
    nand g1694(n186 ,n59[2] ,n133);
    nand g1695(n1623 ,n965 ,n791);
    nand g1696(n582 ,n55[4] ,n374);
    dff g1697(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1750), .Q(n25[0]));
    dff g1698(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1654), .Q(n42[5]));
    nand g1699(n1646 ,n988 ,n693);
    xor g1700(n1945 ,n57[3] ,n69);
    nand g1701(n988 ,n4[3] ,n712);
    nand g1702(n1631 ,n973 ,n621);
    dff g1703(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1847), .Q(n36[1]));
    nand g1704(n1141 ,n810 ,n808);
    nand g1705(n764 ,n46[3] ,n485);
    not g1706(n132 ,n36[4]);
    not g1707(n130 ,n40[1]);
    nand g1708(n1610 ,n1063 ,n774);
    nand g1709(n918 ,n52[5] ,n484);
    nand g1710(n259 ,n148 ,n209);
    dff g1711(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n957), .Q(n41[0]));
    dff g1712(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1790), .Q(n33[0]));
    dff g1713(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1774), .Q(n22[0]));
    nand g1714(n1363 ,n170 ,n1104);
    nand g1715(n1467 ,n25[0] ,n1106);
    dff g1716(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1613), .Q(n48[1]));
    dff g1717(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1782), .Q(n34[0]));
    dff g1718(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n363), .Q(n39[6]));
    nand g1719(n966 ,n4[4] ,n716);
    nand g1720(n1530 ,n31[3] ,n1098);
    dff g1721(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1628), .Q(n45[7]));
    nand g1722(n1126 ,n898 ,n938);
    nor g1723(n298 ,n179 ,n243);
    nand g1724(n1599 ,n1010 ,n583);
    nor g1725(n63 ,n36[2] ,n61);
    or g1726(n1267 ,n156 ,n1097);
    nand g1727(n888 ,n60[4] ,n396);
    dff g1728(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1724), .Q(n30[2]));
    nand g1729(n920 ,n54[1] ,n394);
    nor g1730(n147 ,n111 ,n42[0]);
    or g1731(n1409 ,n181 ,n1109);
    nor g1732(n254 ,n40[1] ,n232);
    nand g1733(n769 ,n33[4] ,n404);
    nor g1734(n91 ,n59[1] ,n59[0]);
    nand g1735(n1151 ,n839 ,n641);
    nor g1736(n321 ,n111 ,n244);
    nand g1737(n450 ,n18[2] ,n345);
    nand g1738(n857 ,n23[1] ,n413);
    nor g1739(n528 ,n325 ,n468);
    nand g1740(n621 ,n45[4] ,n382);
    nand g1741(n1744 ,n1461 ,n1369);
    nand g1742(n1065 ,n4[2] ,n707);
    nand g1743(n610 ,n51[4] ,n401);
    nand g1744(n1837 ,n1662 ,n1307);
    nand g1745(n1427 ,n182 ,n1090);
    nand g1746(n1751 ,n1468 ,n1426);
    dff g1747(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n202), .Q(n7[1]));
    nand g1748(n1856 ,n1675 ,n1313);
    nor g1749(n1484 ,n704 ,n1088);
    nand g1750(n821 ,n56[4] ,n476);
    nor g1751(n240 ,n59[0] ,n235);
    dff g1752(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1781), .Q(n34[1]));
    nand g1753(n1515 ,n33[2] ,n1109);
    nor g1754(n485 ,n219 ,n344);
    dff g1755(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1835), .Q(n21[3]));
    nand g1756(n833 ,n28[2] ,n487);
    nand g1757(n736 ,n30[5] ,n399);
    buf g1758(n10[2], 1'b0);
    or g1759(n194 ,n117 ,n38[2]);
    or g1760(n1408 ,n175 ,n1109);
    nand g1761(n1524 ,n32[1] ,n1101);
    dff g1762(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1831), .Q(n21[7]));
    dff g1763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1651), .Q(n42[7]));
    nand g1764(n932 ,n42[0] ,n403);
    nand g1765(n878 ,n33[5] ,n404);
    dff g1766(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1725), .Q(n30[1]));
    nand g1767(n778 ,n32[3] ,n414);
    dff g1768(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1681), .Q(n37[1]));
    dff g1769(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1919), .Q(n60[0]));
    nand g1770(n1365 ,n176 ,n1104);
    nand g1771(n452 ,n57[2] ,n316);
    nand g1772(n1842 ,n326 ,n1689);
    nand g1773(n1607 ,n1060 ,n768);
    nand g1774(n1781 ,n1508 ,n1404);
    nand g1775(n1053 ,n4[7] ,n708);
    nand g1776(n625 ,n45[5] ,n397);
    nand g1777(n1549 ,n1038 ,n567);
    nor g1778(n1922 ,n93 ,n91);
    dff g1779(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1767), .Q(n22[7]));
    nand g1780(n690 ,n56[5] ,n378);
    dff g1781(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1827), .Q(n28[3]));
    dff g1782(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1639), .Q(n44[3]));
    or g1783(n1396 ,n177 ,n1087);
    or g1784(n1402 ,n175 ,n1102);
    nand g1785(n1652 ,n21[5] ,n1095);
    dff g1786(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1745), .Q(n25[5]));
    nand g1787(n1642 ,n984 ,n639);
    nand g1788(n1048 ,n4[5] ,n713);
    nand g1789(n1851 ,n1931 ,n1485);
    nor g1790(n354 ,n112 ,n250);
    nor g1791(n1333 ,n1129 ,n1131);
    or g1792(n1275 ,n179 ,n1097);
    or g1793(n213 ,n37[1] ,n200);
    nand g1794(n964 ,n4[6] ,n716);
    nand g1795(n1746 ,n1463 ,n1371);
    nand g1796(n583 ,n50[1] ,n380);
    dff g1797(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n437), .Q(n59[0]));
    not g1798(n247 ,n248);
    nand g1799(n658 ,n43[5] ,n419);
    nand g1800(n181 ,n39[1] ,n1);
    nand g1801(n1026 ,n4[5] ,n720);
    nand g1802(n526 ,n303 ,n433);
    not g1803(n109 ,n108);
    nand g1804(n1004 ,n4[1] ,n709);
    nand g1805(n1156 ,n458 ,n660);
    nand g1806(n1584 ,n1023 ,n568);
    nor g1807(n1872 ,n1706 ,n1705);
    nand g1808(n1633 ,n975 ,n647);
    nand g1809(n185 ,n59[1] ,n59[2]);
    nand g1810(n749 ,n30[4] ,n399);
    or g1811(n1345 ,n1231 ,n1230);
    nand g1812(n633 ,n26[2] ,n393);
    nand g1813(n1232 ,n924 ,n921);
    nand g1814(n1443 ,n30[0] ,n1094);
    nand g1815(n535 ,n56[1] ,n378);
    nand g1816(n685 ,n41[0] ,n400);
    nand g1817(n104 ,n38[1] ,n38[0]);
    nand g1818(n1229 ,n919 ,n842);
    dff g1819(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1912), .Q(n6[1]));
    nor g1820(n1295 ,n1228 ,n1227);
    dff g1821(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1593), .Q(n50[7]));
    nor g1822(n210 ,n36[3] ,n160);
    nor g1823(n1895 ,n1246 ,n1887);
    not g1824(n1106 ,n1107);
    nand g1825(n1171 ,n865 ,n946);
    dff g1826(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1625), .Q(n46[3]));
    nand g1827(n1542 ,n1034 ,n537);
    nand g1828(n800 ,n50[6] ,n412);
    dff g1829(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1644), .Q(n43[5]));
    nand g1830(n1118 ,n754 ,n659);
    nand g1831(n1552 ,n29[4] ,n1097);
    nor g1832(n708 ,n157 ,n488);
    nand g1833(n1446 ,n27[5] ,n1091);
    nor g1834(n301 ,n183 ,n243);
    nand g1835(n1789 ,n1516 ,n1410);
    nand g1836(n790 ,n46[6] ,n480);
    nand g1837(n679 ,n24[1] ,n410);
    nand g1838(n1724 ,n1441 ,n1355);
    nand g1839(n1463 ,n25[4] ,n1106);
    nand g1840(n1043 ,n4[3] ,n714);
    nand g1841(n1016 ,n4[3] ,n720);
    nand g1842(n1018 ,n4[1] ,n720);
    nand g1843(n1708 ,n1325 ,n1322);
    nand g1844(n1540 ,n1030 ,n691);
    nand g1845(n1582 ,n28[0] ,n1096);
    nand g1846(n862 ,n29[7] ,n407);
    nand g1847(n171 ,n39[5] ,n1);
    nand g1848(n527 ,n227 ,n364);
    nand g1849(n846 ,n22[7] ,n409);
    nand g1850(n188 ,n40[1] ,n1);
    dff g1851(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1848), .Q(n36[2]));
    nand g1852(n1372 ,n174 ,n1107);
    dff g1853(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1814), .Q(n35[0]));
    nand g1854(n930 ,n60[0] ,n396);
    nand g1855(n1029 ,n4[3] ,n705);
    nand g1856(n871 ,n54[7] ,n394);
    dff g1857(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1914), .Q(n6[5]));
    nand g1858(n1472 ,n24[3] ,n1099);
    nor g1859(n99 ,n58[1] ,n58[0]);
    nand g1860(n1210 ,n575 ,n638);
    dff g1861(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1918), .Q(n60[1]));
    nand g1862(n158 ,n130 ,n119);
    nand g1863(n1074 ,n4[1] ,n706);
    nand g1864(n638 ,n41[2] ,n400);
    not g1865(n385 ,n386);
    nand g1866(n1121 ,n753 ,n751);
    dff g1867(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1621), .Q(n46[7]));
    nand g1868(n1777 ,n1504 ,n1400);
    nor g1869(n503 ,n150 ,n479);
    or g1870(n256 ,n111 ,n207);
    nand g1871(n939 ,n30[0] ,n399);
    nor g1872(n511 ,n154 ,n475);
    nand g1873(n1840 ,n322 ,n1691);
    nand g1874(n471 ,n58[2] ,n313);
    nor g1875(n1149 ,n111 ,n948);
    nand g1876(n1688 ,n36[0] ,n1110);
    nand g1877(n277 ,n12 ,n229);
    nand g1878(n701 ,n20[6] ,n405);
    dff g1879(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1753), .Q(n24[5]));
    nand g1880(n575 ,n45[2] ,n397);
    nand g1881(n1595 ,n1007 ,n540);
    nand g1882(n590 ,n49[2] ,n388);
    nand g1883(n1230 ,n787 ,n685);
    nand g1884(n783 ,n28[3] ,n487);
    nor g1885(n476 ,n239 ,n344);
    nand g1886(n1438 ,n30[5] ,n1094);
    dff g1887(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1640), .Q(n44[2]));
    nor g1888(n1323 ,n1224 ,n1175);
    dff g1889(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1877), .Q(n38[2]));
    dff g1890(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1622), .Q(n46[6]));
    dff g1891(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1562), .Q(n54[2]));
    nand g1892(n475 ,n258 ,n352);
    nand g1893(n1454 ,n26[5] ,n1103);
    nand g1894(n594 ,n43[0] ,n419);
    dff g1895(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1598), .Q(n50[2]));
    nand g1896(n902 ,n60[3] ,n396);
    nand g1897(n834 ,n52[1] ,n484);
    not g1898(n121 ,n13);
    not g1899(n159 ,n158);
    or g1900(n1882 ,n1188 ,n1868);
    nand g1901(n1613 ,n1066 ,n777);
    dff g1902(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1601), .Q(n49[6]));
    nand g1903(n1756 ,n1473 ,n1379);
    nand g1904(n1891 ,n698 ,n1871);
    nand g1905(n686 ,n56[3] ,n378);
    nand g1906(n1750 ,n1467 ,n1256);
    nand g1907(n806 ,n29[0] ,n407);
    xor g1908(n1934 ,n36[4] ,n66);
    or g1909(n1277 ,n175 ,n1097);
    dff g1910(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1586), .Q(n51[7]));
    nor g1911(n724 ,n111 ,n472);
    nand g1912(n599 ,n25[7] ,n415);
    nand g1913(n1448 ,n27[3] ,n1091);
    or g1914(n1305 ,n175 ,n1095);
    nand g1915(n175 ,n39[2] ,n1);
    nand g1916(n1196 ,n671 ,n665);
    nand g1917(n1742 ,n1459 ,n1255);
    not g1918(n134 ,n38[0]);
    nor g1919(n307 ,n17[0] ,n253);
    dff g1920(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1915), .Q(n6[7]));
    dff g1921(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n950), .Q(n45[0]));
    nand g1922(n819 ,n49[1] ,n418);
    not g1923(n155 ,n156);
    nor g1924(n1349 ,n1243 ,n1242);
    nand g1925(n1797 ,n1524 ,n1416);
    nor g1926(n332 ,n191 ,n279);
    nand g1927(n62 ,n36[1] ,n36[0]);
    or g1928(n1310 ,n171 ,n1105);
    nand g1929(n913 ,n23[6] ,n413);
    nand g1930(n884 ,n42[5] ,n403);
    nand g1931(n634 ,n43[2] ,n376);
    xnor g1932(n1927 ,n37[3] ,n98);
    nor g1933(n163 ,n58[1] ,n58[2]);
    nand g1934(n1769 ,n1668 ,n1309);
    nand g1935(n1057 ,n4[3] ,n708);
    nand g1936(n1828 ,n1576 ,n1287);
    or g1937(n428 ,n59[3] ,n319);
    not g1938(n430 ,n429);
    nand g1939(n201 ,n8[1] ,n1);
    nor g1940(n715 ,n186 ,n428);
    nand g1941(n810 ,n30[3] ,n399);
    nand g1942(n1804 ,n1531 ,n1421);
    nand g1943(n553 ,n53[5] ,n370);
    dff g1944(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1760), .Q(n23[6]));
    or g1945(n347 ,n37[3] ,n281);
    nand g1946(n382 ,n256 ,n314);
    xnor g1947(n1923 ,n59[2] ,n92);
    nand g1948(n1852 ,n1932 ,n1485);
    nand g1949(n827 ,n49[7] ,n418);
    dff g1950(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1680), .Q(n37[2]));
    nand g1951(n699 ,n27[6] ,n486);
    nor g1952(n150 ,n111 ,n46[0]);
    dff g1953(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1807), .Q(n35[7]));
    nand g1954(n309 ,n1 ,n245);
    nand g1955(n1148 ,n636 ,n823);
    nand g1956(n1369 ,n170 ,n1107);
    nand g1957(n1123 ,n544 ,n757);
    nand g1958(n816 ,n23[3] ,n413);
    dff g1959(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1796), .Q(n32[2]));
    nor g1960(n364 ,n40[0] ,n288);
    nand g1961(n928 ,n46[0] ,n485);
    nand g1962(n914 ,n29[6] ,n407);
    nand g1963(n342 ,n1946 ,n254);
    nand g1964(n947 ,n55[0] ,n416);
    dff g1965(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1766), .Q(n23[0]));
    dff g1966(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1792), .Q(n32[6]));
    nand g1967(n603 ,n55[5] ,n416);
    nor g1968(n286 ,n173 ,n244);
    nand g1969(n1570 ,n1075 ,n654);
    nand g1970(n1912 ,n1350 ,n1898);
    not g1971(n113 ,n59[3]);
    nand g1972(n1541 ,n1031 ,n535);
    nand g1973(n1785 ,n1512 ,n1406);
    nand g1974(n235 ,n59[3] ,n159);
    nand g1975(n1567 ,n1041 ,n673);
    dff g1976(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1555), .Q(n54[6]));
    nand g1977(n894 ,n44[4] ,n398);
    nand g1978(n1877 ,n1845 ,n1852);
    nor g1979(n295 ,n171 ,n243);
    nand g1980(n659 ,n43[7] ,n419);
    nand g1981(n1193 ,n821 ,n820);
    nand g1982(n876 ,n33[7] ,n404);
    nand g1983(n817 ,n47[4] ,n417);
    nand g1984(n515 ,n153 ,n381);
    dff g1985(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1813), .Q(n35[1]));
    nand g1986(n1248 ,n765 ,n736);
    buf g1987(n14, n13);
    nand g1988(n1739 ,n1456 ,n1366);
    nand g1989(n627 ,n26[3] ,n393);
    nand g1990(n643 ,n55[4] ,n416);
    nand g1991(n523 ,n153 ,n391);
    not g1992(n228 ,n229);
    not g1993(n205 ,n204);
    nand g1994(n1357 ,n170 ,n1092);
    nand g1995(n667 ,n60[4] ,n420);
    nor g1996(n328 ,n132 ,n260);
    not g1997(n218 ,n217);
    nand g1998(n1471 ,n24[4] ,n1099);
    nand g1999(n1760 ,n1477 ,n1382);
    nand g2000(n1491 ,n22[1] ,n1108);
    nand g2001(n1246 ,n453 ,n548);
    nand g2002(n677 ,n41[5] ,n400);
    nand g2003(n912 ,n35[6] ,n481);
    nand g2004(n1710 ,n1326 ,n1338);
    dff g2005(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1720), .Q(n30[6]));
    dff g2006(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1607), .Q(n48[7]));
    nor g2007(n1348 ,n1211 ,n1210);
    nand g2008(n866 ,n44[7] ,n398);
    nand g2009(n1523 ,n32[2] ,n1101);
    dff g2010(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1722), .Q(n30[4]));
    dff g2011(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n959), .Q(n49[0]));
    dff g2012(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1549), .Q(n55[2]));
    nand g2013(n763 ,n44[0] ,n398);
    nand g2014(n773 ,n54[5] ,n394);
    nand g2015(n922 ,n32[4] ,n414);
    nand g2016(n689 ,n54[7] ,n392);
    nand g2017(n1686 ,n336 ,n1222);
    nor g2018(n507 ,n154 ,n478);
    dff g2019(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1738), .Q(n26[4]));
    nand g2020(n514 ,n153 ,n377);
    dff g2021(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1435), .Q(n40[0]));
    nand g2022(n772 ,n50[2] ,n412);
    nand g2023(n900 ,n48[3] ,n395);
    dff g2024(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n954), .Q(n47[0]));
    nor g2025(n1338 ,n1184 ,n1144);
    xnor g2026(n304 ,n15 ,n216);
    nand g2027(n893 ,n28[6] ,n487);
    nand g2028(n795 ,n46[2] ,n480);
    nand g2029(n669 ,n20[1] ,n405);
    nand g2030(n1795 ,n1522 ,n1414);
    nand g2031(n1876 ,n1846 ,n1853);
    nand g2032(n1627 ,n969 ,n797);
    nand g2033(n1656 ,n21[4] ,n1095);
    nor g2034(n961 ,n111 ,n528);
    nor g2035(n1308 ,n1151 ,n1150);
    nand g2036(n1112 ,n758 ,n662);
    nand g2037(n226 ,n13 ,n189);
    or g2038(n1352 ,n179 ,n1094);
    nor g2039(n1928 ,n101 ,n99);
    nand g2040(n177 ,n39[3] ,n1);
    nand g2041(n576 ,n51[1] ,n386);
    nand g2042(n1503 ,n34[6] ,n1102);
    not g2043(n432 ,n431);
    dff g2044(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n526), .Q(n37[0]));
    nand g2045(n464 ,n57[1] ,n316);
    nand g2046(n1754 ,n1471 ,n1377);
    dff g2047(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1794), .Q(n32[4]));
    nand g2048(n1067 ,n4[6] ,n711);
    nand g2049(n370 ,n256 ,n318);
    nand g2050(n874 ,n60[6] ,n396);
    nand g2051(n1203 ,n752 ,n580);
    nand g2052(n1025 ,n4[3] ,n719);
    nand g2053(n1819 ,n1554 ,n1277);
    nor g2054(n1326 ,n1194 ,n1185);
    dff g2055(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1542), .Q(n55[7]));
    dff g2056(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1920), .Q(n6[6]));
    nand g2057(n1265 ,n155 ,n1092);
    dff g2058(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1723), .Q(n30[3]));
    dff g2059(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1560), .Q(n54[3]));
    nand g2060(n378 ,n257 ,n317);
    dff g2061(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1908), .Q(n60[5]));
    dff g2062(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1784), .Q(n33[6]));
    nand g2063(n702 ,n153 ,n373);
    nand g2064(n1883 ,n1332 ,n1873);
    nand g2065(n82 ,n36[2] ,n81);
    dff g2066(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1785), .Q(n33[5]));
    nand g2067(n157 ,n133 ,n115);
    or g2068(n494 ,n143 ,n379);
    not g2069(n114 ,n58[1]);
    nand g2070(n1475 ,n24[0] ,n1099);
    or g2071(n239 ,n131 ,n195);
    or g2072(n1433 ,n183 ,n1098);
    dff g2073(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1821), .Q(n29[1]));
    nand g2074(n1839 ,n1487 ,n1389);
    nor g2075(n423 ,n111 ,n292);
    not g2076(n116 ,n37[1]);
    dff g2077(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1630), .Q(n45[5]));
    nand g2078(n908 ,n47[5] ,n417);
    nand g2079(n1558 ,n1015 ,n546);
    nand g2080(n552 ,n25[5] ,n415);
    nand g2081(n1256 ,n155 ,n1107);
    nand g2082(n751 ,n31[4] ,n402);
    nor g2083(n292 ,n191 ,n282);
    or g2084(n1355 ,n181 ,n1094);
    dff g2085(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1574), .Q(n53[2]));
    nand g2086(n341 ,n1944 ,n248);
    nand g2087(n1753 ,n1470 ,n1376);
    nand g2088(n694 ,n43[4] ,n376);
    nand g2089(n1254 ,n1929 ,n726);
    nor g2090(n331 ,n1921 ,n270);
    nor g2091(n502 ,n154 ,n480);
    dff g2092(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1730), .Q(n27[4]));
    nor g2093(n1867 ,n1183 ,n1708);
    nand g2094(n692 ,n45[1] ,n397);
    or g2095(n518 ,n152 ,n391);
    nand g2096(n1581 ,n1022 ,n564);
    nand g2097(n519 ,n153 ,n387);
    not g2098(n371 ,n372);
    nand g2099(n696 ,n21[4] ,n406);
    dff g2100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1610), .Q(n48[4]));
    nand g2101(n1447 ,n27[4] ,n1091);
    nand g2102(n936 ,n46[6] ,n485);
    nor g2103(n1297 ,n1119 ,n1176);
    xnor g2104(n1926 ,n37[2] ,n96);
    dff g2105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1869), .Q(n38[1]));
    dff g2106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1596), .Q(n50[4]));
    nand g2107(n1757 ,n1474 ,n1380);
    dff g2108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n167), .Q(n10[6]));
    or g2109(n318 ,n111 ,n240);
    nand g2110(n1119 ,n800 ,n746);
    nand g2111(n910 ,n32[1] ,n414);
    dff g2112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1735), .Q(n26[7]));
    nand g2113(n1061 ,n4[6] ,n707);
    nand g2114(n586 ,n24[4] ,n410);
    nand g2115(n1915 ,n1334 ,n1900);
    nor g2116(n718 ,n157 ,n489);
    dff g2117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1570), .Q(n53[4]));
    dff g2118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1590), .Q(n51[3]));
    nor g2119(n1330 ,n1193 ,n1145);
    or g2120(n1405 ,n171 ,n1109);
    nand g2121(n1166 ,n889 ,n541);
    nand g2122(n1603 ,n1056 ,n587);
    nand g2123(n1641 ,n983 ,n818);
    nand g2124(n856 ,n44[2] ,n478);
    nand g2125(n1762 ,n1479 ,n1384);
    nor g2126(n77 ,n36[2] ,n36[0]);
    nand g2127(n791 ,n46[5] ,n480);
    nand g2128(n782 ,n29[3] ,n407);
    nand g2129(n1782 ,n1509 ,n1261);
    dff g2130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1614), .Q(n47[7]));
    or g2131(n1263 ,n156 ,n1101);
    nand g2132(n598 ,n21[3] ,n406);
    nor g2133(n1325 ,n1177 ,n1172);
    nand g2134(n380 ,n317 ,n258);
    dff g2135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n943), .Q(n58[0]));
    nand g2136(n1766 ,n1266 ,n1258);
    nand g2137(n1097 ,n424 ,n723);
    nand g2138(n938 ,n47[3] ,n417);
    nor g2139(n1299 ,n1148 ,n1146);
    nor g2140(n481 ,n231 ,n351);
    nand g2141(n1489 ,n22[3] ,n1108);
    nand g2142(n1660 ,n21[2] ,n1095);
    nand g2143(n1122 ,n738 ,n853);
    nand g2144(n1244 ,n732 ,n729);
    nand g2145(n1096 ,n426 ,n723);
    nand g2146(n547 ,n51[6] ,n386);
    nand g2147(n1587 ,n1047 ,n547);
    nand g2148(n607 ,n21[7] ,n406);
    nand g2149(n792 ,n34[3] ,n411);
    nor g2150(n401 ,n222 ,n311);
    nand g2151(n1704 ,n1308 ,n1299);
    nor g2152(n1322 ,n1168 ,n1164);
    or g2153(n76 ,n36[4] ,n36[1]);
    or g2154(n1271 ,n183 ,n1097);
    nand g2155(n1179 ,n886 ,n941);
    nand g2156(n809 ,n450 ,n443);
    nand g2157(n340 ,n1934 ,n246);
    dff g2158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n302), .Q(n40[1]));
    nand g2159(n1211 ,n906 ,n772);
    nand g2160(n372 ,n258 ,n314);
    nand g2161(n539 ,n55[3] ,n374);
    buf g2162(n9[1], 1'b0);
    or g2163(n1712 ,n1196 ,n1331);
    nand g2164(n558 ,n55[3] ,n416);
    nor g2165(n1951 ,n109 ,n107);
    nor g2166(n1280 ,n1226 ,n1235);
    or g2167(n353 ,n38[1] ,n264);
    nand g2168(n335 ,n1949 ,n246);
    nand g2169(n1437 ,n30[6] ,n1094);
    nand g2170(n869 ,n48[5] ,n395);
    nor g2171(n1350 ,n1232 ,n1202);
    nand g2172(n915 ,n56[1] ,n476);
    nand g2173(n640 ,n41[3] ,n400);
    nand g2174(n1531 ,n31[2] ,n1098);
    nand g2175(n1790 ,n1517 ,n1262);
    nand g2176(n1021 ,n4[5] ,n719);
    nand g2177(n548 ,n21[5] ,n406);
    not g2178(n375 ,n376);
    nand g2179(n1532 ,n31[1] ,n1098);
    nand g2180(n1202 ,n910 ,n679);
    nand g2181(n1614 ,n1068 ,n600);
    buf g2182(n10[3], n7[1]);
    nand g2183(n233 ,n37[1] ,n164);
    nand g2184(n683 ,n51[5] ,n401);
    nand g2185(n675 ,n60[1] ,n420);
    or g2186(n1304 ,n177 ,n1095);
    or g2187(n67 ,n57[1] ,n57[0]);
    nand g2188(n1589 ,n1049 ,n565);
    not g2189(n369 ,n370);
    or g2190(n956 ,n495 ,n511);
    not g2191(n491 ,n469);
    nand g2192(n1654 ,n993 ,n832);
    nand g2193(n1225 ,n920 ,n804);
    nand g2194(n1722 ,n1439 ,n1353);
    nand g2195(n1598 ,n1011 ,n581);
    nand g2196(n250 ,n1 ,n215);
    nor g2197(n439 ,n275 ,n307);
    nand g2198(n1460 ,n25[7] ,n1106);
    or g2199(n1417 ,n171 ,n1098);
    nand g2200(n543 ,n50[7] ,n380);
    nand g2201(n253 ,n189 ,n232);
    dff g2202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1637), .Q(n44[5]));
    nor g2203(n720 ,n186 ,n489);
    not g2204(n1094 ,n1093);
    nand g2205(n1805 ,n1532 ,n1422);
    nor g2206(n1897 ,n1124 ,n1894);
    nand g2207(n1359 ,n176 ,n1092);
    nand g2208(n1125 ,n748 ,n928);
    or g2209(n1279 ,n173 ,n1097);
    nand g2210(n1510 ,n33[7] ,n1109);
    nand g2211(n200 ,n37[2] ,n128);
    nand g2212(n572 ,n51[5] ,n386);
    nand g2213(n1576 ,n28[2] ,n1096);
    nand g2214(n1813 ,n1500 ,n1398);
    nand g2215(n753 ,n35[4] ,n481);
    nand g2216(n560 ,n20[4] ,n405);
    nand g2217(n1238 ,n933 ,n554);
    nand g2218(n1105 ,n430 ,n723);
    nand g2219(n944 ,n26[6] ,n393);
    nor g2220(n405 ,n214 ,n346);
    not g2221(n1696 ,n1682);
    or g2222(n1353 ,n177 ,n1094);
    nand g2223(n468 ,n342 ,n278);
    nand g2224(n1650 ,n21[6] ,n1095);
    nand g2225(n760 ,n48[6] ,n483);
    nor g2226(n148 ,n57[1] ,n57[2]);
    nand g2227(n602 ,n47[5] ,n390);
    nand g2228(n173 ,n39[0] ,n1);
    nand g2229(n1050 ,n4[3] ,n713);
    nand g2230(n1663 ,n998 ,n649);
    nand g2231(n1477 ,n23[6] ,n1089);
    not g2232(n389 ,n390);
    nand g2233(n1143 ,n816 ,n627);
    dff g2234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1786), .Q(n33[4]));
    nand g2235(n1535 ,n1033 ,n700);
    nand g2236(n1681 ,n435 ,n1009);
    xnor g2237(n1935 ,n36[2] ,n80);
    nand g2238(n536 ,n55[1] ,n374);
    nand g2239(n1499 ,n35[2] ,n1087);
    dff g2240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1540), .Q(n56[2]));
    nor g2241(n215 ,n190 ,n158);
    nand g2242(n1548 ,n29[6] ,n1097);
    nand g2243(n195 ,n58[1] ,n58[3]);
    nor g2244(n472 ,n194 ,n355);
    nand g2245(n1041 ,n4[6] ,n714);
    dff g2246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n366), .Q(n39[1]));
    nand g2247(n997 ,n4[1] ,n710);
    nand g2248(n651 ,n53[3] ,n370);
    nand g2249(n616 ,n45[7] ,n382);
endmodule
