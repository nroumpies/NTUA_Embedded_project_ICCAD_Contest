module top (n0, n1, n2, n3, n5, n8, n6, n9, n4, n7, n10, n11, n12, n13);
    input n0, n1;
    input [15:0] n2;
    input [7:0] n3, n4;
    input [3:0] n5, n6, n7;
    input [5:0] n8;
    input [1:0] n9;
    output [7:0] n10;
    output [3:0] n11;
    output [1:0] n12;
    output n13;
    wire n0, n1;
    wire [15:0] n2;
    wire [7:0] n3, n4;
    wire [3:0] n5, n6, n7;
    wire [5:0] n8;
    wire [1:0] n9;
    wire [7:0] n10;
    wire [3:0] n11;
    wire [1:0] n12;
    wire n13;
    wire [7:0] n14;
    wire [2:0] n15;
    wire [15:0] n16;
    wire [7:0] n17;
    wire [7:0] n18;
    wire [15:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [15:0] n23;
    wire [15:0] n24;
    wire [15:0] n25;
    wire [15:0] n26;
    wire [7:0] n27;
    wire [7:0] n28;
    wire [7:0] n29;
    wire [7:0] n30;
    wire [15:0] n31;
    wire [7:0] n32;
    wire [15:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [7:0] n36;
    wire [15:0] n37;
    wire [2:0] n38;
    wire [7:0] n39;
    wire [7:0] n40;
    wire [7:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [7:0] n44;
    wire [7:0] n45;
    wire [7:0] n46;
    wire [7:0] n47;
    wire n48, n49, n50, n51, n52, n53, n54, n55;
    wire n56, n57, n58, n59, n60, n61, n62, n63;
    wire n64, n65, n66, n67, n68, n69, n70, n71;
    wire n72, n73, n74, n75, n76, n77, n78, n79;
    wire n80, n81, n82, n83, n84, n85, n86, n87;
    wire n88, n89, n90, n91, n92, n93, n94, n95;
    wire n96, n97, n98, n99, n100, n101, n102, n103;
    wire n104, n105, n106, n107, n108, n109, n110, n111;
    wire n112, n113, n114, n115, n116, n117, n118, n119;
    wire n120, n121, n122, n123, n124, n125, n126, n127;
    wire n128, n129, n130, n131, n132, n133, n134, n135;
    wire n136, n137, n138, n139, n140, n141, n142, n143;
    wire n144, n145, n146, n147, n148, n149, n150, n151;
    wire n152, n153, n154, n155, n156, n157, n158, n159;
    wire n160, n161, n162, n163, n164, n165, n166, n167;
    wire n168, n169, n170, n171, n172, n173, n174, n175;
    wire n176, n177, n178, n179, n180, n181, n182, n183;
    wire n184, n185, n186, n187, n188, n189, n190, n191;
    wire n192, n193, n194, n195, n196, n197, n198, n199;
    wire n200, n201, n202, n203, n204, n205, n206, n207;
    wire n208, n209, n210, n211, n212, n213, n214, n215;
    wire n216, n217, n218, n219, n220, n221, n222, n223;
    wire n224, n225, n226, n227, n228, n229, n230, n231;
    wire n232, n233, n234, n235, n236, n237, n238, n239;
    wire n240, n241, n242, n243, n244, n245, n246, n247;
    wire n248, n249, n250, n251, n252, n253, n254, n255;
    wire n256, n257, n258, n259, n260, n261, n262, n263;
    wire n264, n265, n266, n267, n268, n269, n270, n271;
    wire n272, n273, n274, n275, n276, n277, n278, n279;
    wire n280, n281, n282, n283, n284, n285, n286, n287;
    wire n288, n289, n290, n291, n292, n293, n294, n295;
    wire n296, n297, n298, n299, n300, n301, n302, n303;
    wire n304, n305, n306, n307, n308, n309, n310, n311;
    wire n312, n313, n314, n315, n316, n317, n318, n319;
    wire n320, n321, n322, n323, n324, n325, n326, n327;
    wire n328, n329, n330, n331, n332, n333, n334, n335;
    wire n336, n337, n338, n339, n340, n341, n342, n343;
    wire n344, n345, n346, n347, n348, n349, n350, n351;
    wire n352, n353, n354, n355, n356, n357, n358, n359;
    wire n360, n361, n362, n363, n364, n365, n366, n367;
    wire n368, n369, n370, n371, n372, n373, n374, n375;
    wire n376, n377, n378, n379, n380, n381, n382, n383;
    wire n384, n385, n386, n387, n388, n389, n390, n391;
    wire n392, n393, n394, n395, n396, n397, n398, n399;
    wire n400, n401, n402, n403, n404, n405, n406, n407;
    wire n408, n409, n410, n411, n412, n413, n414, n415;
    wire n416, n417, n418, n419, n420, n421, n422, n423;
    nor g0(n151 ,n64 ,n149);
    nand g1(n231 ,n25[7] ,n200);
    or g2(n247 ,n208 ,n203);
    nand g3(n323 ,n269 ,n268);
    nand g4(n294 ,n240 ,n239);
    xnor g5(n122 ,n2[1] ,n3[1]);
    nand g6(n271 ,n23[2] ,n202);
    xor g7(n145 ,n6[1] ,n40[3]);
    dff g8(.RN(n1), .SN(1'b1), .CK(n0), .D(n134), .Q(n18[2]));
    nand g9(n149 ,n60 ,n59);
    dff g10(.RN(n1), .SN(1'b1), .CK(n0), .D(n24[1]), .Q(n24[3]));
    dff g11(.RN(n1), .SN(1'b1), .CK(n0), .D(n83), .Q(n42[1]));
    nand g12(n163 ,n61 ,n151);
    nand g13(n387 ,n366 ,n386);
    nand g14(n262 ,n23[7] ,n202);
    dff g15(.RN(n1), .SN(1'b1), .CK(n0), .D(n167), .Q(n36[0]));
    nand g16(n309 ,n261 ,n225);
    nand g17(n413 ,n47[1] ,n47[3]);
    nor g18(n376 ,n317 ,n374);
    dff g19(.RN(n1), .SN(1'b1), .CK(n0), .D(n88), .Q(n40[2]));
    nor g20(n366 ,n297 ,n357);
    nand g21(n62 ,n37[12] ,n54);
    dff g22(.RN(n1), .SN(1'b1), .CK(n0), .D(n141), .Q(n37[7]));
    not g23(n55 ,n37[8]);
    dff g24(.RN(n1), .SN(1'b1), .CK(n0), .D(n31[7]), .Q(n30[7]));
    not g25(n204 ,n205);
    dff g26(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[5]), .Q(n26[7]));
    xor g27(n103 ,n8[0] ,n35[0]);
    xor g28(n93 ,n9[0] ,n39[2]);
    dff g29(.RN(n1), .SN(1'b1), .CK(n0), .D(n84), .Q(n41[3]));
    dff g30(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[3]), .Q(n23[5]));
    xor g31(n134 ,n26[2] ,n40[2]);
    xnor g32(n159 ,n109 ,n32[3]);
    dff g33(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[11]), .Q(n33[1]));
    nand g34(n396 ,n330 ,n325);
    dff g35(.RN(n1), .SN(1'b1), .CK(n0), .D(n92), .Q(n39[3]));
    nor g36(n202 ,n15[0] ,n182);
    not g37(n176 ,n15[0]);
    nand g38(n315 ,n271 ,n222);
    nand g39(n420 ,n416 ,n411);
    nor g40(n207 ,n175 ,n178);
    nand g41(n245 ,n17[6] ,n208);
    dff g42(.RN(n1), .SN(1'b1), .CK(n0), .D(n174), .Q(n29[2]));
    xnor g43(n194 ,n37[2] ,n16[2]);
    nor g44(n243 ,n388 ,n204);
    nand g45(n274 ,n22[0] ,n200);
    dff g46(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[7]), .Q(n18[7]));
    not g47(n388 ,n14[6]);
    buf g48(n12[0], 1'b0);
    nor g49(n337 ,n243 ,n293);
    nand g50(n280 ,n20[1] ,n201);
    not g51(n56 ,n37[14]);
    dff g52(.RN(n1), .SN(1'b1), .CK(n0), .D(n157), .Q(n37[0]));
    xor g53(n143 ,n16[1] ,n42[1]);
    xor g54(n96 ,n7[0] ,n39[0]);
    nand g55(n237 ,n22[1] ,n200);
    xnor g56(n173 ,n163 ,n29[3]);
    xor g57(n89 ,n4[1] ,n40[1]);
    or g58(n178 ,n15[0] ,n15[1]);
    nand g59(n269 ,n25[2] ,n200);
    xor g60(n153 ,n119 ,n120);
    dff g61(.RN(n1), .SN(1'b1), .CK(n0), .D(n138), .Q(n37[6]));
    dff g62(.RN(n1), .SN(1'b1), .CK(n0), .D(n77), .Q(n45[2]));
    xor g63(n126 ,n19[2] ,n39[2]);
    xnor g64(n193 ,n16[1] ,n37[1]);
    xor g65(n102 ,n23[2] ,n45[2]);
    or g66(n340 ,n304 ,n398);
    nand g67(n218 ,n30[6] ,n207);
    nand g68(n214 ,n33[7] ,n206);
    nand g69(n284 ,n14[3] ,n205);
    nand g70(n285 ,n17[1] ,n208);
    dff g71(.RN(n1), .SN(1'b1), .CK(n0), .D(n37[6]), .Q(n37[14]));
    dff g72(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[1]), .Q(n23[3]));
    nand g73(n253 ,n19[6] ,n201);
    nand g74(n311 ,n265 ,n264);
    nor g75(n336 ,n321 ,n320);
    dff g76(.RN(n1), .SN(1'b1), .CK(n0), .D(n86), .Q(n30[2]));
    dff g77(.RN(n1), .SN(1'b1), .CK(n0), .D(n159), .Q(n21[3]));
    dff g78(.RN(n1), .SN(1'b1), .CK(n0), .D(n90), .Q(n40[0]));
    nand g79(n288 ,n230 ,n284);
    dff g80(.RN(n1), .SN(1'b1), .CK(n0), .D(n79), .Q(n44[2]));
    nor g81(n384 ,n365 ,n379);
    nand g82(n302 ,n252 ,n251);
    nand g83(n320 ,n224 ,n280);
    not g84(n407 ,n1);
    xor g85(n87 ,n8[5] ,n35[5]);
    dff g86(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[5]), .Q(n25[7]));
    dff g87(.RN(n1), .SN(1'b1), .CK(n0), .D(n162), .Q(n22[3]));
    xnor g88(n342 ,n186 ,n393);
    nand g89(n215 ,n30[2] ,n207);
    nor g90(n65 ,n57 ,n37[15]);
    or g91(n397 ,n298 ,n295);
    dff g92(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[3]), .Q(n16[5]));
    dff g93(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[2]), .Q(n16[4]));
    or g94(n392 ,n308 ,n339);
    xor g95(n99 ,n8[1] ,n35[1]);
    xnor g96(n71 ,n8[2] ,n35[2]);
    dff g97(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[4]), .Q(n25[6]));
    dff g98(.RN(n1), .SN(1'b1), .CK(n0), .D(n158), .Q(n33[0]));
    nand g99(n306 ,n258 ,n219);
    xnor g100(n121 ,n5[2] ,n21[2]);
    dff g101(.RN(n1), .SN(1'b1), .CK(n0), .D(n38[0]), .Q(n15[0]));
    dff g102(.RN(n1), .SN(1'b1), .CK(n0), .D(n161), .Q(n21[2]));
    dff g103(.RN(n1), .SN(1'b1), .CK(n0), .D(n31[4]), .Q(n31[6]));
    xor g104(n125 ,n19[3] ,n39[3]);
    nand g105(n380 ,n208 ,n370);
    xnor g106(n183 ,n21[1] ,n22[1]);
    xor g107(n88 ,n9[1] ,n40[2]);
    xnor g108(n111 ,n2[3] ,n3[3]);
    nand g109(n246 ,n29[3] ,n207);
    dff g110(.RN(n1), .SN(1'b1), .CK(n0), .D(n31[6]), .Q(n30[6]));
    dff g111(.RN(n1), .SN(1'b1), .CK(n0), .D(n392), .Q(n10[7]));
    xor g112(n132 ,n5[1] ,n21[1]);
    nor g113(n199 ,n176 ,n177);
    nand g114(n276 ,n20[7] ,n201);
    xnor g115(n353 ,n189 ,n344);
    dff g116(.RN(n1), .SN(1'b1), .CK(n0), .D(n145), .Q(n40[3]));
    not g117(n354 ,n353);
    nor g118(n329 ,n303 ,n302);
    dff g119(.RN(n1), .SN(1'b1), .CK(n0), .D(n155), .Q(n26[0]));
    xor g120(n345 ,n198 ,n389);
    xnor g121(n368 ,n187 ,n356);
    nand g122(n236 ,n21[1] ,n202);
    nand g123(n229 ,n30[3] ,n207);
    dff g124(.RN(n408), .SN(1'b1), .CK(n0), .D(n404), .Q(n47[0]));
    xnor g125(n116 ,n2[4] ,n3[2]);
    nand g126(n304 ,n255 ,n210);
    xor g127(n141 ,n2[7] ,n3[7]);
    xor g128(n155 ,n113 ,n114);
    dff g129(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[7]), .Q(n28[7]));
    nor g130(n326 ,n309 ,n307);
    xor g131(n79 ,n7[1] ,n44[2]);
    dff g132(.RN(n408), .SN(1'b1), .CK(n0), .D(n401), .Q(n47[3]));
    dff g133(.RN(n1), .SN(1'b1), .CK(n0), .D(n154), .Q(n24[0]));
    nand g134(n349 ,n201 ,n342);
    dff g135(.RN(n1), .SN(1'b1), .CK(n0), .D(n95), .Q(n39[1]));
    nand g136(n268 ,n24[2] ,n208);
    xnor g137(n369 ,n193 ,n359);
    dff g138(.RN(n1), .SN(1'b1), .CK(n0), .D(n24[7]), .Q(n17[7]));
    xor g139(n92 ,n6[0] ,n39[3]);
    dff g140(.RN(n1), .SN(1'b1), .CK(n0), .D(n38[2]), .Q(n15[2]));
    dff g141(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[13]), .Q(n23[1]));
    nand g142(n182 ,n15[2] ,n15[1]);
    or g143(n421 ,n419 ,n420);
    nand g144(n415 ,n398 ,n400);
    nor g145(n410 ,n47[0] ,n47[2]);
    dff g146(.RN(n1), .SN(1'b1), .CK(n0), .D(n97), .Q(n25[0]));
    xor g147(n123 ,n4[7] ,n46[3]);
    not g148(n54 ,n37[11]);
    xnor g149(n117 ,n3[2] ,n22[2]);
    xnor g150(n157 ,n5[0] ,n108);
    nand g151(n385 ,n367 ,n380);
    xnor g152(n343 ,n190 ,n395);
    dff g153(.RN(n1), .SN(1'b1), .CK(n0), .D(n102), .Q(n28[2]));
    dff g154(.RN(n1), .SN(1'b1), .CK(n0), .D(n127), .Q(n20[1]));
    xor g155(n139 ,n24[2] ,n41[2]);
    nor g156(n375 ,n291 ,n373);
    nand g157(n257 ,n28[6] ,n202);
    dff g158(.RN(n1), .SN(1'b1), .CK(n0), .D(n33[1]), .Q(n33[3]));
    xnor g159(n160 ,n8[4] ,n70);
    nand g160(n233 ,n18[0] ,n203);
    nand g161(n394 ,n324 ,n336);
    dff g162(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[3]), .Q(n11[3]));
    nand g163(n213 ,n31[7] ,n207);
    dff g164(.RN(n408), .SN(1'b1), .CK(n0), .D(n400), .Q(n47[4]));
    nand g165(n281 ,n20[3] ,n201);
    xnor g166(n158 ,n8[5] ,n69);
    nand g167(n314 ,n267 ,n285);
    dff g168(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[5]), .Q(n19[7]));
    nand g169(n283 ,n18[1] ,n203);
    xor g170(n156 ,n112 ,n108);
    nor g171(n330 ,n292 ,n290);
    xnor g172(n69 ,n2[10] ,n3[5]);
    dff g173(.RN(n1), .SN(1'b1), .CK(n0), .D(n31[0]), .Q(n31[2]));
    xnor g174(n110 ,n2[2] ,n3[2]);
    nand g175(n232 ,n18[3] ,n203);
    xor g176(n73 ,n3[0] ,n22[0]);
    dff g177(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[3]), .Q(n26[5]));
    nand g178(n299 ,n248 ,n227);
    dff g179(.RN(n1), .SN(1'b1), .CK(n0), .D(n24[0]), .Q(n24[2]));
    xor g180(n72 ,n6[3] ,n36[3]);
    xnor g181(n115 ,n5[2] ,n8[2]);
    nand g182(n305 ,n242 ,n241);
    xnor g183(n67 ,n8[3] ,n35[3]);
    nand g184(n196 ,n35[5] ,n178);
    xor g185(n107 ,n7[2] ,n41[1]);
    dff g186(.RN(n1), .SN(1'b1), .CK(n0), .D(n85), .Q(n41[2]));
    not g187(n52 ,n37[7]);
    nand g188(n266 ,n14[7] ,n205);
    xnor g189(n189 ,n35[3] ,n36[3]);
    xor g190(n82 ,n4[3] ,n42[2]);
    xor g191(n74 ,n6[2] ,n36[2]);
    dff g192(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[2]), .Q(n26[4]));
    xor g193(n129 ,n4[4] ,n43[3]);
    nand g194(n403 ,n375 ,n381);
    nand g195(n222 ,n33[2] ,n206);
    dff g196(.RN(n1), .SN(1'b1), .CK(n0), .D(n24[6]), .Q(n17[6]));
    not g197(n51 ,n37[1]);
    dff g198(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[0]), .Q(n25[2]));
    nand g199(n270 ,n24[6] ,n208);
    nand g200(n300 ,n250 ,n249);
    dff g201(.RN(n1), .SN(1'b1), .CK(n0), .D(n101), .Q(n28[3]));
    nor g202(n60 ,n51 ,n37[0]);
    not g203(n408 ,n407);
    nand g204(n303 ,n216 ,n215);
    dff g205(.RN(n1), .SN(1'b1), .CK(n0), .D(n74), .Q(n36[2]));
    dff g206(.RN(n1), .SN(1'b1), .CK(n0), .D(n168), .Q(n37[1]));
    nand g207(n398 ,n245 ,n337);
    dff g208(.RN(n1), .SN(1'b1), .CK(n0), .D(n142), .Q(n17[3]));
    nor g209(n177 ,n16[3] ,n37[3]);
    xor g210(n76 ,n4[6] ,n45[3]);
    xnor g211(n162 ,n118 ,n29[3]);
    dff g212(.RN(n1), .SN(1'b1), .CK(n0), .D(n391), .Q(n10[6]));
    or g213(n339 ,n306 ,n397);
    nand g214(n360 ,n247 ,n356);
    dff g215(.RN(n408), .SN(1'b1), .CK(n0), .D(n403), .Q(n47[1]));
    xnor g216(n118 ,n3[3] ,n22[3]);
    nor g217(n409 ,n47[4] ,n47[6]);
    dff g218(.RN(n1), .SN(1'b1), .CK(n0), .D(n130), .Q(n18[1]));
    dff g219(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[0]), .Q(n16[2]));
    nor g220(n411 ,n397 ,n403);
    nand g221(n389 ,n335 ,n326);
    nand g222(n217 ,n33[6] ,n206);
    nand g223(n261 ,n16[6] ,n205);
    nand g224(n298 ,n266 ,n244);
    dff g225(.RN(n1), .SN(1'b1), .CK(n0), .D(n31[1]), .Q(n31[3]));
    dff g226(.RN(n1), .SN(1'b1), .CK(n0), .D(n99), .Q(n35[1]));
    or g227(n402 ,n385 ,n387);
    nor g228(n335 ,n316 ,n311);
    xor g229(n154 ,n115 ,n116);
    nand g230(n277 ,n21[3] ,n202);
    dff g231(.RN(n1), .SN(1'b1), .CK(n0), .D(n129), .Q(n43[3]));
    nand g232(n321 ,n283 ,n228);
    dff g233(.RN(n1), .SN(1'b1), .CK(n0), .D(n37[7]), .Q(n37[15]));
    xor g234(n406 ,n38[1] ,n38[0]);
    dff g235(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[1]), .Q(n25[3]));
    nand g236(n390 ,n338 ,n327);
    nand g237(n313 ,n286 ,n221);
    xor g238(n95 ,n4[0] ,n39[1]);
    dff g239(.RN(n1), .SN(1'b1), .CK(n0), .D(n133), .Q(n21[0]));
    dff g240(.RN(n1), .SN(1'b1), .CK(n0), .D(n31[5]), .Q(n31[7]));
    or g241(n372 ,n181 ,n363);
    dff g242(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[2]), .Q(n11[2]));
    nor g243(n63 ,n55 ,n37[9]);
    dff g244(.RN(n1), .SN(1'b1), .CK(n0), .D(n150), .Q(n14[3]));
    nor g245(n324 ,n287 ,n314);
    nor g246(n423 ,n422 ,n421);
    xnor g247(n167 ,n9[0] ,n68);
    dff g248(.RN(n1), .SN(1'b1), .CK(n0), .D(n390), .Q(n10[5]));
    xor g249(n104 ,n33[3] ,n44[3]);
    dff g250(.RN(n1), .SN(1'b1), .CK(n0), .D(n125), .Q(n20[3]));
    xnor g251(n185 ,n32[2] ,n29[2]);
    xnor g252(n68 ,n6[0] ,n36[0]);
    or g253(n358 ,n318 ,n352);
    nand g254(n287 ,n259 ,n254);
    dff g255(.RN(n1), .SN(1'b1), .CK(n0), .D(n132), .Q(n21[1]));
    xnor g256(n170 ,n5[3] ,n111);
    xor g257(n138 ,n2[6] ,n3[6]);
    xnor g258(n184 ,n21[3] ,n22[3]);
    xor g259(n135 ,n26[3] ,n40[3]);
    dff g260(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[1]), .Q(n19[3]));
    xor g261(n84 ,n6[2] ,n41[3]);
    nand g262(n211 ,n34[3] ,n206);
    nand g263(n224 ,n33[3] ,n206);
    dff g264(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[4]), .Q(n26[6]));
    xor g265(n124 ,n26[0] ,n40[0]);
    nand g266(n234 ,n28[3] ,n202);
    nand g267(n273 ,n21[0] ,n202);
    xor g268(n140 ,n3[1] ,n22[1]);
    dff g269(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[4]), .Q(n19[6]));
    dff g270(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[5]), .Q(n24[1]));
    xor g271(n77 ,n7[2] ,n45[2]);
    nand g272(n248 ,n17[2] ,n208);
    nand g273(n295 ,n279 ,n276);
    xnor g274(n112 ,n5[0] ,n8[0]);
    xor g275(n136 ,n2[5] ,n3[5]);
    nand g276(n419 ,n410 ,n409);
    nand g277(n251 ,n20[2] ,n201);
    nand g278(n230 ,n27[3] ,n200);
    nor g279(n206 ,n175 ,n179);
    nand g280(n254 ,n14[1] ,n205);
    nand g281(n393 ,n334 ,n333);
    dff g282(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[1]), .Q(n16[3]));
    nand g283(n278 ,n20[6] ,n201);
    nor g284(n338 ,n310 ,n301);
    dff g285(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[7]), .Q(n27[7]));
    xnor g286(n190 ,n21[2] ,n22[2]);
    not g287(n350 ,n348);
    dff g288(.RN(n1), .SN(1'b1), .CK(n0), .D(n33[2]), .Q(n33[4]));
    dff g289(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[6]), .Q(n14[6]));
    dff g290(.RN(n1), .SN(1'b1), .CK(n0), .D(n82), .Q(n42[2]));
    xor g291(n150 ,n16[3] ,n42[3]);
    dff g292(.RN(n1), .SN(1'b1), .CK(n0), .D(n31[3]), .Q(n31[5]));
    dff g293(.RN(n1), .SN(1'b1), .CK(n0), .D(n173), .Q(n29[3]));
    xnor g294(n66 ,n6[1] ,n36[1]);
    nand g295(n220 ,n34[7] ,n206);
    dff g296(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[7]), .Q(n14[7]));
    dff g297(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[3]), .Q(n19[5]));
    xor g298(n148 ,n29[2] ,n32[2]);
    dff g299(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[4]), .Q(n23[6]));
    nand g300(n279 ,n17[7] ,n208);
    xnor g301(n113 ,n5[1] ,n8[1]);
    dff g302(.RN(n1), .SN(1'b1), .CK(n0), .D(n49), .Q(n38[0]));
    xor g303(n128 ,n19[0] ,n39[0]);
    xor g304(n137 ,n24[1] ,n41[1]);
    dff g305(.RN(n1), .SN(1'b1), .CK(n0), .D(n165), .Q(n22[2]));
    nand g306(n291 ,n237 ,n236);
    xnor g307(n186 ,n21[0] ,n22[0]);
    nand g308(n386 ,n378 ,n383);
    xnor g309(n70 ,n2[8] ,n3[4]);
    nand g310(n317 ,n274 ,n273);
    xor g311(n98 ,n25[3] ,n46[3]);
    xnor g312(n174 ,n164 ,n29[2]);
    xor g313(n81 ,n6[3] ,n42[3]);
    dff g314(.RN(n1), .SN(1'b1), .CK(n0), .D(n73), .Q(n22[0]));
    nor g315(n334 ,n315 ,n323);
    nand g316(n301 ,n214 ,n213);
    nand g317(n264 ,n26[6] ,n203);
    nand g318(n216 ,n34[2] ,n206);
    nor g319(n383 ,n204 ,n377);
    nand g320(n382 ,n205 ,n368);
    dff g321(.RN(n1), .SN(1'b1), .CK(n0), .D(n104), .Q(n34[3]));
    nand g322(n348 ,n201 ,n343);
    xor g323(n106 ,n31[3] ,n43[3]);
    xor g324(n91 ,n8[4] ,n35[4]);
    nand g325(n351 ,n201 ,n344);
    nand g326(n296 ,n257 ,n218);
    nand g327(n364 ,n203 ,n353);
    dff g328(.RN(n1), .SN(1'b1), .CK(n0), .D(n140), .Q(n22[1]));
    not g329(n332 ,n331);
    dff g330(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[1]), .Q(n19[1]));
    nand g331(n226 ,n32[3] ,n206);
    dff g332(.RN(n408), .SN(1'b1), .CK(n0), .D(n423), .Q(n13));
    or g333(n391 ,n296 ,n340);
    nand g334(n164 ,n58 ,n152);
    xnor g335(n165 ,n117 ,n29[2]);
    nand g336(n244 ,n18[7] ,n203);
    nand g337(n219 ,n30[7] ,n207);
    xor g338(n127 ,n19[1] ,n39[1]);
    nand g339(n255 ,n27[6] ,n200);
    nand g340(n181 ,n15[1] ,n175);
    xnor g341(n169 ,n71 ,n32[2]);
    dff g342(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[2]), .Q(n19[4]));
    nand g343(n146 ,n63 ,n65);
    dff g344(.RN(n1), .SN(1'b1), .CK(n0), .D(n395), .Q(n10[2]));
    nand g345(n263 ,n25[6] ,n200);
    dff g346(.RN(n1), .SN(1'b1), .CK(n0), .D(n171), .Q(n37[2]));
    nand g347(n225 ,n31[6] ,n207);
    xor g348(n78 ,n4[5] ,n44[3]);
    or g349(n179 ,n176 ,n15[1]);
    nand g350(n310 ,n262 ,n256);
    dff g351(.RN(n1), .SN(1'b1), .CK(n0), .D(n75), .Q(n46[2]));
    nand g352(n316 ,n263 ,n270);
    dff g353(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[2]), .Q(n23[4]));
    dff g354(.RN(n1), .SN(1'b1), .CK(n0), .D(n33[3]), .Q(n33[5]));
    dff g355(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[4]), .Q(n16[6]));
    nor g356(n201 ,n15[2] ,n178);
    dff g357(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[1]), .Q(n26[3]));
    nor g358(n58 ,n56 ,n37[13]);
    dff g359(.RN(n1), .SN(1'b1), .CK(n0), .D(n139), .Q(n17[2]));
    dff g360(.RN(n1), .SN(1'b1), .CK(n0), .D(n153), .Q(n16[0]));
    nand g361(n249 ,n14[2] ,n205);
    dff g362(.RN(n1), .SN(1'b1), .CK(n0), .D(n37[5]), .Q(n37[13]));
    dff g363(.RN(n1), .SN(1'b1), .CK(n0), .D(n128), .Q(n20[0]));
    dff g364(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[5]), .Q(n23[7]));
    dff g365(.RN(n1), .SN(1'b1), .CK(n0), .D(n96), .Q(n39[0]));
    dff g366(.RN(n1), .SN(1'b1), .CK(n0), .D(n33[7]), .Q(n34[7]));
    xor g367(n100 ,n25[2] ,n46[2]);
    nand g368(n322 ,n229 ,n281);
    xor g369(n83 ,n7[3] ,n42[1]);
    nand g370(n252 ,n27[2] ,n200);
    or g371(n378 ,n195 ,n370);
    not g372(n195 ,n194);
    dff g373(.RN(n1), .SN(1'b1), .CK(n0), .D(n131), .Q(n37[4]));
    nor g374(n325 ,n288 ,n322);
    dff g375(.RN(n1), .SN(1'b1), .CK(n0), .D(n107), .Q(n41[1]));
    xnor g376(n370 ,n185 ,n355);
    dff g377(.RN(n408), .SN(1'b1), .CK(n0), .D(n402), .Q(n47[2]));
    xor g378(n85 ,n4[2] ,n41[2]);
    nand g379(n414 ,n402 ,n404);
    nor g380(n200 ,n176 ,n182);
    xor g381(n80 ,n7[0] ,n43[2]);
    dff g382(.RN(n1), .SN(1'b1), .CK(n0), .D(n126), .Q(n20[2]));
    nand g383(n180 ,n16[3] ,n37[3]);
    xnor g384(n108 ,n2[0] ,n3[0]);
    xnor g385(n168 ,n5[1] ,n122);
    xnor g386(n359 ,n197 ,n341);
    dff g387(.RN(n1), .SN(1'b1), .CK(n0), .D(n389), .Q(n10[4]));
    buf g388(n11[1], 1'b0);
    nand g389(n227 ,n18[2] ,n203);
    dff g390(.RN(n1), .SN(1'b1), .CK(n0), .D(n76), .Q(n45[3]));
    nand g391(n267 ,n23[3] ,n202);
    nor g392(n362 ,n331 ,n354);
    nand g393(n361 ,n247 ,n359);
    xnor g394(n344 ,n184 ,n396);
    nand g395(n401 ,n364 ,n384);
    nand g396(n241 ,n21[2] ,n202);
    dff g397(.RN(n1), .SN(1'b1), .CK(n0), .D(n31[2]), .Q(n31[4]));
    xnor g398(n197 ,n35[1] ,n36[1]);
    xor g399(n97 ,n2[14] ,n3[7]);
    dff g400(.RN(n1), .SN(1'b1), .CK(n0), .D(n87), .Q(n35[5]));
    dff g401(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[15]), .Q(n25[1]));
    dff g402(.RN(n1), .SN(1'b1), .CK(n0), .D(n33[0]), .Q(n33[2]));
    xor g403(n133 ,n5[0] ,n21[0]);
    xnor g404(n188 ,n32[3] ,n29[3]);
    nor g405(n418 ,n415 ,n414);
    xnor g406(n192 ,n35[0] ,n36[0]);
    dff g407(.RN(n1), .SN(1'b1), .CK(n0), .D(n105), .Q(n34[2]));
    nand g408(n292 ,n211 ,n238);
    dff g409(.RN(n1), .SN(1'b1), .CK(n0), .D(n91), .Q(n35[4]));
    dff g410(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[2]), .Q(n25[4]));
    dff g411(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[6]), .Q(n18[6]));
    nand g412(n282 ,n19[7] ,n201);
    nand g413(n256 ,n26[7] ,n203);
    dff g414(.RN(n1), .SN(1'b1), .CK(n0), .D(n37[3]), .Q(n37[11]));
    nor g415(n377 ,n194 ,n371);
    dff g416(.RN(n1), .SN(1'b1), .CK(n0), .D(n24[3]), .Q(n24[5]));
    nand g417(n286 ,n16[2] ,n205);
    xnor g418(n356 ,n192 ,n342);
    xnor g419(n119 ,n5[3] ,n8[3]);
    nand g420(n289 ,n231 ,n282);
    nand g421(n319 ,n277 ,n246);
    nand g422(n240 ,n16[7] ,n205);
    nor g423(n399 ,n15[2] ,n346);
    nand g424(n221 ,n31[2] ,n207);
    nand g425(n258 ,n28[7] ,n202);
    dff g426(.RN(n1), .SN(1'b1), .CK(n0), .D(n135), .Q(n18[3]));
    nand g427(n381 ,n205 ,n369);
    nand g428(n64 ,n37[5] ,n53);
    nor g429(n152 ,n62 ,n146);
    dff g430(.RN(n1), .SN(1'b1), .CK(n0), .D(n147), .Q(n32[3]));
    nand g431(n275 ,n22[3] ,n200);
    nand g432(n260 ,n27[7] ,n200);
    dff g433(.RN(n1), .SN(1'b1), .CK(n0), .D(n37[0]), .Q(n37[8]));
    nand g434(n250 ,n28[2] ,n202);
    dff g435(.RN(n1), .SN(1'b1), .CK(n0), .D(n166), .Q(n36[1]));
    dff g436(.RN(n1), .SN(1'b1), .CK(n0), .D(n72), .Q(n36[3]));
    dff g437(.RN(n1), .SN(1'b1), .CK(n0), .D(n123), .Q(n46[3]));
    nor g438(n417 ,n413 ,n412);
    dff g439(.RN(n1), .SN(1'b1), .CK(n0), .D(n89), .Q(n40[1]));
    dff g440(.RN(n1), .SN(1'b1), .CK(n0), .D(n33[5]), .Q(n33[7]));
    dff g441(.RN(n1), .SN(1'b1), .CK(n0), .D(n106), .Q(n30[3]));
    dff g442(.RN(n1), .SN(1'b1), .CK(n0), .D(n170), .Q(n37[3]));
    xor g443(n105 ,n33[2] ,n44[2]);
    xor g444(n94 ,n2[12] ,n3[6]);
    xor g445(n101 ,n23[3] ,n45[3]);
    nor g446(n205 ,n176 ,n181);
    nand g447(n198 ,n35[4] ,n178);
    not g448(n57 ,n37[10]);
    xor g449(n147 ,n29[3] ,n32[3]);
    xnor g450(n166 ,n9[1] ,n66);
    or g451(n357 ,n305 ,n350);
    xor g452(n90 ,n7[1] ,n40[0]);
    xor g453(n346 ,n196 ,n390);
    dff g454(.RN(n1), .SN(1'b1), .CK(n0), .D(n94), .Q(n23[0]));
    nor g455(n379 ,n362 ,n372);
    dff g456(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[0]), .Q(n23[2]));
    nand g457(n412 ,n47[5] ,n47[7]);
    nand g458(n422 ,n417 ,n418);
    xnor g459(n161 ,n121 ,n32[2]);
    dff g460(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[5]), .Q(n16[7]));
    nand g461(n223 ,n29[2] ,n207);
    xnor g462(n172 ,n67 ,n32[3]);
    dff g463(.RN(n1), .SN(1'b1), .CK(n0), .D(n80), .Q(n43[2]));
    dff g464(.RN(n1), .SN(1'b1), .CK(n0), .D(n37[4]), .Q(n37[12]));
    nand g465(n259 ,n25[3] ,n200);
    dff g466(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[6]), .Q(n20[6]));
    dff g467(.RN(n1), .SN(1'b1), .CK(n0), .D(n100), .Q(n27[2]));
    dff g468(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[3]), .Q(n25[5]));
    nand g469(n297 ,n212 ,n223);
    nand g470(n373 ,n347 ,n361);
    xor g471(n131 ,n2[4] ,n3[4]);
    dff g472(.RN(n1), .SN(1'b1), .CK(n0), .D(n38[1]), .Q(n15[1]));
    nand g473(n209 ,n180 ,n199);
    nor g474(n327 ,n294 ,n289);
    nor g475(n208 ,n15[0] ,n181);
    buf g476(n12[1], 1'b0);
    dff g477(.RN(n408), .SN(1'b1), .CK(n0), .D(n398), .Q(n47[6]));
    nor g478(n333 ,n313 ,n312);
    nand g479(n374 ,n349 ,n360);
    dff g480(.RN(n1), .SN(1'b1), .CK(n0), .D(n98), .Q(n27[3]));
    dff g481(.RN(n408), .SN(1'b1), .CK(n0), .D(n397), .Q(n47[7]));
    nand g482(n265 ,n23[6] ,n202);
    dff g483(.RN(n1), .SN(1'b1), .CK(n0), .D(n37[2]), .Q(n37[10]));
    nand g484(n228 ,n31[3] ,n207);
    nor g485(n416 ,n399 ,n401);
    dff g486(.RN(n1), .SN(1'b1), .CK(n0), .D(n172), .Q(n35[3]));
    dff g487(.RN(n1), .SN(1'b1), .CK(n0), .D(n156), .Q(n19[0]));
    dff g488(.RN(n1), .SN(1'b1), .CK(n0), .D(n405), .Q(n38[2]));
    xnor g489(n114 ,n2[2] ,n3[1]);
    not g490(n49 ,n38[0]);
    nand g491(n293 ,n235 ,n278);
    nand g492(n242 ,n22[2] ,n200);
    dff g493(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[7]), .Q(n16[1]));
    dff g494(.RN(n1), .SN(1'b1), .CK(n0), .D(n33[6]), .Q(n34[6]));
    dff g495(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[0]), .Q(n26[2]));
    dff g496(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[7]), .Q(n20[7]));
    dff g497(.RN(n1), .SN(1'b1), .CK(n0), .D(n143), .Q(n14[1]));
    nor g498(n61 ,n52 ,n37[6]);
    xor g499(n130 ,n26[1] ,n40[1]);
    nand g500(n212 ,n32[2] ,n206);
    dff g501(.RN(n1), .SN(1'b1), .CK(n0), .D(n103), .Q(n35[0]));
    nand g502(n239 ,n24[7] ,n208);
    nand g503(n307 ,n217 ,n253);
    not g504(n175 ,n15[2]);
    dff g505(.RN(n1), .SN(1'b1), .CK(n0), .D(n406), .Q(n38[1]));
    nand g506(n318 ,n275 ,n226);
    xnor g507(n171 ,n5[2] ,n110);
    or g508(n365 ,n319 ,n358);
    not g509(n50 ,n37[3]);
    nand g510(n312 ,n233 ,n272);
    dff g511(.RN(n1), .SN(1'b1), .CK(n0), .D(n93), .Q(n39[2]));
    dff g512(.RN(n1), .SN(1'b1), .CK(n0), .D(n124), .Q(n18[0]));
    xor g513(n142 ,n24[3] ,n41[3]);
    dff g514(.RN(n1), .SN(1'b1), .CK(n0), .D(n24[5]), .Q(n24[7]));
    dff g515(.RN(n1), .SN(1'b1), .CK(n0), .D(n394), .Q(n10[1]));
    nand g516(n308 ,n260 ,n220);
    nand g517(n48 ,n38[1] ,n38[0]);
    nor g518(n203 ,n15[2] ,n179);
    dff g519(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[3]), .Q(n26[1]));
    dff g520(.RN(n1), .SN(1'b1), .CK(n0), .D(n169), .Q(n35[2]));
    nor g521(n59 ,n50 ,n37[2]);
    xnor g522(n341 ,n183 ,n394);
    xnor g523(n191 ,n35[2] ,n36[2]);
    nand g524(n404 ,n376 ,n382);
    dff g525(.RN(n1), .SN(1'b1), .CK(n0), .D(n393), .Q(n10[0]));
    xor g526(n75 ,n7[3] ,n46[2]);
    dff g527(.RN(n1), .SN(1'b1), .CK(n0), .D(n78), .Q(n44[3]));
    dff g528(.RN(n1), .SN(1'b1), .CK(n0), .D(n24[4]), .Q(n24[6]));
    dff g529(.RN(n1), .SN(1'b1), .CK(n0), .D(n148), .Q(n32[2]));
    nand g530(n290 ,n234 ,n232);
    nand g531(n395 ,n329 ,n328);
    dff g532(.RN(n1), .SN(1'b1), .CK(n0), .D(n144), .Q(n14[2]));
    dff g533(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[6]), .Q(n27[6]));
    xnor g534(n355 ,n191 ,n343);
    nand g535(n272 ,n20[0] ,n201);
    xnor g536(n331 ,n188 ,n209);
    buf g537(n11[0], 1'b0);
    not g538(n53 ,n37[4]);
    xnor g539(n405 ,n38[2] ,n48);
    xnor g540(n109 ,n5[3] ,n21[3]);
    dff g541(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[0]), .Q(n19[2]));
    nand g542(n238 ,n17[3] ,n208);
    not g543(n352 ,n351);
    dff g544(.RN(n1), .SN(1'b1), .CK(n0), .D(n37[1]), .Q(n37[9]));
    xor g545(n86 ,n31[2] ,n43[2]);
    not g546(n371 ,n370);
    dff g547(.RN(n1), .SN(1'b1), .CK(n0), .D(n160), .Q(n31[0]));
    xnor g548(n187 ,n16[0] ,n37[0]);
    dff g549(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[6]), .Q(n28[6]));
    xnor g550(n120 ,n2[6] ,n3[3]);
    dff g551(.RN(n1), .SN(1'b1), .CK(n0), .D(n396), .Q(n10[3]));
    nand g552(n210 ,n34[6] ,n206);
    nand g553(n347 ,n201 ,n341);
    dff g554(.RN(n1), .SN(1'b1), .CK(n0), .D(n81), .Q(n42[3]));
    xor g555(n144 ,n16[2] ,n42[2]);
    nand g556(n367 ,n203 ,n355);
    nand g557(n235 ,n18[6] ,n203);
    dff g558(.RN(n408), .SN(1'b1), .CK(n0), .D(n399), .Q(n47[5]));
    dff g559(.RN(n1), .SN(1'b1), .CK(n0), .D(n136), .Q(n37[5]));
    nor g560(n400 ,n15[2] ,n345);
    nor g561(n363 ,n332 ,n353);
    dff g562(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[9]), .Q(n31[1]));
    nor g563(n328 ,n300 ,n299);
    dff g564(.RN(n1), .SN(1'b1), .CK(n0), .D(n33[4]), .Q(n33[6]));
    dff g565(.RN(n1), .SN(1'b1), .CK(n0), .D(n137), .Q(n17[1]));
    dff g566(.RN(n1), .SN(1'b1), .CK(n0), .D(n24[2]), .Q(n24[4]));
endmodule
