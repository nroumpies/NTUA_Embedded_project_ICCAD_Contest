module top (n0, n1, n2, n3);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3;
    wire [15:0] n4;
    wire [7:0] n5;
    wire [7:0] n6;
    wire [3:0] n7;
    wire [31:0] n8;
    wire [63:0] n9;
    wire [3:0] n10;
    wire [3:0] n11;
    wire [7:0] n12;
    wire [7:0] n13;
    wire [15:0] n14;
    wire [15:0] n15;
    wire [3:0] n16;
    wire n17, n18, n19, n20, n21, n22, n23, n24;
    wire n25, n26, n27, n28, n29, n30, n31, n32;
    wire n33, n34, n35, n36, n37, n38, n39, n40;
    wire n41, n42, n43, n44, n45, n46, n47, n48;
    wire n49, n50, n51, n52, n53, n54, n55, n56;
    wire n57, n58, n59, n60, n61, n62, n63, n64;
    wire n65, n66, n67, n68, n69, n70, n71, n72;
    wire n73, n74, n75, n76, n77, n78, n79, n80;
    wire n81, n82, n83, n84, n85, n86, n87, n88;
    wire n89, n90, n91, n92, n93, n94, n95, n96;
    wire n97, n98, n99, n100, n101, n102, n103, n104;
    wire n105, n106, n107, n108, n109, n110, n111, n112;
    wire n113, n114, n115, n116, n117, n118, n119, n120;
    wire n121, n122, n123, n124, n125, n126, n127, n128;
    wire n129, n130, n131, n132, n133, n134, n135, n136;
    wire n137, n138, n139, n140, n141, n142, n143, n144;
    wire n145, n146, n147, n148, n149, n150, n151, n152;
    wire n153, n154, n155, n156, n157, n158, n159, n160;
    wire n161, n162, n163, n164, n165, n166, n167, n168;
    wire n169, n170, n171, n172, n173, n174, n175, n176;
    wire n177, n178, n179, n180, n181, n182, n183, n184;
    wire n185, n186, n187, n188, n189, n190, n191, n192;
    wire n193, n194, n195, n196, n197, n198, n199, n200;
    wire n201, n202, n203, n204, n205, n206, n207, n208;
    wire n209, n210, n211, n212, n213, n214, n215, n216;
    wire n217, n218, n219, n220, n221, n222, n223, n224;
    wire n225, n226, n227, n228, n229, n230, n231, n232;
    wire n233, n234, n235, n236, n237, n238, n239, n240;
    wire n241, n242, n243, n244, n245, n246, n247, n248;
    wire n249, n250, n251, n252, n253, n254, n255, n256;
    wire n257, n258, n259, n260, n261, n262, n263, n264;
    wire n265, n266, n267, n268, n269, n270, n271, n272;
    wire n273, n274, n275, n276, n277, n278, n279, n280;
    wire n281, n282, n283, n284, n285, n286, n287, n288;
    wire n289, n290, n291, n292, n293, n294, n295, n296;
    wire n297, n298, n299, n300, n301, n302, n303, n304;
    wire n305, n306, n307, n308, n309, n310, n311, n312;
    wire n313, n314, n315, n316, n317, n318, n319, n320;
    wire n321, n322, n323, n324, n325, n326, n327, n328;
    wire n329, n330, n331, n332, n333, n334, n335, n336;
    wire n337, n338, n339, n340, n341, n342, n343, n344;
    wire n345, n346, n347, n348, n349, n350, n351, n352;
    wire n353, n354, n355, n356, n357, n358, n359, n360;
    wire n361, n362, n363, n364, n365, n366, n367, n368;
    wire n369, n370, n371, n372, n373, n374, n375, n376;
    wire n377, n378, n379, n380, n381, n382, n383, n384;
    wire n385, n386, n387, n388, n389, n390, n391, n392;
    wire n393, n394, n395, n396;
    or g0(n191 ,n13[0] ,n164);
    nand g1(n385 ,n1 ,n16[0]);
    nand g2(n228 ,n368 ,n165);
    not g3(n138 ,n350);
    nor g4(n244 ,n131 ,n185);
    nor g5(n176 ,n122 ,n336);
    not g6(n146 ,n15[0]);
    nor g7(n304 ,n251 ,n297);
    nand g8(n94 ,n14[1] ,n14[0]);
    buf g9(n3[43], n3[63]);
    buf g10(n3[52], n3[63]);
    dff g11(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n393), .Q(n16[2]));
    xnor g12(n302 ,n278 ,n396);
    dff g13(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n218), .Q(n14[7]));
    not g14(n143 ,n7[0]);
    not g15(n102 ,n101);
    buf g16(n3[36], n3[63]);
    nor g17(n71 ,n62 ,n70);
    xnor g18(n343 ,n14[3] ,n96);
    nand g19(n320 ,n313 ,n316);
    buf g20(n3[18], n3[63]);
    or g21(n21 ,n15[13] ,n15[12]);
    dff g22(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n321), .Q(n9[0]));
    or g23(n42 ,n14[4] ,n41);
    nand g24(n108 ,n14[9] ,n106);
    nand g25(n56 ,n47 ,n52);
    dff g26(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n292), .Q(n7[2]));
    nand g27(n238 ,n364 ,n165);
    buf g28(n3[62], n3[63]);
    nand g29(n226 ,n366 ,n165);
    nor g30(n359 ,n120 ,n118);
    xnor g31(n358 ,n10[2] ,n119);
    not g32(n377 ,n334);
    not g33(n116 ,n115);
    nor g34(n45 ,n37 ,n44);
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n183), .Q(n5[5]));
    xnor g36(n357 ,n10[3] ,n121);
    nor g37(n319 ,n305 ,n315);
    xnor g38(n348 ,n14[8] ,n105);
    nor g39(n271 ,n122 ,n190);
    not g40(n140 ,n13[0]);
    nand g41(n208 ,n15[2] ,n186);
    buf g42(n3[28], n3[63]);
    buf g43(n3[47], n3[63]);
    nand g44(n289 ,n358 ,n268);
    not g45(n389 ,n384);
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n271), .Q(n7[1]));
    nand g47(n361 ,n20 ,n31);
    nor g48(n79 ,n15[9] ,n78);
    nand g49(n266 ,n206 ,n233);
    nor g50(n93 ,n14[1] ,n14[0]);
    nand g51(n332 ,n5[5] ,n331);
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n256), .Q(n15[3]));
    nand g53(n269 ,n1 ,n223);
    buf g54(n3[4], n3[63]);
    nand g55(n173 ,n6[2] ,n337);
    buf g56(n3[55], n3[63]);
    buf g57(n3[40], n3[63]);
    nor g58(n192 ,n339 ,n155);
    buf g59(n3[51], n3[63]);
    nor g60(n378 ,n388 ,n2[0]);
    not g61(n153 ,n5[6]);
    not g62(n337 ,n340);
    xnor g63(n393 ,n390 ,n381);
    nor g64(n353 ,n114 ,n116);
    nand g65(n280 ,n144 ,n268);
    buf g66(n3[34], n3[63]);
    nor g67(n395 ,n380 ,n378);
    nand g68(n285 ,n10[2] ,n270);
    nand g69(n356 ,n58 ,n61);
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n264), .Q(n15[6]));
    nor g71(n291 ,n161 ,n250);
    not g72(n120 ,n119);
    nor g73(n211 ,n134 ,n185);
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n177), .Q(n5[4]));
    buf g75(n3[9], n3[63]);
    nand g76(n290 ,n10[3] ,n270);
    nand g77(n163 ,n339 ,n123);
    xnor g78(n333 ,n329 ,n330);
    nor g79(n309 ,n122 ,n306);
    nor g80(n253 ,n170 ,n192);
    nand g81(n70 ,n15[3] ,n69);
    not g82(n139 ,n351);
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n215), .Q(n14[13]));
    not g84(n95 ,n94);
    nor g85(n220 ,n125 ,n185);
    buf g86(n3[33], n3[63]);
    nand g87(n87 ,n15[13] ,n85);
    xnor g88(n324 ,n11[0] ,n12[0]);
    buf g89(n3[1], n3[63]);
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n275), .Q(n15[14]));
    nand g91(n248 ,n374 ,n165);
    buf g92(n3[53], n3[63]);
    nor g93(n49 ,n15[13] ,n15[12]);
    nand g94(n274 ,n241 ,n236);
    not g95(n170 ,n169);
    nor g96(n160 ,n143 ,n122);
    nor g97(n372 ,n72 ,n74);
    nand g98(n310 ,n283 ,n307);
    buf g99(n3[49], n3[63]);
    nand g100(n259 ,n219 ,n226);
    nand g101(n260 ,n199 ,n227);
    nor g102(n161 ,n142 ,n6[0]);
    nand g103(n383 ,n390 ,n382);
    nand g104(n40 ,n33 ,n34);
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n300), .Q(n10[1]));
    buf g106(n3[50], n3[63]);
    nand g107(n275 ,n240 ,n237);
    xnor g108(n370 ,n15[7] ,n75);
    not g109(n91 ,n14[8]);
    nand g110(n219 ,n15[11] ,n186);
    not g111(n28 ,n27);
    nor g112(n215 ,n128 ,n185);
    buf g113(n3[17], n3[63]);
    buf g114(n3[37], n3[63]);
    nor g115(n247 ,n136 ,n185);
    nand g116(n276 ,n225 ,n238);
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n220), .Q(n14[5]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n214), .Q(n14[11]));
    or g119(n322 ,n6[2] ,n5[4]);
    xnor g120(n362 ,n89 ,n15[15]);
    not g121(n128 ,n353);
    nand g122(n205 ,n15[5] ,n186);
    buf g123(n3[21], n3[63]);
    not g124(n184 ,n185);
    nand g125(n267 ,n10[3] ,n197);
    not g126(n270 ,n269);
    nor g127(n57 ,n15[2] ,n56);
    not g128(n32 ,n14[3]);
    nand g129(n241 ,n15[15] ,n186);
    buf g130(n3[48], n3[63]);
    buf g131(n3[44], n3[63]);
    not g132(n81 ,n80);
    nand g133(n96 ,n14[2] ,n95);
    nor g134(n179 ,n151 ,n122);
    buf g135(n3[26], n3[63]);
    nand g136(n239 ,n365 ,n165);
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n244), .Q(n14[6]));
    nand g138(n73 ,n15[5] ,n71);
    nor g139(n35 ,n14[15] ,n14[14]);
    nand g140(n286 ,n10[1] ,n270);
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n272), .Q(n15[1]));
    buf g142(n3[22], n3[63]);
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n265), .Q(n15[5]));
    xnor g144(n350 ,n14[10] ,n108);
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n176), .Q(n4[0]));
    xnor g146(n363 ,n15[14] ,n87);
    buf g147(n3[0], n3[63]);
    xnor g148(n329 ,n326 ,n323);
    or g149(n297 ,n13[2] ,n281);
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n394), .Q(n16[1]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n274), .Q(n15[15]));
    nor g152(n183 ,n150 ,n122);
    nand g153(n159 ,n7[0] ,n10[0]);
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n212), .Q(n14[15]));
    nand g155(n210 ,n15[0] ,n186);
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n261), .Q(n15[9]));
    buf g157(n3[14], n3[63]);
    nand g158(n29 ,n15[5] ,n28);
    nor g159(n106 ,n91 ,n105);
    not g160(n97 ,n96);
    nand g161(n312 ,n13[0] ,n309);
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n296), .Q(n10[0]));
    buf g163(n3[54], n3[63]);
    not g164(n90 ,n14[4]);
    xnor g165(n190 ,n13[0] ,n13[1]);
    nor g166(n169 ,n7[0] ,n7[2]);
    not g167(n132 ,n355);
    nor g168(n224 ,n7[3] ,n169);
    nand g169(n360 ,n35 ,n46);
    nor g170(n86 ,n15[13] ,n85);
    xnor g171(n351 ,n14[11] ,n110);
    nor g172(n50 ,n15[7] ,n15[6]);
    nand g173(n256 ,n207 ,n248);
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n392), .Q(n396));
    nand g175(n112 ,n14[11] ,n111);
    nand g176(n250 ,n156 ,n224);
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n263), .Q(n15[7]));
    buf g178(n3[39], n3[63]);
    nor g179(n107 ,n14[9] ,n106);
    nand g180(n207 ,n15[3] ,n186);
    nand g181(n278 ,n154 ,n257);
    nand g182(n66 ,n15[1] ,n15[0]);
    nand g183(n308 ,n171 ,n306);
    nand g184(n237 ,n363 ,n165);
    nor g185(n198 ,n13[2] ,n167);
    xnor g186(n338 ,n4[0] ,n339);
    nand g187(n257 ,n159 ,n196);
    not g188(n104 ,n103);
    not g189(n142 ,n7[2]);
    nand g190(n121 ,n10[2] ,n120);
    not g191(n111 ,n110);
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n189), .Q(n14[0]));
    buf g193(n3[15], n3[63]);
    xnor g194(n355 ,n117 ,n14[15]);
    or g195(n195 ,n187 ,n168);
    nand g196(n223 ,n13[2] ,n167);
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n317), .Q(n13[0]));
    nor g198(n51 ,n15[11] ,n15[10]);
    buf g199(n3[10], n3[63]);
    nand g200(n200 ,n15[9] ,n186);
    nand g201(n52 ,n15[1] ,n15[0]);
    nor g202(n318 ,n304 ,n311);
    buf g203(n3[27], n3[63]);
    not g204(n145 ,n6[0]);
    nor g205(n175 ,n152 ,n122);
    nor g206(n114 ,n14[13] ,n113);
    not g207(n67 ,n66);
    nand g208(n236 ,n362 ,n165);
    buf g209(n3[31], n3[63]);
    not g210(n92 ,n14[12]);
    nand g211(n234 ,n375 ,n165);
    buf g212(n3[20], n3[63]);
    buf g213(n3[5], n3[63]);
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n318), .Q(n13[2]));
    nor g215(n58 ,n15[15] ,n55);
    nor g216(n197 ,n144 ,n168);
    xnor g217(n325 ,n9[0] ,n10[0]);
    nand g218(n313 ,n13[1] ,n309);
    nand g219(n43 ,n14[9] ,n42);
    nand g220(n119 ,n10[1] ,n10[0]);
    nor g221(n303 ,n279 ,n294);
    buf g222(n3[60], n3[63]);
    nor g223(n281 ,n13[0] ,n254);
    nand g224(n288 ,n357 ,n268);
    nor g225(n204 ,n129 ,n185);
    xnor g226(n367 ,n15[10] ,n80);
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n262), .Q(n15[8]));
    nor g228(n46 ,n40 ,n45);
    nand g229(n115 ,n14[13] ,n113);
    not g230(n151 ,n6[1]);
    not g231(n74 ,n73);
    nor g232(n311 ,n292 ,n309);
    nand g233(n68 ,n15[2] ,n67);
    not g234(n152 ,n5[5]);
    nor g235(n18 ,n15[15] ,n15[14]);
    buf g236(n3[30], n3[63]);
    not g237(n122 ,n1);
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n213), .Q(n14[14]));
    buf g239(n3[11], n3[63]);
    xnor g240(n347 ,n14[7] ,n103);
    xnor g241(n365 ,n15[12] ,n84);
    nand g242(n166 ,n13[0] ,n13[1]);
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n180), .Q(n6[1]));
    nor g244(n65 ,n15[1] ,n15[0]);
    nand g245(n225 ,n15[13] ,n186);
    nand g246(n27 ,n15[6] ,n26);
    nor g247(n33 ,n14[13] ,n14[12]);
    xnor g248(n392 ,n391 ,n383);
    nor g249(n213 ,n133 ,n185);
    not g250(n150 ,n5[4]);
    xnor g251(n323 ,n13[0] ,n14[0]);
    nor g252(n158 ,n122 ,n123);
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n259), .Q(n15[11]));
    nor g254(n180 ,n145 ,n122);
    nor g255(n254 ,n162 ,n193);
    not g256(n125 ,n345);
    nand g257(n105 ,n14[7] ,n104);
    buf g258(n3[8], n3[63]);
    not g259(n129 ,n348);
    nor g260(n118 ,n10[1] ,n10[0]);
    nand g261(n24 ,n15[2] ,n17);
    not g262(n148 ,n7[3]);
    nand g263(n98 ,n14[3] ,n97);
    nor g264(n212 ,n132 ,n185);
    nor g265(n293 ,n396 ,n291);
    or g266(n60 ,n54 ,n59);
    nand g267(n55 ,n49 ,n51);
    or g268(n17 ,n15[1] ,n15[0]);
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n266), .Q(n15[4]));
    nor g270(n100 ,n14[5] ,n99);
    nand g271(n77 ,n15[7] ,n76);
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n249), .Q(n11[0]));
    nor g273(n20 ,n15[9] ,n15[8]);
    dff g274(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n243), .Q(n14[1]));
    buf g275(n3[2], n3[63]);
    nor g276(n321 ,n122 ,n319);
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n320), .Q(n13[1]));
    not g278(n76 ,n75);
    buf g279(n3[35], n3[63]);
    nand g280(n82 ,n15[10] ,n81);
    nor g281(n188 ,n166 ,n187);
    nor g282(n376 ,n67 ,n65);
    xnor g283(n330 ,n324 ,n325);
    xnor g284(n373 ,n15[4] ,n70);
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n204), .Q(n14[8]));
    nand g286(n298 ,n290 ,n288);
    nor g287(n99 ,n90 ,n98);
    nor g288(n246 ,n127 ,n185);
    nand g289(n53 ,n15[5] ,n15[4]);
    nor g290(n61 ,n15[14] ,n60);
    nand g291(n201 ,n15[8] ,n186);
    nand g292(n299 ,n285 ,n289);
    or g293(n44 ,n38 ,n43);
    not g294(n141 ,n13[1]);
    nand g295(n381 ,n389 ,n380);
    dff g296(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n298), .Q(n10[3]));
    nor g297(n59 ,n53 ,n57);
    nor g298(n177 ,n149 ,n122);
    nand g299(n185 ,n1 ,n2[0]);
    not g300(n149 ,n5[3]);
    xnor g301(n369 ,n15[8] ,n77);
    nand g302(n379 ,n388 ,n2[0]);
    nand g303(n38 ,n14[8] ,n14[5]);
    buf g304(n3[45], n3[63]);
    dff g305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n246), .Q(n14[2]));
    nor g306(n165 ,n122 ,n377);
    nor g307(n334 ,n322 ,n332);
    not g308(n137 ,n344);
    buf g309(n3[13], n3[63]);
    nand g310(n181 ,n6[0] ,n13[1]);
    nand g311(n384 ,n1 ,n16[1]);
    nor g312(n171 ,n122 ,n13[0]);
    nand g313(n386 ,n1 ,n16[2]);
    buf g314(n3[41], n3[63]);
    buf g315(n3[42], n3[63]);
    dff g316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n158), .Q(n8[0]));
    buf g317(n3[56], n3[63]);
    nor g318(n279 ,n172 ,n267);
    nor g319(n193 ,n181 ,n173);
    not g320(n336 ,n338);
    nand g321(n182 ,n7[1] ,n148);
    dff g322(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n175), .Q(n5[6]));
    nand g323(n261 ,n200 ,n228);
    not g324(n380 ,n379);
    nand g325(n283 ,n163 ,n253);
    not g326(n167 ,n166);
    nand g327(n242 ,n15[12] ,n186);
    nand g328(n101 ,n14[5] ,n99);
    buf g329(n3[46], n3[63]);
    nor g330(n364 ,n86 ,n88);
    buf g331(n3[58], n3[63]);
    xnor g332(n371 ,n15[6] ,n73);
    nor g333(n221 ,n137 ,n185);
    nor g334(n31 ,n15[7] ,n30);
    xnor g335(n352 ,n14[12] ,n112);
    nand g336(n231 ,n371 ,n165);
    nor g337(n306 ,n304 ,n303);
    nand g338(n262 ,n201 ,n229);
    nand g339(n255 ,n210 ,n194);
    dff g340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n268), .Q(n7[3]));
    xnor g341(n374 ,n15[3] ,n68);
    nand g342(n387 ,n1 ,n396);
    nand g343(n110 ,n14[10] ,n109);
    nor g344(n292 ,n198 ,n269);
    nor g345(n214 ,n139 ,n185);
    xnor g346(n354 ,n14[14] ,n115);
    buf g347(n3[7], n3[63]);
    nor g348(n174 ,n153 ,n122);
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n211), .Q(n14[9]));
    nand g350(n282 ,n10[0] ,n270);
    nand g351(n265 ,n205 ,n232);
    not g352(n135 ,n352);
    nor g353(n162 ,n335 ,n13[1]);
    nand g354(n80 ,n15[9] ,n78);
    nor g355(n196 ,n142 ,n157);
    or g356(n156 ,n7[2] ,n2[0]);
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n174), .Q(n5[7]));
    nand g358(n84 ,n15[11] ,n83);
    nand g359(n300 ,n286 ,n284);
    nand g360(n316 ,n271 ,n312);
    dff g361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n260), .Q(n15[10]));
    not g362(n124 ,n377);
    dff g363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n276), .Q(n15[13]));
    nand g364(n273 ,n2[0] ,n188);
    nor g365(n218 ,n126 ,n185);
    dff g366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n277), .Q(n15[2]));
    nand g367(n194 ,n146 ,n165);
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n160), .Q(n12[0]));
    nand g369(n75 ,n15[6] ,n74);
    nand g370(n263 ,n202 ,n230);
    dff g371(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n247), .Q(n14[3]));
    nand g372(n307 ,n224 ,n302);
    nand g373(n251 ,n245 ,n195);
    not g374(n133 ,n354);
    nand g375(n301 ,n182 ,n295);
    nand g376(n339 ,n356 ,n334);
    not g377(n64 ,n15[12]);
    dff g378(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n179), .Q(n6[2]));
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n171), .Q(n7[0]));
    nor g380(n39 ,n14[1] ,n36);
    nand g381(n245 ,n360 ,n167);
    nor g382(n368 ,n79 ,n81);
    nor g383(n34 ,n14[11] ,n14[10]);
    buf g384(n3[59], n3[63]);
    not g385(n131 ,n346);
    nor g386(n252 ,n377 ,n191);
    xnor g387(n344 ,n14[4] ,n98);
    nand g388(n54 ,n48 ,n50);
    dff g389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n184), .Q(n6[0]));
    nor g390(n22 ,n15[11] ,n15[10]);
    buf g391(n3[16], n3[63]);
    buf g392(n3[19], n3[63]);
    nand g393(n187 ,n2[2] ,n2[1]);
    or g394(n154 ,n14[0] ,n7[2]);
    nand g395(n264 ,n203 ,n231);
    not g396(n47 ,n15[3]);
    nor g397(n249 ,n122 ,n222);
    nor g398(n113 ,n92 ,n112);
    dff g399(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n178), .Q(n5[3]));
    nor g400(n349 ,n107 ,n109);
    not g401(n382 ,n381);
    nor g402(n78 ,n63 ,n77);
    not g403(n126 ,n347);
    xnor g404(n326 ,n7[0] ,n8[0]);
    not g405(n130 ,n341);
    nand g406(n296 ,n282 ,n280);
    xnor g407(n346 ,n14[6] ,n101);
    not g408(n109 ,n108);
    xnor g409(n342 ,n14[2] ,n94);
    buf g410(n3[57], n3[63]);
    nor g411(n189 ,n14[0] ,n185);
    nor g412(n268 ,n122 ,n223);
    not g413(n388 ,n385);
    not g414(n62 ,n15[4]);
    nand g415(n209 ,n15[1] ,n186);
    not g416(n134 ,n349);
    nor g417(n164 ,n141 ,n356);
    nand g418(n272 ,n209 ,n235);
    nand g419(n277 ,n208 ,n234);
    not g420(n335 ,n361);
    nor g421(n341 ,n95 ,n93);
    xnor g422(n366 ,n15[11] ,n82);
    dff g423(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n258), .Q(n15[12]));
    buf g424(n3[6], n3[63]);
    nand g425(n26 ,n19 ,n24);
    nor g426(n186 ,n122 ,n124);
    nor g427(n25 ,n21 ,n23);
    nand g428(n232 ,n372 ,n165);
    not g429(n144 ,n10[0]);
    nand g430(n230 ,n370 ,n165);
    or g431(n36 ,n14[2] ,n14[0]);
    not g432(n127 ,n342);
    nand g433(n233 ,n373 ,n165);
    nor g434(n243 ,n130 ,n185);
    nand g435(n103 ,n14[6] ,n102);
    dff g436(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n216), .Q(n14[12]));
    xnor g437(n394 ,n389 ,n379);
    nor g438(n305 ,n293 ,n301);
    xnor g439(n375 ,n15[2] ,n66);
    buf g440(n3[25], n3[63]);
    nand g441(n340 ,n5[3] ,n6[1]);
    dff g442(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n299), .Q(n10[2]));
    nand g443(n117 ,n14[14] ,n116);
    not g444(n391 ,n387);
    nand g445(n229 ,n369 ,n165);
    nor g446(n157 ,n140 ,n7[0]);
    not g447(n83 ,n82);
    nand g448(n30 ,n25 ,n29);
    nand g449(n284 ,n359 ,n268);
    or g450(n294 ,n252 ,n287);
    nand g451(n172 ,n10[1] ,n10[2]);
    nand g452(n168 ,n13[0] ,n141);
    nand g453(n314 ,n7[1] ,n310);
    xnor g454(n222 ,n396 ,n11[0]);
    dff g455(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n395), .Q(n16[0]));
    not g456(n136 ,n343);
    not g457(n147 ,n6[2]);
    nand g458(n287 ,n13[2] ,n273);
    not g459(n390 ,n386);
    nor g460(n345 ,n100 ,n102);
    not g461(n63 ,n15[8]);
    buf g462(n3[29], n3[63]);
    buf g463(n3[23], n3[63]);
    dff g464(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n221), .Q(n14[4]));
    nor g465(n41 ,n32 ,n39);
    not g466(n315 ,n314);
    nand g467(n295 ,n396 ,n291);
    nor g468(n331 ,n6[0] ,n328);
    nor g469(n327 ,n5[6] ,n340);
    nand g470(n23 ,n18 ,n22);
    nor g471(n178 ,n147 ,n122);
    buf g472(n3[24], n3[63]);
    xnor g473(n3[63] ,n338 ,n333);
    nand g474(n258 ,n242 ,n239);
    nor g475(n72 ,n15[5] ,n71);
    nor g476(n155 ,n7[3] ,n396);
    nand g477(n227 ,n367 ,n165);
    buf g478(n3[61], n3[63]);
    buf g479(n3[3], n3[63]);
    nor g480(n19 ,n15[4] ,n15[3]);
    dff g481(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n217), .Q(n14[10]));
    nor g482(n48 ,n15[9] ,n15[8]);
    nand g483(n317 ,n312 ,n308);
    not g484(n123 ,n396);
    buf g485(n3[12], n3[63]);
    nor g486(n85 ,n64 ,n84);
    buf g487(n3[32], n3[63]);
    nand g488(n202 ,n15[7] ,n186);
    nand g489(n203 ,n15[6] ,n186);
    buf g490(n3[38], n3[63]);
    not g491(n69 ,n68);
    nor g492(n217 ,n138 ,n185);
    nand g493(n235 ,n376 ,n165);
    nand g494(n328 ,n5[7] ,n327);
    nand g495(n89 ,n15[14] ,n88);
    nor g496(n216 ,n135 ,n185);
    nand g497(n240 ,n15[14] ,n186);
    nand g498(n199 ,n15[10] ,n186);
    not g499(n88 ,n87);
    dff g500(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n255), .Q(n15[0]));
    nand g501(n206 ,n15[4] ,n186);
    nand g502(n37 ,n14[7] ,n14[6]);
endmodule
