module top (n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [3:0] n6;
    wire [31:0] n7;
    wire [31:0] n8;
    wire [1:0] n9;
    wire [31:0] n10;
    wire n11, n12, n13, n14, n15, n16, n17, n18;
    wire n19, n20, n21, n22, n23, n24, n25, n26;
    wire n27, n28, n29, n30, n31, n32, n33, n34;
    wire n35, n36, n37, n38, n39, n40, n41, n42;
    wire n43, n44, n45, n46, n47, n48, n49, n50;
    wire n51, n52, n53, n54, n55, n56, n57, n58;
    wire n59, n60, n61, n62, n63, n64, n65, n66;
    wire n67, n68, n69, n70, n71, n72, n73, n74;
    wire n75, n76, n77, n78, n79, n80, n81, n82;
    wire n83, n84, n85, n86, n87, n88, n89, n90;
    wire n91, n92, n93, n94, n95, n96, n97, n98;
    wire n99, n100, n101, n102, n103, n104, n105, n106;
    wire n107, n108, n109, n110, n111, n112, n113, n114;
    wire n115, n116, n117, n118, n119, n120, n121, n122;
    wire n123, n124, n125, n126, n127, n128, n129, n130;
    wire n131, n132, n133, n134, n135, n136, n137, n138;
    wire n139, n140, n141, n142, n143, n144, n145, n146;
    wire n147, n148, n149, n150, n151, n152, n153, n154;
    wire n155, n156, n157, n158, n159, n160, n161, n162;
    wire n163, n164, n165, n166, n167, n168, n169, n170;
    wire n171, n172, n173, n174, n175, n176, n177, n178;
    wire n179, n180, n181, n182, n183, n184, n185, n186;
    wire n187, n188, n189, n190, n191, n192, n193, n194;
    wire n195, n196, n197, n198, n199, n200, n201, n202;
    wire n203, n204, n205, n206, n207, n208, n209, n210;
    wire n211, n212, n213, n214, n215, n216, n217, n218;
    wire n219, n220, n221, n222, n223, n224, n225, n226;
    wire n227, n228, n229, n230, n231, n232, n233, n234;
    wire n235, n236, n237, n238, n239, n240, n241, n242;
    wire n243, n244, n245, n246, n247, n248, n249, n250;
    wire n251, n252, n253, n254, n255, n256, n257, n258;
    wire n259, n260, n261, n262, n263, n264, n265, n266;
    wire n267, n268, n269, n270, n271, n272, n273, n274;
    wire n275, n276, n277, n278, n279, n280, n281, n282;
    wire n283, n284, n285, n286, n287, n288, n289, n290;
    wire n291, n292, n293, n294, n295, n296, n297, n298;
    wire n299, n300, n301, n302, n303, n304, n305, n306;
    wire n307, n308, n309, n310, n311, n312, n313, n314;
    wire n315, n316, n317, n318, n319, n320, n321, n322;
    wire n323, n324, n325, n326, n327, n328, n329, n330;
    wire n331, n332, n333, n334, n335, n336, n337, n338;
    wire n339, n340, n341, n342, n343, n344, n345, n346;
    wire n347, n348, n349, n350, n351, n352, n353, n354;
    wire n355, n356, n357, n358, n359, n360, n361, n362;
    wire n363, n364, n365, n366, n367, n368, n369, n370;
    wire n371, n372, n373, n374, n375, n376, n377, n378;
    wire n379, n380, n381, n382, n383, n384, n385, n386;
    wire n387, n388, n389, n390, n391, n392, n393, n394;
    wire n395, n396, n397, n398, n399, n400, n401, n402;
    wire n403, n404, n405, n406, n407, n408, n409, n410;
    wire n411, n412, n413, n414, n415, n416, n417, n418;
    wire n419, n420, n421, n422, n423, n424, n425, n426;
    wire n427, n428, n429, n430, n431, n432, n433, n434;
    wire n435, n436, n437, n438, n439, n440, n441, n442;
    wire n443, n444, n445, n446, n447, n448, n449, n450;
    wire n451, n452, n453, n454, n455, n456, n457, n458;
    wire n459, n460, n461, n462, n463, n464, n465, n466;
    wire n467, n468, n469, n470, n471, n472, n473, n474;
    wire n475, n476, n477, n478, n479, n480, n481, n482;
    wire n483, n484, n485, n486, n487, n488, n489, n490;
    wire n491, n492, n493, n494, n495, n496, n497, n498;
    wire n499, n500, n501, n502, n503, n504, n505, n506;
    wire n507, n508, n509, n510, n511, n512, n513, n514;
    wire n515, n516, n517, n518, n519, n520, n521, n522;
    wire n523, n524, n525, n526, n527, n528, n529, n530;
    wire n531, n532, n533, n534, n535, n536, n537, n538;
    wire n539, n540, n541, n542, n543, n544, n545, n546;
    wire n547, n548, n549, n550, n551, n552, n553, n554;
    wire n555, n556, n557, n558, n559, n560, n561, n562;
    wire n563, n564, n565, n566, n567, n568, n569, n570;
    wire n571, n572, n573, n574, n575, n576, n577, n578;
    wire n579, n580, n581, n582, n583, n584, n585, n586;
    wire n587, n588, n589, n590, n591, n592, n593, n594;
    wire n595, n596, n597, n598, n599, n600, n601, n602;
    wire n603, n604, n605, n606, n607, n608, n609, n610;
    wire n611, n612, n613, n614, n615, n616, n617, n618;
    wire n619, n620, n621, n622, n623, n624, n625, n626;
    wire n627, n628, n629, n630, n631, n632, n633, n634;
    wire n635, n636, n637, n638, n639, n640, n641, n642;
    wire n643, n644, n645, n646, n647, n648, n649, n650;
    wire n651, n652, n653, n654, n655, n656, n657, n658;
    wire n659, n660, n661, n662, n663, n664, n665, n666;
    wire n667, n668, n669, n670, n671, n672, n673, n674;
    wire n675, n676, n677, n678, n679, n680, n681, n682;
    wire n683, n684, n685, n686, n687, n688, n689, n690;
    wire n691, n692, n693, n694, n695, n696, n697, n698;
    wire n699, n700, n701, n702, n703, n704, n705, n706;
    wire n707, n708, n709, n710, n711, n712, n713, n714;
    wire n715, n716, n717, n718, n719, n720, n721, n722;
    wire n723, n724, n725, n726, n727, n728, n729, n730;
    wire n731, n732, n733, n734, n735, n736, n737, n738;
    wire n739, n740, n741, n742, n743, n744, n745, n746;
    wire n747, n748, n749, n750, n751, n752, n753, n754;
    wire n755, n756, n757, n758, n759, n760, n761, n762;
    wire n763, n764, n765, n766, n767, n768, n769, n770;
    wire n771, n772, n773, n774, n775, n776, n777, n778;
    wire n779, n780, n781, n782, n783, n784, n785, n786;
    wire n787, n788, n789, n790, n791, n792, n793, n794;
    wire n795, n796, n797, n798, n799, n800, n801, n802;
    wire n803, n804, n805, n806, n807, n808, n809, n810;
    wire n811, n812, n813, n814, n815, n816, n817, n818;
    wire n819, n820, n821, n822, n823, n824, n825, n826;
    wire n827, n828, n829, n830, n831, n832, n833, n834;
    wire n835, n836, n837, n838, n839, n840, n841, n842;
    wire n843, n844, n845, n846, n847, n848, n849, n850;
    wire n851, n852, n853, n854, n855, n856, n857, n858;
    wire n859, n860, n861, n862, n863, n864, n865, n866;
    wire n867, n868, n869, n870, n871, n872, n873, n874;
    wire n875, n876, n877, n878, n879, n880, n881, n882;
    wire n883, n884, n885, n886, n887, n888, n889, n890;
    wire n891, n892, n893, n894, n895, n896, n897, n898;
    wire n899, n900, n901, n902, n903, n904, n905, n906;
    wire n907, n908, n909, n910, n911, n912, n913, n914;
    wire n915, n916, n917, n918, n919, n920, n921, n922;
    wire n923, n924, n925, n926, n927, n928, n929, n930;
    wire n931, n932, n933, n934, n935, n936, n937, n938;
    wire n939, n940, n941, n942, n943, n944, n945, n946;
    wire n947, n948, n949, n950, n951, n952, n953, n954;
    wire n955, n956, n957, n958, n959, n960, n961, n962;
    wire n963, n964, n965, n966, n967, n968, n969, n970;
    wire n971, n972, n973, n974, n975, n976, n977, n978;
    wire n979, n980, n981, n982, n983, n984, n985, n986;
    wire n987, n988, n989, n990, n991, n992, n993, n994;
    wire n995, n996, n997, n998, n999, n1000, n1001, n1002;
    wire n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010;
    wire n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018;
    wire n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
    wire n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
    wire n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
    wire n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050;
    wire n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058;
    wire n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066;
    wire n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074;
    wire n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082;
    wire n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090;
    wire n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098;
    wire n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106;
    wire n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114;
    wire n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122;
    wire n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130;
    wire n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138;
    wire n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146;
    wire n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154;
    wire n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162;
    wire n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170;
    wire n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178;
    wire n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186;
    wire n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194;
    wire n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202;
    wire n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210;
    wire n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218;
    wire n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226;
    wire n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234;
    wire n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242;
    wire n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250;
    wire n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258;
    wire n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266;
    wire n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274;
    wire n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282;
    wire n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290;
    wire n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298;
    wire n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306;
    wire n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314;
    wire n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322;
    wire n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330;
    wire n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338;
    wire n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346;
    wire n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354;
    wire n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362;
    wire n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370;
    wire n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378;
    wire n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386;
    wire n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394;
    wire n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402;
    wire n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410;
    wire n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418;
    wire n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426;
    wire n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434;
    wire n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442;
    wire n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450;
    wire n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458;
    wire n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466;
    wire n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474;
    wire n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482;
    wire n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490;
    wire n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498;
    wire n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506;
    wire n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514;
    wire n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522;
    wire n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530;
    wire n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538;
    wire n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546;
    wire n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554;
    wire n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562;
    wire n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570;
    wire n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578;
    wire n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586;
    wire n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594;
    wire n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602;
    wire n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610;
    wire n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618;
    wire n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626;
    wire n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634;
    wire n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642;
    wire n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650;
    wire n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658;
    wire n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666;
    wire n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674;
    wire n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682;
    wire n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690;
    wire n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698;
    wire n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706;
    wire n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714;
    wire n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722;
    wire n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730;
    wire n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738;
    wire n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746;
    wire n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754;
    wire n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762;
    wire n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770;
    wire n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778;
    wire n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786;
    wire n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794;
    wire n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802;
    wire n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810;
    wire n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818;
    wire n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826;
    wire n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834;
    wire n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842;
    wire n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850;
    wire n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858;
    wire n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866;
    wire n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874;
    wire n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882;
    wire n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890;
    wire n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898;
    wire n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906;
    wire n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914;
    wire n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922;
    wire n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930;
    wire n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938;
    wire n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946;
    wire n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954;
    wire n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962;
    wire n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970;
    wire n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978;
    wire n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986;
    wire n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994;
    wire n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002;
    wire n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010;
    wire n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018;
    wire n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026;
    wire n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034;
    wire n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042;
    wire n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050;
    wire n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058;
    wire n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066;
    wire n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074;
    wire n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082;
    wire n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090;
    wire n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098;
    wire n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106;
    wire n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114;
    wire n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122;
    wire n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130;
    wire n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138;
    wire n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146;
    wire n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154;
    wire n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162;
    wire n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170;
    wire n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178;
    wire n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186;
    wire n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194;
    wire n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202;
    wire n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210;
    wire n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218;
    wire n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226;
    wire n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234;
    wire n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242;
    wire n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250;
    wire n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258;
    wire n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266;
    wire n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274;
    wire n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282;
    wire n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290;
    wire n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298;
    wire n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306;
    wire n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314;
    wire n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322;
    wire n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330;
    wire n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338;
    wire n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346;
    wire n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354;
    wire n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362;
    wire n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370;
    wire n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378;
    wire n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386;
    wire n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394;
    wire n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402;
    wire n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410;
    wire n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418;
    wire n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426;
    wire n2427, n2428, n2429;
    nor g0(n948 ,n492 ,n875);
    nor g1(n1338 ,n5[4] ,n1040);
    nand g2(n630 ,n8[4] ,n2359);
    nor g3(n1766 ,n1352 ,n1260);
    nand g4(n1943 ,n5[15] ,n1631);
    nor g5(n958 ,n373 ,n875);
    nand g6(n2101 ,n1974 ,n1973);
    nor g7(n185 ,n39 ,n184);
    not g8(n1692 ,n1607);
    nand g9(n2074 ,n1741 ,n1739);
    dff g10(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2284), .Q(n3[6]));
    nand g11(n2426 ,n2424 ,n2425);
    nand g12(n1741 ,n4[21] ,n1462);
    xnor g13(n2353 ,n80 ,n195);
    nor g14(n838 ,n526 ,n804);
    dff g15(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2161), .Q(n5[26]));
    nand g16(n1625 ,n756 ,n948);
    not g17(n1259 ,n1131);
    nand g18(n1744 ,n4[20] ,n1464);
    nand g19(n2213 ,n3[45] ,n1878);
    or g20(n1484 ,n810 ,n1046);
    dff g21(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2123), .Q(n4[36]));
    nor g22(n1400 ,n4[52] ,n1024);
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2308), .Q(n3[50]));
    nor g24(n1853 ,n1384 ,n1217);
    nor g25(n410 ,n8[9] ,n2[41]);
    nor g26(n1792 ,n1363 ,n1672);
    nor g27(n1973 ,n1518 ,n1684);
    nand g28(n2149 ,n1801 ,n1797);
    or g29(n1477 ,n807 ,n1065);
    not g30(n1326 ,n1198);
    nor g31(n450 ,n8[23] ,n2[23]);
    xnor g32(n2372 ,n98 ,n233);
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2292), .Q(n3[34]));
    nor g34(n918 ,n449 ,n804);
    nor g35(n1330 ,n3[23] ,n1028);
    nor g36(n908 ,n476 ,n804);
    nor g37(n42 ,n2[9] ,n2[73]);
    nand g38(n2311 ,n1836 ,n2205);
    nand g39(n2112 ,n1906 ,n2004);
    not g40(n338 ,n2388);
    nor g41(n500 ,n8[22] ,n2[86]);
    or g42(n1475 ,n807 ,n1055);
    nor g43(n591 ,n296 ,n1);
    or g44(n875 ,n801 ,n806);
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n556), .Q(n7[6]));
    nor g46(n372 ,n8[5] ,n2360);
    nand g47(n1084 ,n640 ,n818);
    nand g48(n1151 ,n710 ,n892);
    not g49(n1307 ,n1179);
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n535), .Q(n7[8]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n543), .Q(n7[13]));
    nor g52(n1912 ,n1437 ,n1273);
    nor g53(n1530 ,n5[9] ,n1012);
    nor g54(n510 ,n8[24] ,n2[88]);
    not g55(n1677 ,n1592);
    nor g56(n973 ,n507 ,n269);
    nand g57(n616 ,n8[2] ,n2325);
    nand g58(n2023 ,n4[41] ,n1452);
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n585), .Q(n7[7]));
    or g60(n1474 ,n810 ,n1057);
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2166), .Q(n5[21]));
    nand g62(n2222 ,n3[36] ,n1887);
    nor g63(n213 ,n62 ,n212);
    nand g64(n627 ,n8[23] ,n2378);
    nor g65(n446 ,n8[22] ,n2[118]);
    nor g66(n167 ,n18 ,n166);
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2305), .Q(n3[47]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2172), .Q(n5[15]));
    not g69(n1216 ,n1088);
    nor g70(n929 ,n420 ,n805);
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n600), .Q(n7[14]));
    not g72(n1293 ,n1165);
    nor g73(n388 ,n8[7] ,n2362);
    nor g74(n1913 ,n1436 ,n1271);
    nor g75(n194 ,n75 ,n193);
    nand g76(n717 ,n8[20] ,n2[20]);
    not g77(n1305 ,n1177);
    or g78(n1480 ,n807 ,n1061);
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2104), .Q(n4[55]));
    nor g80(n199 ,n68 ,n198);
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2072), .Q(n4[23]));
    nor g82(n1408 ,n3[47] ,n1019);
    nor g83(n1955 ,n1508 ,n1306);
    or g84(n1632 ,n810 ,n1066);
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2301), .Q(n3[43]));
    xnor g86(n123 ,n2[52] ,n2[116]);
    not g87(n334 ,n2[0]);
    nand g88(n1097 ,n645 ,n836);
    nand g89(n2096 ,n1960 ,n1959);
    nor g90(n1439 ,n3[27] ,n1033);
    nor g91(n582 ,n329 ,n1);
    or g92(n1867 ,n1060 ,n1446);
    nor g93(n585 ,n303 ,n1);
    nand g94(n2141 ,n1763 ,n1762);
    nor g95(n443 ,n8[14] ,n2[78]);
    nor g96(n2043 ,n1550 ,n1707);
    not g97(n1257 ,n1129);
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2162), .Q(n4[45]));
    nand g99(n658 ,n2[33] ,n10[1]);
    nor g100(n963 ,n528 ,n875);
    nor g101(n258 ,n113 ,n257);
    nor g102(n896 ,n456 ,n804);
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2187), .Q(n5[57]));
    nor g104(n1966 ,n1516 ,n1209);
    not g105(n1664 ,n1579);
    nor g106(n555 ,n301 ,n1);
    nor g107(n904 ,n469 ,n804);
    nand g108(n1793 ,n4[6] ,n1469);
    nand g109(n659 ,n8[7] ,n2[7]);
    not g110(n1325 ,n1197);
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2169), .Q(n5[18]));
    not g112(n1702 ,n1617);
    nor g113(n1384 ,n5[0] ,n1037);
    nand g114(n676 ,n8[30] ,n2[126]);
    nand g115(n2017 ,n5[58] ,n1483);
    nand g116(n1186 ,n747 ,n925);
    xnor g117(n2375 ,n123 ,n239);
    not g118(n1321 ,n1193);
    nand g119(n2148 ,n1791 ,n1794);
    nor g120(n578 ,n284 ,n1);
    nor g121(n507 ,n8[26] ,n2[122]);
    nand g122(n732 ,n8[13] ,n2[13]);
    nor g123(n2401 ,n7[1] ,n7[0]);
    xnor g124(n103 ,n2[16] ,n2[80]);
    nor g125(n1410 ,n3[45] ,n1017);
    nor g126(n1940 ,n1495 ,n1294);
    nor g127(n1979 ,n1522 ,n1312);
    nor g128(n544 ,n326 ,n1);
    nor g129(n355 ,n8[7] ,n2[71]);
    nand g130(n793 ,n8[30] ,n2385);
    xnor g131(n2327 ,n101 ,n143);
    nor g132(n974 ,n493 ,n875);
    not g133(n1210 ,n1082);
    nor g134(n1975 ,n1520 ,n1685);
    nand g135(n2250 ,n3[8] ,n1883);
    nor g136(n1937 ,n1511 ,n1291);
    nand g137(n649 ,n8[24] ,n2[56]);
    nand g138(n1134 ,n705 ,n932);
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2194), .Q(n5[7]));
    nand g140(n2076 ,n1749 ,n1748);
    xnor g141(n132 ,n2[21] ,n2[85]);
    nor g142(n345 ,n8[31] ,n2[63]);
    nor g143(n1054 ,n8[19] ,n876);
    not g144(n1223 ,n1095);
    nor g145(n214 ,n120 ,n213);
    not g146(n1284 ,n1156);
    nor g147(n1759 ,n1345 ,n1311);
    not g148(n1319 ,n1191);
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2093), .Q(n4[2]));
    or g150(n2416 ,n2413 ,n2402);
    nor g151(n1364 ,n5[38] ,n1011);
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2076), .Q(n4[19]));
    nand g153(n2228 ,n3[30] ,n1861);
    nand g154(n2421 ,n2399 ,n2406);
    xnor g155(n125 ,n2[8] ,n2[72]);
    not g156(n2398 ,n7[25]);
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n559), .Q(n7[21]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2165), .Q(n5[22]));
    nand g159(n1800 ,n4[4] ,n1474);
    nand g160(n1824 ,n5[33] ,n1466);
    nor g161(n436 ,n8[21] ,n2344);
    not g162(n267 ,n266);
    xnor g163(n128 ,n2[53] ,n2[117]);
    xnor g164(n2338 ,n121 ,n165);
    nand g165(n2056 ,n4[31] ,n1482);
    nand g166(n1612 ,n669 ,n960);
    nand g167(n2151 ,n1809 ,n1807);
    nand g168(n1746 ,n5[46] ,n1648);
    nand g169(n2145 ,n1804 ,n1795);
    nand g170(n2010 ,n4[45] ,n1485);
    nand g171(n645 ,n8[26] ,n2[58]);
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n549), .Q(n7[25]));
    nor g173(n188 ,n82 ,n187);
    nand g174(n2211 ,n3[47] ,n1876);
    nor g175(n1359 ,n4[9] ,n1012);
    nand g176(n943 ,n9[1] ,n810);
    nor g177(n164 ,n119 ,n163);
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n541), .Q(n7[12]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2153), .Q(n5[34]));
    nand g180(n1961 ,n4[62] ,n1634);
    xnor g181(n2332 ,n110 ,n153);
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2310), .Q(n3[52]));
    nand g183(n688 ,n8[23] ,n2346);
    nor g184(n1980 ,n1524 ,n1687);
    xnor g185(n2356 ,n97 ,n201);
    nor g186(n186 ,n87 ,n185);
    nor g187(n407 ,n8[11] ,n2[75]);
    nand g188(n2109 ,n1997 ,n1996);
    nand g189(n1994 ,n4[51] ,n1468);
    not g190(n1315 ,n1187);
    nor g191(n1936 ,n1502 ,n1293);
    xnor g192(n2345 ,n134 ,n179);
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2167), .Q(n5[20]));
    nor g194(n1065 ,n8[28] ,n876);
    nand g195(n2270 ,n1928 ,n2238);
    nand g196(n2266 ,n1921 ,n2234);
    xnor g197(n2341 ,n127 ,n171);
    nor g198(n1921 ,n1387 ,n1278);
    nand g199(n1727 ,n4[25] ,n1454);
    xnor g200(n108 ,n2[36] ,n2[100]);
    nand g201(n718 ,n8[8] ,n2[104]);
    not g202(n1674 ,n1589);
    nand g203(n680 ,n8[7] ,n2[39]);
    nor g204(n886 ,n440 ,n804);
    nand g205(n2224 ,n3[34] ,n1889);
    nand g206(n1997 ,n4[50] ,n1647);
    nor g207(n924 ,n490 ,n804);
    nor g208(n939 ,n530 ,n805);
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n550), .Q(n8[13]));
    nand g210(n1039 ,n8[5] ,n877);
    nor g211(n2048 ,n1528 ,n1708);
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2188), .Q(n5[56]));
    nand g213(n2173 ,n1944 ,n1948);
    nand g214(n1030 ,n8[7] ,n877);
    nand g215(n2261 ,n1911 ,n2229);
    nand g216(n1848 ,n5[28] ,n1477);
    nor g217(n893 ,n451 ,n271);
    nand g218(n1801 ,n5[37] ,n1636);
    nand g219(n2316 ,n1829 ,n2200);
    nor g220(n975 ,n494 ,n875);
    nand g221(n1129 ,n683 ,n866);
    nor g222(n1412 ,n5[63] ,n1036);
    nor g223(n1760 ,n1349 ,n1663);
    nand g224(n781 ,n8[22] ,n2377);
    not g225(n330 ,n2[29]);
    nor g226(n1533 ,n4[49] ,n1021);
    nor g227(n1004 ,n510 ,n875);
    nand g228(n710 ,n8[19] ,n2342);
    xnor g229(n2343 ,n130 ,n175);
    nand g230(n2008 ,n4[46] ,n1479);
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2303), .Q(n3[45]));
    nor g232(n827 ,n345 ,n804);
    nand g233(n2012 ,n5[59] ,n1448);
    nor g234(n885 ,n471 ,n805);
    nor g235(n142 ,n99 ,n141);
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2297), .Q(n3[39]));
    xnor g237(n84 ,n2[44] ,n2[108]);
    nand g238(n761 ,n8[19] ,n2[83]);
    nor g239(n1528 ,n4[34] ,n1027);
    nor g240(n819 ,n388 ,n805);
    not g241(n317 ,n2[14]);
    nor g242(n1732 ,n1336 ,n1655);
    nor g243(n1942 ,n1491 ,n1295);
    not g244(n1660 ,n1575);
    nor g245(n144 ,n101 ,n143);
    xnor g246(n2336 ,n118 ,n161);
    nand g247(n643 ,n8[4] ,n2[4]);
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2156), .Q(n5[31]));
    nor g249(n148 ,n136 ,n147);
    not g250(n296 ,n2[43]);
    nand g251(n1133 ,n685 ,n869);
    nand g252(n1128 ,n693 ,n863);
    or g253(n1633 ,n807 ,n1054);
    nand g254(n2188 ,n2032 ,n2030);
    nand g255(n2247 ,n3[11] ,n1880);
    not g256(n1673 ,n1588);
    nand g257(n2137 ,n1740 ,n1726);
    nand g258(n1596 ,n763 ,n977);
    nor g259(n1007 ,n418 ,n875);
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n534), .Q(n8[7]));
    or g261(n1471 ,n807 ,n1067);
    xnor g262(n77 ,n2[28] ,n2[92]);
    nor g263(n2040 ,n1371 ,n1706);
    nor g264(n1417 ,n3[42] ,n1041);
    nor g265(n1051 ,n8[9] ,n876);
    dff g266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2127), .Q(n4[32]));
    dff g267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2291), .Q(n3[33]));
    nand g268(n1976 ,n4[57] ,n1454);
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n572), .Q(n7[5]));
    not g270(n1711 ,n1626);
    or g271(n1647 ,n810 ,n1053);
    not g272(n269 ,n268);
    nand g273(n2191 ,n2052 ,n2047);
    nand g274(n2225 ,n3[33] ,n1874);
    nand g275(n2226 ,n3[32] ,n1859);
    not g276(n1690 ,n1605);
    nor g277(n143 ,n67 ,n142);
    dff g278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2191), .Q(n5[53]));
    nor g279(n529 ,n8[18] ,n2373);
    not g280(n308 ,n2[1]);
    nand g281(n707 ,n8[25] ,n2[25]);
    nor g282(n832 ,n477 ,n804);
    not g283(n2395 ,n7[20]);
    nor g284(n453 ,n338 ,n1);
    not g285(n1275 ,n1147);
    nand g286(n1803 ,n4[3] ,n1478);
    nand g287(n1114 ,n661 ,n849);
    nand g288(n1575 ,n746 ,n999);
    nand g289(n1143 ,n623 ,n882);
    nor g290(n184 ,n86 ,n183);
    nand g291(n2078 ,n1754 ,n1753);
    or g292(n1642 ,n807 ,n1057);
    nor g293(n411 ,n8[27] ,n2350);
    nand g294(n696 ,n8[10] ,n2365);
    nand g295(n622 ,n8[5] ,n2[69]);
    nor g296(n1731 ,n1335 ,n1319);
    xnor g297(n2351 ,n77 ,n191);
    nand g298(n1953 ,n5[13] ,n1646);
    nor g299(n1405 ,n5[59] ,n1033);
    nand g300(n2240 ,n3[18] ,n1873);
    nand g301(n727 ,n8[15] ,n2[15]);
    nand g302(n2157 ,n1837 ,n1834);
    nand g303(n265 ,n6[2] ,n264);
    nand g304(n1136 ,n688 ,n870);
    nand g305(n633 ,n2[65] ,n10[1]);
    nand g306(n2085 ,n1779 ,n1778);
    nand g307(n775 ,n8[25] ,n2[89]);
    not g308(n1324 ,n1196);
    nor g309(n161 ,n31 ,n160);
    nor g310(n1807 ,n1368 ,n1215);
    nor g311(n380 ,n6[0] ,n1);
    not g312(n1203 ,n1075);
    nor g313(n2024 ,n1543 ,n1320);
    nand g314(n2006 ,n5[60] ,n1477);
    nor g315(n1995 ,n1529 ,n1226);
    not g316(n264 ,n263);
    nand g317(n747 ,n8[13] ,n2[45]);
    xnor g318(n2340 ,n124 ,n169);
    nand g319(n1752 ,n5[45] ,n1646);
    or g320(n1877 ,n1048 ,n1446);
    nor g321(n602 ,n278 ,n1);
    dff g322(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2287), .Q(n3[3]));
    nor g323(n1357 ,n4[10] ,n1041);
    nor g324(n1963 ,n1515 ,n1308);
    nor g325(n361 ,n8[2] ,n2[2]);
    not g326(n320 ,n2[54]);
    nor g327(n1827 ,n1386 ,n1224);
    nor g328(n942 ,n529 ,n805);
    nand g329(n1777 ,n5[2] ,n1489);
    nand g330(n1782 ,n5[40] ,n1639);
    nand g331(n2105 ,n1984 ,n1983);
    nor g332(n155 ,n42 ,n154);
    nor g333(n1951 ,n1498 ,n1302);
    not g334(n287 ,n2[20]);
    xnor g335(n117 ,n2[51] ,n2[115]);
    nor g336(n990 ,n505 ,n875);
    nor g337(n1523 ,n5[52] ,n1024);
    nor g338(n905 ,n395 ,n804);
    nand g339(n2257 ,n3[1] ,n1874);
    dff g340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2083), .Q(n4[12]));
    dff g341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2150), .Q(n5[0]));
    nor g342(n1504 ,n5[16] ,n1020);
    nor g343(n1345 ,n5[3] ,n1016);
    nor g344(n1433 ,n5[22] ,n1026);
    nand g345(n2407 ,n7[21] ,n2395);
    nor g346(n395 ,n8[13] ,n2[13]);
    nand g347(n2233 ,n3[25] ,n1866);
    xnor g348(n112 ,n2[10] ,n2[74]);
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2266), .Q(n3[24]));
    not g350(n271 ,n270);
    nand g351(n2058 ,n5[52] ,n1475);
    dff g352(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2320), .Q(n3[62]));
    nor g353(n438 ,n8[8] ,n2[8]);
    nand g354(n1791 ,n5[38] ,n1635);
    nand g355(n1122 ,n752 ,n857);
    nand g356(n2234 ,n3[24] ,n1867);
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2183), .Q(n5[8]));
    nor g358(n960 ,n518 ,n269);
    not g359(n1676 ,n1591);
    xnor g360(n116 ,n2[38] ,n2[102]);
    nand g361(n738 ,n8[29] ,n2384);
    xnor g362(n102 ,n2[34] ,n2[98]);
    nor g363(n367 ,n8[13] ,n2[77]);
    nand g364(n1152 ,n711 ,n891);
    nand g365(n1103 ,n750 ,n841);
    nor g366(n226 ,n78 ,n225);
    nor g367(n1828 ,n1390 ,n1228);
    nor g368(n1444 ,n4[48] ,n1020);
    nor g369(n2065 ,n1564 ,n1714);
    xnor g370(n109 ,n2[50] ,n2[114]);
    xnor g371(n133 ,n2[55] ,n2[119]);
    nand g372(n2150 ,n1784 ,n1853);
    nor g373(n517 ,n8[18] ,n2341);
    nor g374(n897 ,n462 ,n805);
    not g375(n1296 ,n1168);
    nor g376(n2429 ,n2423 ,n2428);
    or g377(n1634 ,n810 ,n1067);
    not g378(n1669 ,n1584);
    nor g379(n899 ,n457 ,n804);
    nand g380(n669 ,n8[13] ,n2[109]);
    nor g381(n1720 ,n1544 ,n1652);
    nand g382(n1811 ,n4[1] ,n1490);
    nor g383(n1383 ,n3[60] ,n1034);
    nor g384(n1964 ,n1354 ,n1681);
    not g385(n310 ,n2[40]);
    nor g386(n895 ,n567 ,n271);
    not g387(n1290 ,n1162);
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2102), .Q(n4[57]));
    not g389(n1277 ,n1149);
    dff g390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2271), .Q(n3[19]));
    dff g391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2103), .Q(n4[56]));
    nor g392(n1069 ,n10[0] ,n876);
    not g393(n1318 ,n1190);
    xnor g394(n124 ,n2[17] ,n2[81]);
    dff g395(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2311), .Q(n3[53]));
    nand g396(n1775 ,n4[11] ,n1487);
    nand g397(n684 ,n8[13] ,n2336);
    nor g398(n224 ,n84 ,n223);
    nor g399(n228 ,n76 ,n227);
    not g400(n1212 ,n1084);
    nand g401(n1992 ,n5[62] ,n1471);
    xnor g402(n2365 ,n131 ,n219);
    nand g403(n652 ,n8[30] ,n2353);
    nand g404(n1170 ,n739 ,n910);
    not g405(n1265 ,n1137);
    nor g406(n1440 ,n5[20] ,n1024);
    nand g407(n606 ,n8[26] ,n2[122]);
    nand g408(n1154 ,n715 ,n895);
    nor g409(n160 ,n115 ,n159);
    nor g410(n231 ,n11 ,n230);
    nor g411(n1424 ,n5[24] ,n1029);
    nand g412(n2298 ,n1891 ,n2218);
    nand g413(n1023 ,n8[19] ,n877);
    not g414(n278 ,n2[35]);
    xnor g415(n2382 ,n100 ,n253);
    nand g416(n704 ,n8[26] ,n2[26]);
    nand g417(n2312 ,n1835 ,n2204);
    nor g418(n997 ,n465 ,n875);
    nand g419(n638 ,n8[7] ,n2362);
    nand g420(n1852 ,n5[27] ,n1448);
    nor g421(n818 ,n369 ,n805);
    not g422(n1313 ,n1185);
    not g423(n1240 ,n1112);
    or g424(n1469 ,n810 ,n1043);
    dff g425(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n584), .Q(n7[23]));
    not g426(n1269 ,n1141);
    nor g427(n1716 ,n1332 ,n1651);
    nor g428(n162 ,n118 ,n161);
    xnor g429(n2333 ,n112 ,n155);
    not g430(n316 ,n2[32]);
    not g431(n298 ,n2[60]);
    xnor g432(n2370 ,n81 ,n229);
    nor g433(n241 ,n44 ,n240);
    nor g434(n890 ,n343 ,n271);
    nand g435(n1118 ,n668 ,n853);
    nor g436(n429 ,n2[32] ,n10[0]);
    nor g437(n1952 ,n1505 ,n1304);
    nor g438(n845 ,n354 ,n804);
    dff g439(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2139), .Q(n5[3]));
    dff g440(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n579), .Q(n8[28]));
    nor g441(n545 ,n293 ,n1);
    nor g442(n475 ,n8[17] ,n2[81]);
    nand g443(n1786 ,n4[8] ,n1453);
    or g444(n1890 ,n1052 ,n1446);
    nand g445(n141 ,n72 ,n140);
    nor g446(n1377 ,n3[63] ,n1036);
    dff g447(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2138), .Q(n5[45]));
    nand g448(n2206 ,n3[52] ,n1871);
    dff g449(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2270), .Q(n3[20]));
    not g450(n326 ,n2[11]);
    not g451(n1683 ,n1598);
    nor g452(n1891 ,n1420 ,n1253);
    nor g453(n1795 ,n1361 ,n1212);
    nor g454(n526 ,n8[25] ,n2[57]);
    nor g455(n536 ,n324 ,n1);
    nand g456(n666 ,n8[27] ,n2350);
    nor g457(n1520 ,n4[57] ,n1031);
    nor g458(n1553 ,n5[53] ,n1025);
    nor g459(n171 ,n41 ,n170);
    or g460(n1860 ,n1044 ,n1446);
    nor g461(n190 ,n79 ,n189);
    or g462(n1482 ,n810 ,n1044);
    nand g463(n1100 ,n647 ,n837);
    nand g464(n794 ,n8[25] ,n2380);
    nand g465(n1201 ,n637 ,n828);
    nand g466(n2310 ,n1838 ,n2206);
    nor g467(n1503 ,n4[18] ,n1022);
    dff g468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2272), .Q(n3[18]));
    nand g469(n2274 ,n1904 ,n2226);
    nand g470(n2118 ,n2023 ,n2022);
    nand g471(n1041 ,n8[10] ,n877);
    nor g472(n466 ,n8[16] ,n2[16]);
    nand g473(n2139 ,n1742 ,n1759);
    nand g474(n754 ,n8[4] ,n2[36]);
    nor g475(n256 ,n94 ,n255);
    nand g476(n2143 ,n1858 ,n1769);
    nor g477(n1914 ,n1439 ,n1274);
    not g478(n329 ,n2[19]);
    not g479(n1703 ,n1618);
    dff g480(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2268), .Q(n3[22]));
    dff g481(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2322), .Q(n3[16]));
    nor g482(n452 ,n8[8] ,n2[104]);
    or g483(n1461 ,n807 ,n1060);
    nand g484(n730 ,n8[14] ,n2[14]);
    nor g485(n2004 ,n1537 ,n1695);
    dff g486(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2088), .Q(n4[7]));
    nor g487(n1539 ,n5[8] ,n1010);
    not g488(n1244 ,n1116);
    nor g489(n1989 ,n1530 ,n1240);
    nand g490(n1808 ,n4[2] ,n1486);
    nor g491(n62 ,n2[38] ,n2[102]);
    dff g492(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2306), .Q(n3[48]));
    nand g493(n646 ,n8[31] ,n2386);
    nor g494(n998 ,n475 ,n875);
    nor g495(n27 ,n2[42] ,n2[106]);
    nor g496(n1446 ,n1 ,n1008);
    nor g497(n2009 ,n1401 ,n1697);
    nor g498(n202 ,n97 ,n201);
    not g499(n1252 ,n1124);
    nor g500(n1495 ,n3[13] ,n1017);
    dff g501(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2164), .Q(n5[23]));
    nand g502(n1603 ,n692 ,n969);
    nand g503(n2116 ,n2029 ,n2016);
    nor g504(n2417 ,n2409 ,n2407);
    not g505(n1697 ,n1612);
    dff g506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2145), .Q(n5[1]));
    nand g507(n1168 ,n769 ,n856);
    not g508(n1705 ,n1620);
    nor g509(n382 ,n8[17] ,n2[113]);
    or g510(n1481 ,n810 ,n1049);
    dff g511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n542), .Q(n8[30]));
    nand g512(n2294 ,n1897 ,n2222);
    nand g513(n2185 ,n2037 ,n2046);
    nand g514(n628 ,n8[3] ,n2[67]);
    not g515(n1242 ,n1114);
    dff g516(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2141), .Q(n5[43]));
    nor g517(n2036 ,n1344 ,n1324);
    nand g518(n660 ,n8[25] ,n2[121]);
    nand g519(n767 ,n8[8] ,n2331);
    nand g520(n795 ,n8[18] ,n2373);
    not g521(n266 ,n805);
    nor g522(n240 ,n123 ,n239);
    nor g523(n575 ,n292 ,n1);
    nand g524(n745 ,n8[6] ,n2361);
    nand g525(n1099 ,n783 ,n838);
    xnor g526(n2378 ,n133 ,n245);
    dff g527(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2294), .Q(n3[36]));
    not g528(n1678 ,n1593);
    nor g529(n1839 ,n1402 ,n1236);
    not g530(n1224 ,n1096);
    nor g531(n1388 ,n4[44] ,n1015);
    nor g532(n1841 ,n1403 ,n1239);
    nand g533(n632 ,n8[2] ,n2[66]);
    nor g534(n342 ,n8[30] ,n2[62]);
    nor g535(n435 ,n8[25] ,n2348);
    nand g536(n728 ,n8[3] ,n2[3]);
    xnor g537(n2379 ,n93 ,n247);
    nor g538(n825 ,n521 ,n805);
    nand g539(n2075 ,n1744 ,n1743);
    nor g540(n253 ,n52 ,n252);
    nor g541(n1535 ,n4[42] ,n1041);
    nand g542(n1584 ,n653 ,n990);
    nor g543(n247 ,n13 ,n246);
    not g544(n1666 ,n1581);
    nand g545(n2069 ,n1721 ,n1720);
    nor g546(n239 ,n36 ,n238);
    nand g547(n2140 ,n1756 ,n1755);
    not g548(n1231 ,n1103);
    xnor g549(n118 ,n2[13] ,n2[77]);
    nand g550(n2183 ,n2021 ,n2015);
    not g551(n273 ,n1);
    nor g552(n843 ,n532 ,n271);
    nand g553(n2114 ,n1895 ,n1893);
    or g554(n1473 ,n810 ,n1052);
    nor g555(n1404 ,n3[49] ,n1021);
    or g556(n1885 ,n1043 ,n1446);
    nor g557(n1402 ,n3[51] ,n1023);
    nor g558(n587 ,n330 ,n1);
    or g559(n1464 ,n810 ,n1055);
    dff g560(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2111), .Q(n4[48]));
    nor g561(n1058 ,n8[22] ,n876);
    nor g562(n1349 ,n4[15] ,n1019);
    dff g563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2147), .Q(n5[39]));
    nor g564(n473 ,n8[23] ,n2[55]);
    nor g565(n1003 ,n503 ,n875);
    nor g566(n1833 ,n1392 ,n1230);
    nor g567(n1898 ,n1424 ,n1257);
    dff g568(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2277), .Q(n3[14]));
    nor g569(n1063 ,n8[8] ,n876);
    nor g570(n481 ,n8[10] ,n2[10]);
    not g571(n1289 ,n1161);
    nor g572(n909 ,n360 ,n267);
    nand g573(n2186 ,n2017 ,n2018);
    nand g574(n1189 ,n767 ,n878);
    nor g575(n2050 ,n1552 ,n1709);
    nand g576(n1144 ,n695 ,n883);
    nor g577(n2007 ,n1538 ,n1696);
    nor g578(n19 ,n2[33] ,n2[97]);
    nor g579(n176 ,n130 ,n175);
    dff g580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n539), .Q(n8[26]));
    dff g581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2319), .Q(n3[61]));
    nand g582(n1965 ,n4[61] ,n1632);
    nor g583(n2389 ,n264 ,n262);
    nand g584(n2295 ,n1896 ,n2221);
    dff g585(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2070), .Q(n4[25]));
    nand g586(n2268 ,n1924 ,n2236);
    nor g587(n1717 ,n1331 ,n1202);
    not g588(n319 ,n2[53]);
    nand g589(n2260 ,n1909 ,n2228);
    not g590(n1278 ,n1150);
    dff g591(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2276), .Q(n3[13]));
    nor g592(n222 ,n135 ,n221);
    nor g593(n1423 ,n3[37] ,n1039);
    nor g594(n146 ,n104 ,n145);
    dff g595(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2173), .Q(n5[14]));
    xnor g596(n129 ,n2[19] ,n2[83]);
    nand g597(n2000 ,n4[49] ,n1473);
    nand g598(n1991 ,n4[52] ,n1464);
    nor g599(n527 ,n8[17] ,n2[49]);
    nor g600(n984 ,n368 ,n269);
    xnor g601(n98 ,n2[49] ,n2[113]);
    nor g602(n31 ,n2[12] ,n2[76]);
    nor g603(n959 ,n397 ,n269);
    not g604(n337 ,n2[17]);
    nand g605(n808 ,n9[1] ,n802);
    nor g606(n12 ,n2[29] ,n2[93]);
    dff g607(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2091), .Q(n4[4]));
    xnor g608(n2380 ,n105 ,n249);
    nor g609(n1420 ,n3[40] ,n1010);
    not g610(n1227 ,n1099);
    nand g611(n2246 ,n3[12] ,n1879);
    dff g612(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2117), .Q(n4[42]));
    nor g613(n1360 ,n5[39] ,n1030);
    nor g614(n2028 ,n1546 ,n1703);
    or g615(n1863 ,n1065 ,n1446);
    nand g616(n1094 ,n743 ,n832);
    nor g617(n49 ,n2[28] ,n2[92]);
    nor g618(n813 ,n511 ,n805);
    not g619(n1248 ,n1120);
    nand g620(n624 ,n2[1] ,n10[1]);
    dff g621(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2100), .Q(n4[59]));
    xnor g622(n2377 ,n85 ,n243);
    nand g623(n1121 ,n673 ,n867);
    xnor g624(n2354 ,n83 ,n197);
    dff g625(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2099), .Q(n4[60]));
    nand g626(n750 ,n8[22] ,n2[54]);
    not g627(n1661 ,n1576);
    nor g628(n52 ,n2[58] ,n2[122]);
    xnor g629(n2350 ,n79 ,n189);
    nor g630(n580 ,n340 ,n1);
    nand g631(n2125 ,n2049 ,n2048);
    nor g632(n966 ,n516 ,n269);
    nand g633(n2263 ,n1914 ,n2231);
    dff g634(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2130), .Q(n4[29]));
    nand g635(n2092 ,n1803 ,n1802);
    nor g636(n1547 ,n5[7] ,n1030);
    nand g637(n779 ,n8[27] ,n2[91]);
    nand g638(n1123 ,n672 ,n854);
    nor g639(n547 ,n310 ,n1);
    nand g640(n711 ,n8[23] ,n2[23]);
    nor g641(n516 ,n8[19] ,n2[115]);
    or g642(n1644 ,n807 ,n1046);
    nor g643(n465 ,n8[16] ,n2[80]);
    nand g644(n139 ,n15 ,n138);
    nand g645(n2111 ,n2002 ,n1920);
    nor g646(n503 ,n8[23] ,n2[87]);
    nor g647(n254 ,n100 ,n253);
    nand g648(n2099 ,n1968 ,n1967);
    nand g649(n712 ,n8[15] ,n2[79]);
    nor g650(n44 ,n2[52] ,n2[116]);
    nand g651(n1619 ,n611 ,n953);
    nand g652(n2002 ,n4[48] ,n1476);
    dff g653(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2154), .Q(n5[33]));
    nor g654(n1414 ,n4[11] ,n1014);
    nor g655(n1856 ,n1416 ,n1251);
    not g656(n1327 ,n1199);
    xnor g657(n137 ,n2[23] ,n2[87]);
    not g658(n876 ,n877);
    dff g659(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2285), .Q(n3[5]));
    nand g660(n789 ,n8[18] ,n2[50]);
    nand g661(n2202 ,n3[56] ,n1867);
    nor g662(n28 ,n2[50] ,n2[114]);
    dff g663(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2315), .Q(n3[57]));
    nor g664(n1500 ,n3[14] ,n1018);
    nor g665(n872 ,n426 ,n271);
    nand g666(n1620 ,n614 ,n952);
    nand g667(n2165 ,n1910 ,n1908);
    nor g668(n961 ,n482 ,n269);
    nor g669(n1817 ,n1377 ,n1204);
    nand g670(n1106 ,n631 ,n843);
    nor g671(n373 ,n8[11] ,n2[107]);
    nand g672(n2181 ,n2003 ,n1989);
    nor g673(n349 ,n8[29] ,n2[61]);
    dff g674(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n453), .Q(n6[2]));
    nor g675(n815 ,n455 ,n805);
    nor g676(n201 ,n43 ,n200);
    nor g677(n1799 ,n1366 ,n1674);
    nor g678(n36 ,n2[51] ,n2[115]);
    nand g679(n785 ,n8[20] ,n2375);
    nor g680(n1560 ,n5[51] ,n1023);
    xnor g681(n85 ,n2[54] ,n2[118]);
    nand g682(n629 ,n8[29] ,n2[93]);
    nor g683(n244 ,n85 ,n243);
    nor g684(n428 ,n8[2] ,n2[34]);
    not g685(n1311 ,n1183);
    nand g686(n2217 ,n3[41] ,n1882);
    or g687(n1650 ,n810 ,n1065);
    dff g688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2181), .Q(n5[9]));
    not g689(n294 ,n2[47]);
    nand g690(n2171 ,n1941 ,n1939);
    nor g691(n1561 ,n4[29] ,n1035);
    xnor g692(n2330 ,n107 ,n149);
    nand g693(n2208 ,n3[50] ,n1873);
    nand g694(n2315 ,n1830 ,n2201);
    dff g695(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2281), .Q(n3[9]));
    dff g696(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n912), .Q(n9[0]));
    nor g697(n1938 ,n1500 ,n1292);
    nand g698(n1580 ,n691 ,n994);
    nand g699(n2287 ,n1958 ,n2255);
    not g700(n1295 ,n1167);
    nor g701(n29 ,n2[10] ,n2[74]);
    xor g702(n2325 ,n96 ,n139);
    nand g703(n1723 ,n5[5] ,n1636);
    nand g704(n1111 ,n789 ,n846);
    nand g705(n2014 ,n4[44] ,n1484);
    nor g706(n1830 ,n1389 ,n1227);
    or g707(n2423 ,n2418 ,n2420);
    nand g708(n2232 ,n3[26] ,n1865);
    nand g709(n1783 ,n4[9] ,n1452);
    dff g710(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2288), .Q(n3[2]));
    nor g711(n1009 ,n409 ,n875);
    nor g712(n1385 ,n3[59] ,n1033);
    dff g713(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2278), .Q(n3[12]));
    nor g714(n837 ,n399 ,n805);
    nor g715(n2066 ,n1521 ,n1686);
    nor g716(n1066 ,n8[29] ,n876);
    or g717(n1639 ,n807 ,n1063);
    nor g718(n223 ,n59 ,n222);
    dff g719(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n544), .Q(n7[11]));
    nand g720(n1601 ,n741 ,n971);
    nor g721(n25 ,n2[8] ,n2[72]);
    nand g722(n1627 ,n749 ,n946);
    dff g723(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2312), .Q(n3[54]));
    nor g724(n2053 ,n1556 ,n1710);
    nand g725(n759 ,n8[4] ,n2[100]);
    dff g726(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2193), .Q(n5[51]));
    nand g727(n2308 ,n1841 ,n2208);
    or g728(n1483 ,n807 ,n1062);
    dff g729(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n944), .Q(n9[1]));
    nor g730(n1838 ,n1399 ,n1235);
    nand g731(n1165 ,n733 ,n906);
    nand g732(n2079 ,n1758 ,n1757);
    nor g733(n951 ,n514 ,n875);
    not g734(n1279 ,n1151);
    nor g735(n420 ,n8[9] ,n2332);
    xnor g736(n2374 ,n117 ,n237);
    nor g737(n1818 ,n1378 ,n1329);
    nor g738(n470 ,n8[19] ,n2[19]);
    nand g739(n1587 ,n617 ,n987);
    nand g740(n2134 ,n1730 ,n1731);
    dff g741(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n599), .Q(n8[1]));
    nor g742(n903 ,n467 ,n267);
    not g743(n1684 ,n1599);
    nor g744(n449 ,n8[6] ,n2[6]);
    nor g745(n852 ,n411 ,n805);
    nand g746(n1779 ,n4[10] ,n1447);
    nand g747(n790 ,n8[5] ,n2328);
    nor g748(n1509 ,n4[50] ,n1022);
    nor g749(n2405 ,n2391 ,n7[18]);
    nand g750(n673 ,n8[9] ,n2364);
    nand g751(n2269 ,n1927 ,n2237);
    nor g752(n1342 ,n4[19] ,n1023);
    nor g753(n531 ,n8[29] ,n2[125]);
    nand g754(n1582 ,n670 ,n992);
    dff g755(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n571), .Q(n8[25]));
    nand g756(n724 ,n8[16] ,n2[16]);
    or g757(n1868 ,n1059 ,n1446);
    nor g758(n579 ,n298 ,n1);
    not g759(n332 ,n2[26]);
    nor g760(n833 ,n390 ,n805);
    nor g761(n1421 ,n3[39] ,n1030);
    nand g762(n1096 ,n731 ,n833);
    nand g763(n1119 ,n651 ,n921);
    nand g764(n1107 ,n620 ,n816);
    nor g765(n67 ,n2[3] ,n2[67]);
    nand g766(n1191 ,n770 ,n811);
    dff g767(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n588), .Q(n7[15]));
    nor g768(n1993 ,n1396 ,n1691);
    dff g769(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2298), .Q(n3[40]));
    nor g770(n945 ,n379 ,n269);
    nor g771(n480 ,n8[18] ,n2[50]);
    nand g772(n2182 ,n2006 ,n2005);
    nor g773(n154 ,n110 ,n153);
    not g774(n1214 ,n1086);
    nand g775(n2179 ,n1992 ,n1995);
    nor g776(n987 ,n408 ,n875);
    nor g777(n1847 ,n1409 ,n1246);
    xnor g778(n79 ,n2[27] ,n2[91]);
    nand g779(n1083 ,n657 ,n848);
    nand g780(n2169 ,n1930 ,n1926);
    nor g781(n1739 ,n1527 ,n1657);
    not g782(n1317 ,n1189);
    nor g783(n999 ,n444 ,n875);
    dff g784(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2282), .Q(n3[8]));
    xnor g785(n2339 ,n103 ,n167);
    or g786(n1645 ,n807 ,n1072);
    xnor g787(n81 ,n2[47] ,n2[111]);
    nand g788(n675 ,n8[9] ,n2[41]);
    nor g789(n2018 ,n1541 ,n1238);
    nand g790(n1120 ,n671 ,n855);
    nand g791(n1842 ,n5[29] ,n1488);
    nor g792(n1416 ,n5[26] ,n1032);
    nand g793(n1742 ,n5[3] ,n1645);
    nand g794(n1604 ,n703 ,n968);
    nand g795(n2167 ,n1919 ,n1917);
    nor g796(n457 ,n8[18] ,n2[18]);
    nor g797(n1928 ,n1549 ,n1284);
    nand g798(n1092 ,n655 ,n831);
    nor g799(n353 ,n8[6] ,n2[102]);
    nor g800(n432 ,n8[31] ,n2[31]);
    xnor g801(n2328 ,n104 ,n145);
    xnor g802(n115 ,n2[12] ,n2[76]);
    nor g803(n468 ,n8[15] ,n2[15]);
    nand g804(n623 ,n8[21] ,n2344);
    nor g805(n403 ,n8[8] ,n2363);
    dff g806(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n563), .Q(n8[23]));
    nor g807(n412 ,n8[11] ,n2[43]);
    not g808(n1304 ,n1176);
    nor g809(n574 ,n302 ,n1);
    nor g810(n992 ,n407 ,n875);
    dff g811(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2179), .Q(n5[62]));
    nor g812(n1929 ,n1548 ,n1285);
    dff g813(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2185), .Q(n5[6]));
    nor g814(n166 ,n121 ,n165);
    nand g815(n1586 ,n634 ,n988);
    nor g816(n912 ,n799 ,n809);
    nor g817(n504 ,n8[5] ,n2328);
    nor g818(n864 ,n423 ,n805);
    xor g819(n2324 ,n91 ,n73);
    nor g820(n396 ,n8[8] ,n2[72]);
    nand g821(n1751 ,n4[18] ,n1647);
    nor g822(n69 ,n2[30] ,n2[94]);
    nand g823(n692 ,n8[22] ,n2[118]);
    nand g824(n2064 ,n5[51] ,n1633);
    not g825(n1322 ,n1194);
    nand g826(n1105 ,n729 ,n935);
    not g827(n270 ,n804);
    nor g828(n447 ,n8[25] ,n2[25]);
    nand g829(n1017 ,n8[13] ,n877);
    dff g830(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2098), .Q(n4[61]));
    nand g831(n2301 ,n1854 ,n2215);
    nand g832(n1804 ,n5[1] ,n1466);
    nand g833(n1628 ,n629 ,n945);
    nor g834(n562 ,n322 ,n1);
    nor g835(n68 ,n2[31] ,n2[95]);
    nor g836(n828 ,n346 ,n805);
    not g837(n1685 ,n1600);
    nor g838(n581 ,n313 ,n1);
    xnor g839(n2346 ,n137 ,n181);
    nand g840(n2214 ,n3[44] ,n1879);
    xnor g841(n94 ,n2[60] ,n2[124]);
    nand g842(n1968 ,n4[60] ,n1650);
    nand g843(n2302 ,n1851 ,n2214);
    nor g844(n871 ,n428 ,n804);
    nor g845(n1429 ,n3[33] ,n1038);
    nor g846(n1908 ,n1433 ,n1269);
    dff g847(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2080), .Q(n4[15]));
    nor g848(n490 ,n8[3] ,n2[3]);
    not g849(n1306 ,n1178);
    nor g850(n389 ,n8[24] ,n2347);
    xnor g851(n80 ,n2[30] ,n2[94]);
    nor g852(n829 ,n342 ,n804);
    or g853(n1649 ,n807 ,n1050);
    nand g854(n699 ,n8[28] ,n2[28]);
    not g855(n312 ,n2[15]);
    not g856(n1663 ,n1578);
    nor g857(n1849 ,n1410 ,n1314);
    nor g858(n1445 ,n3[58] ,n1032);
    not g859(n1253 ,n1125);
    nor g860(n442 ,n8[13] ,n2336);
    nor g861(n595 ,n323 ,n1);
    nor g862(n1365 ,n4[5] ,n1039);
    nand g863(n2297 ,n1892 ,n2219);
    nor g864(n243 ,n58 ,n242);
    nor g865(n1999 ,n1533 ,n1693);
    nor g866(n495 ,n8[21] ,n2[85]);
    nor g867(n1825 ,n1385 ,n1223);
    nand g868(n1600 ,n660 ,n972);
    nor g869(n1006 ,n520 ,n875);
    nor g870(n375 ,n8[30] ,n2353);
    nand g871(n755 ,n8[10] ,n2333);
    nor g872(n1510 ,n3[4] ,n1040);
    not g873(n1680 ,n1595);
    dff g874(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n557), .Q(n7[2]));
    nand g875(n757 ,n8[31] ,n2[31]);
    nor g876(n1726 ,n1338 ,n1318);
    nor g877(n1070 ,n8[2] ,n876);
    nor g878(n811 ,n512 ,n805);
    nand g879(n2122 ,n1734 ,n2035);
    nor g880(n552 ,n280 ,n1);
    nor g881(n1000 ,n489 ,n875);
    nand g882(n1011 ,n8[6] ,n877);
    nor g883(n1527 ,n4[21] ,n1025);
    nand g884(n1098 ,n793 ,n930);
    nor g885(n1334 ,n4[25] ,n1031);
    nor g886(n1555 ,n5[18] ,n1022);
    nor g887(n1850 ,n1411 ,n1245);
    not g888(n1651 ,n1566);
    nand g889(n2235 ,n3[23] ,n1868);
    nand g890(n1772 ,n4[12] ,n1484);
    nand g891(n2313 ,n1833 ,n2203);
    or g892(n1631 ,n807 ,n1049);
    nor g893(n177 ,n51 ,n176);
    nor g894(n1393 ,n3[54] ,n1026);
    dff g895(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2119), .Q(n4[40]));
    nand g896(n1194 ,n781 ,n941);
    nor g897(n485 ,n8[6] ,n2361);
    xnor g898(n121 ,n2[15] ,n2[79]);
    nand g899(n1174 ,n684 ,n914);
    nor g900(n1778 ,n1357 ,n1668);
    not g901(n1256 ,n1128);
    not g902(n1286 ,n1158);
    dff g903(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2097), .Q(n4[62]));
    nor g904(n921 ,n445 ,n804);
    nand g905(n2256 ,n3[2] ,n1889);
    nand g906(n2119 ,n2027 ,n2026);
    nor g907(n518 ,n8[13] ,n2[109]);
    nor g908(n906 ,n472 ,n805);
    nand g909(n2060 ,n4[30] ,n1634);
    nor g910(n197 ,n69 ,n196);
    not g911(n1679 ,n1594);
    nand g912(n2071 ,n1729 ,n1728);
    nor g913(n30 ,n2[37] ,n2[101]);
    nor g914(n1053 ,n8[18] ,n876);
    nand g915(n1715 ,n5[50] ,n1638);
    or g916(n1635 ,n807 ,n1043);
    nand g917(n784 ,n8[10] ,n2[74]);
    nor g918(n1052 ,n8[17] ,n876);
    nor g919(n848 ,n403 ,n805);
    nor g920(n570 ,n321 ,n1);
    nand g921(n2309 ,n1839 ,n2207);
    nor g922(n1920 ,n1444 ,n1694);
    nand g923(n2279 ,n1945 ,n2247);
    not g924(n1701 ,n1616);
    nand g925(n1074 ,n795 ,n942);
    nand g926(n2414 ,n7[7] ,n2396);
    nand g927(n1756 ,n5[44] ,n1644);
    not g928(n1239 ,n1111);
    not g929(n276 ,n2[37]);
    nand g930(n694 ,n8[30] ,n2[30]);
    nor g931(n178 ,n132 ,n177);
    nand g932(n2133 ,n1723 ,n1719);
    not g933(n311 ,n2[58]);
    nor g934(n920 ,n513 ,n804);
    not g935(n282 ,n2[21]);
    nor g936(n1840 ,n1398 ,n1237);
    nand g937(n715 ,n8[21] ,n2[21]);
    nand g938(n1182 ,n790 ,n940);
    nor g939(n413 ,n8[8] ,n2[40]);
    nor g940(n471 ,n8[2] ,n2325);
    xnor g941(n119 ,n2[14] ,n2[78]);
    nor g942(n242 ,n128 ,n241);
    nor g943(n1990 ,n1400 ,n1690);
    nand g944(n1721 ,n4[26] ,n1451);
    nor g945(n882 ,n436 ,n805);
    nand g946(n2095 ,n1816 ,n1814);
    nor g947(n55 ,n2[7] ,n2[71]);
    nand g948(n664 ,n8[15] ,n2[47]);
    nand g949(n687 ,n8[2] ,n2[34]);
    nand g950(n2128 ,n2056 ,n2055);
    nand g951(n2288 ,n1962 ,n2256);
    nand g952(n2044 ,n4[35] ,n1478);
    nand g953(n2098 ,n1965 ,n1964);
    nor g954(n250 ,n105 ,n249);
    not g955(n2392 ,n7[22]);
    nor g956(n2424 ,n2422 ,n2419);
    nor g957(n1409 ,n3[46] ,n1018);
    xnor g958(n2342 ,n129 ,n173);
    nand g959(n1172 ,n740 ,n911);
    nor g960(n417 ,n8[3] ,n2[35]);
    or g961(n1638 ,n807 ,n1053);
    nand g962(n2249 ,n3[9] ,n1882);
    not g963(n1211 ,n1083);
    nand g964(n2126 ,n2051 ,n2050);
    nand g965(n1025 ,n8[21] ,n877);
    nor g966(n206 ,n89 ,n205);
    nand g967(n1981 ,n4[55] ,n1458);
    nor g968(n1750 ,n1503 ,n1660);
    nor g969(n1524 ,n4[55] ,n1028);
    dff g970(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n575), .Q(n7[4]));
    nand g971(n1590 ,n628 ,n984);
    nor g972(n502 ,n8[9] ,n2[9]);
    nor g973(n351 ,n8[3] ,n2358);
    nor g974(n1045 ,n8[10] ,n876);
    nand g975(n2300 ,n1855 ,n2216);
    nand g976(n1905 ,n5[23] ,n1463);
    nand g977(n760 ,n8[22] ,n2[86]);
    not g978(n1329 ,n1201);
    nor g979(n401 ,n8[28] ,n2351);
    nand g980(n2291 ,n1903 ,n2225);
    nor g981(n534 ,n325 ,n1);
    nor g982(n235 ,n24 ,n234);
    nand g983(n1113 ,n792 ,n847);
    or g984(n10[0] ,n8[0] ,n2429);
    nand g985(n1110 ,n772 ,n835);
    or g986(n1450 ,n810 ,n1064);
    nor g987(n952 ,n392 ,n875);
    nor g988(n43 ,n2[32] ,n2[96]);
    nor g989(n180 ,n134 ,n179);
    nor g990(n814 ,n487 ,n805);
    nand g991(n2034 ,n4[38] ,n1469);
    not g992(n1288 ,n1160);
    nand g993(n2129 ,n2060 ,n2059);
    nor g994(n225 ,n53 ,n224);
    nand g995(n2230 ,n3[28] ,n1863);
    nor g996(n1366 ,n4[4] ,n1040);
    nor g997(n989 ,n396 ,n875);
    nand g998(n2177 ,n1982 ,n1971);
    dff g999(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n553), .Q(n8[21]));
    nor g1000(n1044 ,n8[31] ,n876);
    nand g1001(n2187 ,n2025 ,n2024);
    nand g1002(n1768 ,n4[13] ,n1485);
    nand g1003(n605 ,n6[2] ,n6[3]);
    not g1004(n323 ,n2[46]);
    nor g1005(n431 ,n8[22] ,n2345);
    dff g1006(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2113), .Q(n4[46]));
    not g1007(n1226 ,n1098);
    nor g1008(n179 ,n54 ,n178);
    not g1009(n313 ,n2[22]);
    dff g1010(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n601), .Q(n8[0]));
    nor g1011(n1998 ,n1534 ,n1316);
    nand g1012(n1031 ,n8[25] ,n877);
    or g1013(n1468 ,n810 ,n1054);
    nor g1014(n211 ,n30 ,n210);
    nand g1015(n1815 ,n5[35] ,n1645);
    not g1016(n1291 ,n1163);
    nor g1017(n1563 ,n5[43] ,n1014);
    nand g1018(n2135 ,n1738 ,n1737);
    nand g1019(n1969 ,n5[11] ,n1472);
    nor g1020(n1909 ,n1434 ,n1270);
    nor g1021(n1773 ,n1355 ,n1249);
    nor g1022(n461 ,n8[28] ,n2[124]);
    nor g1023(n252 ,n122 ,n251);
    nor g1024(n561 ,n290 ,n1);
    nor g1025(n1797 ,n1367 ,n1214);
    nor g1026(n230 ,n81 ,n229);
    nand g1027(n740 ,n8[9] ,n2[9]);
    nor g1028(n425 ,n8[21] ,n2[117]);
    nand g1029(n1167 ,n734 ,n907);
    dff g1030(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2313), .Q(n3[55]));
    nand g1031(n2168 ,n1925 ,n1923);
    nor g1032(n1386 ,n5[32] ,n1037);
    nor g1033(n378 ,n8[8] ,n2331);
    dff g1034(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2131), .Q(n5[50]));
    nor g1035(n826 ,n361 ,n271);
    nand g1036(n2194 ,n2039 ,n2031);
    nand g1037(n787 ,n8[28] ,n2[92]);
    dff g1038(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n560), .Q(n8[19]));
    nor g1039(n946 ,n352 ,n875);
    nor g1040(n835 ,n393 ,n805);
    nand g1041(n1578 ,n712 ,n996);
    dff g1042(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2186), .Q(n5[58]));
    dff g1043(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n538), .Q(n7[10]));
    not g1044(n1271 ,n1143);
    dff g1045(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2170), .Q(n5[17]));
    nor g1046(n1071 ,n8[7] ,n876);
    nor g1047(n1548 ,n3[19] ,n1023);
    nand g1048(n2174 ,n1953 ,n1951);
    nor g1049(n512 ,n8[16] ,n2371);
    nor g1050(n418 ,n8[27] ,n2[91]);
    nor g1051(n364 ,n8[23] ,n2378);
    dff g1052(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n586), .Q(n8[15]));
    not g1053(n318 ,n2[34]);
    nor g1054(n467 ,n8[16] ,n2339);
    not g1055(n1668 ,n1583);
    nand g1056(n1574 ,n761 ,n1000);
    xnor g1057(n2348 ,n87 ,n185);
    nand g1058(n786 ,n8[31] ,n2[95]);
    nor g1059(n371 ,n8[12] ,n2[76]);
    nand g1060(n2081 ,n1765 ,n1764);
    nor g1061(n1835 ,n1393 ,n1231);
    or g1062(n1458 ,n810 ,n1059);
    nand g1063(n2254 ,n3[4] ,n1887);
    nor g1064(n1434 ,n3[30] ,n1013);
    nand g1065(n2253 ,n3[5] ,n1886);
    or g1066(n1889 ,n1070 ,n1446);
    nor g1067(n957 ,n523 ,n875);
    nand g1068(n1598 ,n796 ,n975);
    not g1069(n1303 ,n1175);
    nand g1070(n2108 ,n1994 ,n1993);
    nor g1071(n964 ,n382 ,n875);
    xnor g1072(n99 ,n2[3] ,n2[67]);
    nand g1073(n1163 ,n727 ,n902);
    nor g1074(n594 ,n285 ,n1);
    nand g1075(n1837 ,n5[30] ,n1471);
    nand g1076(n656 ,n8[29] ,n2352);
    nor g1077(n58 ,n2[53] ,n2[117]);
    nor g1078(n831 ,n349 ,n804);
    nor g1079(n572 ,n288 ,n1);
    not g1080(n1281 ,n1153);
    nor g1081(n415 ,n8[20] ,n2[116]);
    nand g1082(n1594 ,n674 ,n979);
    nand g1083(n2204 ,n3[54] ,n1869);
    not g1084(n1255 ,n1127);
    dff g1085(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2175), .Q(n5[12]));
    dff g1086(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n578), .Q(n8[17]));
    nand g1087(n1142 ,n694 ,n881);
    nor g1088(n343 ,n8[24] ,n2[24]);
    nand g1089(n2418 ,n2405 ,n2411);
    nor g1090(n498 ,n8[4] ,n2[4]);
    nand g1091(n1581 ,n686 ,n993);
    nand g1092(n1178 ,n608 ,n919);
    nor g1093(n1496 ,n4[41] ,n1012);
    xnor g1094(n91 ,n2[1] ,n2[65]);
    xor g1095(n2323 ,n2[0] ,n2[64]);
    nor g1096(n525 ,n8[29] ,n2[29]);
    nor g1097(n888 ,n370 ,n805);
    or g1098(n1884 ,n1071 ,n1446);
    or g1099(n1460 ,n810 ,n1058);
    nor g1100(n1521 ,n4[56] ,n1029);
    nor g1101(n1545 ,n5[56] ,n1029);
    dff g1102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2084), .Q(n4[11]));
    nor g1103(n262 ,n6[1] ,n6[0]);
    nor g1104(n387 ,n2356 ,n10[1]);
    nor g1105(n486 ,n8[9] ,n2364);
    nor g1106(n1398 ,n5[29] ,n1035);
    nor g1107(n63 ,n2[27] ,n2[91]);
    nand g1108(n1608 ,n667 ,n964);
    not g1109(n1225 ,n1097);
    nor g1110(n156 ,n112 ,n155);
    nor g1111(n1361 ,n5[1] ,n1038);
    nor g1112(n217 ,n20 ,n216);
    or g1113(n1455 ,n810 ,n1069);
    not g1114(n1709 ,n1624);
    dff g1115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2177), .Q(n5[10]));
    nand g1116(n641 ,n8[11] ,n2334);
    dff g1117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2105), .Q(n4[54]));
    nand g1118(n1957 ,n5[12] ,n1644);
    or g1119(n1883 ,n1063 ,n1446);
    nor g1120(n48 ,n2[62] ,n2[126]);
    dff g1121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2140), .Q(n5[44]));
    or g1122(n1637 ,n807 ,n1071);
    nor g1123(n458 ,n8[4] ,n2327);
    nand g1124(n603 ,n8[9] ,n2332);
    nor g1125(n854 ,n424 ,n805);
    nand g1126(n1091 ,n638 ,n819);
    not g1127(n1204 ,n1076);
    nor g1128(n1519 ,n4[20] ,n1024);
    dff g1129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2125), .Q(n4[34]));
    nand g1130(n769 ,n8[27] ,n2382);
    nor g1131(n1499 ,n3[8] ,n1010);
    nand g1132(n2073 ,n1736 ,n1735);
    nand g1133(n2255 ,n3[3] ,n1888);
    nor g1134(n1917 ,n1440 ,n1275);
    dff g1135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n597), .Q(n7[27]));
    nor g1136(n1983 ,n1438 ,n1688);
    nand g1137(n1577 ,n722 ,n997);
    dff g1138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2143), .Q(n5[42]));
    or g1139(n140 ,n96 ,n139);
    nor g1140(n416 ,n8[13] ,n2[45]);
    not g1141(n1298 ,n1170);
    nand g1142(n1758 ,n4[16] ,n1476);
    nor g1143(n1042 ,n8[5] ,n876);
    nand g1144(n2127 ,n2054 ,n2053);
    nor g1145(n1498 ,n5[13] ,n1017);
    dff g1146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2114), .Q(n5[25]));
    nor g1147(n1970 ,n1340 ,n1683);
    nor g1148(n923 ,n430 ,n267);
    nor g1149(n1854 ,n1415 ,n1248);
    xnor g1150(n110 ,n2[9] ,n2[73]);
    nand g1151(n2259 ,n1907 ,n2227);
    dff g1152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2155), .Q(n5[32]));
    not g1153(n1694 ,n1609);
    dff g1154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2124), .Q(n4[35]));
    not g1155(n272 ,n1);
    not g1156(n339 ,n2387);
    nor g1157(n1896 ,n1423 ,n1258);
    nor g1158(n916 ,n501 ,n804);
    nor g1159(n39 ,n2[24] ,n2[88]);
    xnor g1160(n114 ,n2[11] ,n2[75]);
    nor g1161(n932 ,n341 ,n267);
    dff g1162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2316), .Q(n3[58]));
    nand g1163(n2248 ,n3[10] ,n1881);
    nor g1164(n937 ,n499 ,n267);
    not g1165(n1654 ,n1569);
    nand g1166(n801 ,n9[0] ,n798);
    nor g1167(n1630 ,n5[19] ,n1023);
    nor g1168(n1374 ,n4[1] ,n1038);
    nor g1169(n2030 ,n1545 ,n1233);
    or g1170(n1874 ,n1068 ,n1446);
    nand g1171(n1895 ,n5[25] ,n1480);
    nor g1172(n1857 ,n1418 ,n1252);
    nor g1173(n34 ,n2[13] ,n2[77]);
    nor g1174(n940 ,n504 ,n805);
    nor g1175(n376 ,n8[5] ,n2[69]);
    dff g1176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n581), .Q(n7[22]));
    not g1177(n1234 ,n1106);
    nor g1178(n2412 ,n2398 ,n7[24]);
    nor g1179(n192 ,n77 ,n191);
    nor g1180(n183 ,n14 ,n182);
    xnor g1181(n2383 ,n94 ,n255);
    or g1182(n1643 ,n807 ,n1052);
    nor g1183(n354 ,n8[19] ,n2[51]);
    nor g1184(n1428 ,n5[23] ,n1028);
    nor g1185(n489 ,n8[19] ,n2[83]);
    nand g1186(n1104 ,n652 ,n842);
    not g1187(n1699 ,n1614);
    nor g1188(n812 ,n496 ,n805);
    nor g1189(n514 ,n8[4] ,n2[100]);
    nand g1190(n1158 ,n721 ,n899);
    not g1191(n321 ,n2[36]);
    nand g1192(n661 ,n8[28] ,n2351);
    nor g1193(n474 ,n8[12] ,n2[12]);
    nand g1194(n1576 ,n735 ,n998);
    nor g1195(n596 ,n300 ,n1);
    dff g1196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2128), .Q(n4[31]));
    nor g1197(n1379 ,n4[8] ,n1010);
    nor g1198(n2011 ,n1405 ,n1296);
    not g1199(n1310 ,n1182);
    or g1200(n1472 ,n807 ,n1056);
    nor g1201(n861 ,n413 ,n271);
    nand g1202(n1749 ,n4[19] ,n1468);
    nand g1203(n756 ,n2[96] ,n10[0]);
    xnor g1204(n2357 ,n102 ,n203);
    nor g1205(n14 ,n2[23] ,n2[87]);
    nor g1206(n1836 ,n1395 ,n1234);
    nor g1207(n589 ,n334 ,n1);
    nand g1208(n791 ,n8[19] ,n2374);
    nand g1209(n1135 ,n687 ,n871);
    nand g1210(n2070 ,n1727 ,n1725);
    nand g1211(n803 ,n9[1] ,n798);
    nor g1212(n2059 ,n1558 ,n1712);
    or g1213(n1862 ,n1066 ,n1446);
    nand g1214(n1617 ,n718 ,n955);
    nor g1215(n463 ,n8[10] ,n2[42]);
    nand g1216(n1919 ,n5[20] ,n1475);
    nand g1217(n1145 ,n699 ,n884);
    nor g1218(n1534 ,n5[61] ,n1035);
    nor g1219(n476 ,n8[11] ,n2[11]);
    nor g1220(n902 ,n468 ,n804);
    nor g1221(n1522 ,n3[0] ,n1037);
    or g1222(n1866 ,n1061 ,n1446);
    or g1223(n1470 ,n810 ,n1042);
    nand g1224(n662 ,n8[16] ,n2[48]);
    nor g1225(n444 ,n8[18] ,n2[82]);
    nand g1226(n1021 ,n8[17] ,n877);
    nand g1227(n2273 ,n1932 ,n2241);
    nand g1228(n1115 ,n662 ,n850);
    nor g1229(n195 ,n12 ,n194);
    nor g1230(n441 ,n8[4] ,n2[36]);
    nor g1231(n1893 ,n1419 ,n1255);
    dff g1232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2302), .Q(n3[44]));
    nand g1233(n773 ,n2[97] ,n10[1]);
    not g1234(n297 ,n2[3]);
    nand g1235(n2091 ,n1800 ,n1799);
    nand g1236(n1180 ,n641 ,n923);
    nand g1237(n1567 ,n780 ,n1006);
    nor g1238(n1376 ,n4[0] ,n1037);
    nor g1239(n1762 ,n1563 ,n1208);
    nor g1240(n1805 ,n1514 ,n1680);
    nor g1241(n386 ,n8[23] ,n2[119]);
    nor g1242(n856 ,n365 ,n805);
    dff g1243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2314), .Q(n3[56]));
    nor g1244(n881 ,n383 ,n804);
    not g1245(n1206 ,n1078);
    nor g1246(n2019 ,n1535 ,n1700);
    nor g1247(n1541 ,n5[58] ,n1032);
    not g1248(n1696 ,n1611);
    xnor g1249(n2335 ,n115 ,n159);
    not g1250(n810 ,n809);
    xnor g1251(n2364 ,n126 ,n217);
    nor g1252(n1538 ,n4[46] ,n1018);
    nand g1253(n1088 ,n635 ,n823);
    nor g1254(n1372 ,n4[2] ,n1027);
    not g1255(n1263 ,n1135);
    nor g1256(n1806 ,n1372 ,n1676);
    nand g1257(n1027 ,n8[2] ,n877);
    nor g1258(n1344 ,n5[55] ,n1028);
    dff g1259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n583), .Q(n6[3]));
    nand g1260(n2244 ,n3[14] ,n1877);
    nor g1261(n2057 ,n1523 ,n1327);
    nand g1262(n1149 ,n707 ,n889);
    nor g1263(n566 ,n308 ,n1);
    nor g1264(n423 ,n8[31] ,n2386);
    dff g1265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2087), .Q(n4[8]));
    xnor g1266(n2344 ,n132 ,n177);
    xnor g1267(n2362 ,n120 ,n213);
    xnor g1268(n2360 ,n111 ,n209);
    xnor g1269(n2326 ,n99 ,n141);
    nand g1270(n1137 ,n696 ,n880);
    nor g1271(n168 ,n103 ,n167);
    nor g1272(n931 ,n533 ,n267);
    not g1273(n335 ,n2[30]);
    nand g1274(n2272 ,n1931 ,n2240);
    nor g1275(n1341 ,n4[37] ,n1039);
    nand g1276(n1176 ,n788 ,n918);
    nand g1277(n1607 ,n681 ,n965);
    nor g1278(n986 ,n376 ,n875);
    nor g1279(n798 ,n639 ,n605);
    nor g1280(n1948 ,n1494 ,n1299);
    nor g1281(n535 ,n289 ,n1);
    or g1282(n1476 ,n810 ,n1050);
    nand g1283(n2086 ,n1783 ,n1781);
    nor g1284(n1005 ,n515 ,n875);
    nor g1285(n1843 ,n1404 ,n1241);
    nor g1286(n205 ,n21 ,n204);
    nor g1287(n1002 ,n500 ,n875);
    nand g1288(n2283 ,n1950 ,n2251);
    nand g1289(n1020 ,n8[16] ,n877);
    nand g1290(n2245 ,n3[13] ,n1878);
    nor g1291(n414 ,n8[7] ,n2[39]);
    nor g1292(n844 ,n348 ,n805);
    nor g1293(n873 ,n431 ,n805);
    nand g1294(n2120 ,n1812 ,n2028);
    nor g1295(n1505 ,n3[6] ,n1011);
    nand g1296(n2178 ,n1988 ,n1987);
    not g1297(n1250 ,n1122);
    nor g1298(n1962 ,n1362 ,n1210);
    nor g1299(n541 ,n279 ,n1);
    nand g1300(n1906 ,n4[47] ,n1481);
    nand g1301(n2189 ,n2038 ,n2036);
    nand g1302(n2262 ,n1912 ,n2230);
    nand g1303(n2221 ,n3[37] ,n1886);
    nand g1304(n1611 ,n698 ,n962);
    or g1305(n1886 ,n1042 ,n1446);
    not g1306(n333 ,n2[42]);
    nand g1307(n1196 ,n627 ,n817);
    nand g1308(n735 ,n8[17] ,n2[81]);
    nor g1309(n402 ,n8[10] ,n2[74]);
    nor g1310(n863 ,n437 ,n804);
    nor g1311(n900 ,n464 ,n804);
    nor g1312(n559 ,n282 ,n1);
    nor g1313(n550 ,n314 ,n1);
    nand g1314(n1915 ,n5[21] ,n1467);
    dff g1315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n596), .Q(n8[31]));
    xnor g1316(n2352 ,n75 ,n193);
    nand g1317(n2172 ,n1943 ,n1936);
    nand g1318(n2068 ,n1718 ,n1716);
    nor g1319(n549 ,n274 ,n1);
    nor g1320(n1834 ,n1394 ,n1232);
    nand g1321(n776 ,n8[3] ,n2[99]);
    nand g1322(n2041 ,n4[36] ,n1474);
    not g1323(n289 ,n2[8]);
    nand g1324(n1035 ,n8[29] ,n877);
    nor g1325(n1904 ,n1431 ,n1267);
    nor g1326(n949 ,n497 ,n875);
    nor g1327(n2046 ,n1554 ,n1325);
    nand g1328(n796 ,n8[27] ,n2[123]);
    nor g1329(n23 ,n2[6] ,n2[70]);
    not g1330(n1276 ,n1148);
    not g1331(n1229 ,n1101);
    nor g1332(n1753 ,n1346 ,n1661);
    nand g1333(n653 ,n8[9] ,n2[73]);
    nand g1334(n2107 ,n1991 ,n1990);
    not g1335(n1235 ,n1107);
    nand g1336(n1109 ,n656 ,n844);
    nand g1337(n744 ,n8[24] ,n2[88]);
    nand g1338(n1734 ,n4[37] ,n1470);
    nor g1339(n41 ,n2[17] ,n2[81]);
    nor g1340(n981 ,n347 ,n875);
    nor g1341(n2408 ,n2390 ,n7[2]);
    nand g1342(n1087 ,n630 ,n822);
    nand g1343(n2049 ,n4[34] ,n1486);
    nand g1344(n614 ,n8[5] ,n2[101]);
    nand g1345(n2154 ,n1824 ,n1822);
    nand g1346(n2402 ,n7[14] ,n2393);
    nor g1347(n1536 ,n5[60] ,n1034);
    or g1348(n1489 ,n807 ,n1070);
    nor g1349(n1518 ,n4[58] ,n1032);
    xnor g1350(n105 ,n2[57] ,n2[121]);
    nor g1351(n938 ,n398 ,n267);
    nor g1352(n799 ,n9[0] ,n798);
    nor g1353(n1554 ,n5[6] ,n1011);
    nor g1354(n1735 ,n1531 ,n1656);
    nor g1355(n1947 ,n1497 ,n1300);
    or g1356(n1462 ,n810 ,n1073);
    or g1357(n1865 ,n1062 ,n1446);
    nor g1358(n359 ,n8[26] ,n2[26]);
    nand g1359(n2203 ,n3[55] ,n1868);
    nand g1360(n1147 ,n618 ,n888);
    not g1361(n1213 ,n1085);
    nand g1362(n1602 ,n713 ,n970);
    nor g1363(n1987 ,n1412 ,n1315);
    nor g1364(n822 ,n381 ,n267);
    not g1365(n2390 ,n7[3]);
    nor g1366(n1043 ,n8[6] ,n876);
    nor g1367(n560 ,n281 ,n1);
    nor g1368(n1392 ,n3[55] ,n1028);
    nand g1369(n655 ,n8[29] ,n2[61]);
    nand g1370(n611 ,n8[6] ,n2[102]);
    nor g1371(n56 ,n2[46] ,n2[110]);
    dff g1372(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2115), .Q(n4[44]));
    nand g1373(n1978 ,n4[28] ,n1650);
    nor g1374(n1491 ,n3[12] ,n1015);
    nor g1375(n1719 ,n1562 ,n1310);
    nor g1376(n956 ,n509 ,n269);
    nor g1377(n532 ,n8[21] ,n2[53]);
    nor g1378(n1340 ,n4[59] ,n1033);
    nor g1379(n1442 ,n4[40] ,n1010);
    nor g1380(n523 ,n8[10] ,n2[106]);
    nor g1381(n1851 ,n1413 ,n1247);
    nor g1382(n598 ,n335 ,n1);
    nor g1383(n2016 ,n1397 ,n1699);
    nor g1384(n1516 ,n3[1] ,n1038);
    not g1385(n1686 ,n1601);
    nor g1386(n366 ,n8[14] ,n2[46]);
    nor g1387(n352 ,n8[30] ,n2[94]);
    nor g1388(n1370 ,n4[38] ,n1011);
    nor g1389(n1506 ,n4[53] ,n1025);
    nand g1390(n639 ,n6[0] ,n6[1]);
    dff g1391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2109), .Q(n4[50]));
    nand g1392(n637 ,n8[2] ,n2357);
    nand g1393(n701 ,n8[14] ,n2[78]);
    nand g1394(n689 ,n8[5] ,n2[5]);
    nand g1395(n2276 ,n1940 ,n2245);
    nor g1396(n1924 ,n1565 ,n1281);
    nand g1397(n2097 ,n1961 ,n1805);
    nor g1398(n928 ,n344 ,n804);
    nand g1399(n2271 ,n1929 ,n2239);
    nor g1400(n169 ,n16 ,n168);
    xnor g1401(n134 ,n2[22] ,n2[86]);
    nor g1402(n421 ,n8[23] ,n2346);
    not g1403(n1246 ,n1118);
    nor g1404(n158 ,n114 ,n157);
    nor g1405(n977 ,n531 ,n875);
    dff g1406(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n562), .Q(n8[18]));
    not g1407(n1309 ,n1181);
    nand g1408(n2184 ,n2012 ,n2011);
    dff g1409(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2260), .Q(n3[30]));
    nor g1410(n1047 ,n8[13] ,n876);
    nor g1411(n238 ,n117 ,n237);
    not g1412(n301 ,n2[41]);
    nand g1413(n657 ,n8[8] ,n2363);
    dff g1414(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n574), .Q(n7[16]));
    xnor g1415(n82 ,n2[26] ,n2[90]);
    nor g1416(n968 ,n425 ,n875);
    nor g1417(n493 ,n8[20] ,n2[84]);
    nand g1418(n2136 ,n1746 ,n1745);
    dff g1419(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2112), .Q(n4[47]));
    xnor g1420(n2361 ,n116 ,n211);
    nor g1421(n1396 ,n4[51] ,n1023);
    not g1422(n299 ,n2[2]);
    dff g1423(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2095), .Q(n4[0]));
    dff g1424(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2182), .Q(n5[60]));
    dff g1425(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2304), .Q(n3[46]));
    nor g1426(n926 ,n433 ,n804);
    nand g1427(n774 ,n8[2] ,n2[98]);
    nor g1428(n1060 ,n8[24] ,n876);
    or g1429(n1873 ,n1053 ,n1446);
    nand g1430(n1008 ,n876 ,n804);
    or g1431(n1861 ,n1067 ,n1446);
    xnor g1432(n2368 ,n78 ,n225);
    nand g1433(n642 ,n8[8] ,n2[72]);
    or g1434(n1452 ,n810 ,n1051);
    nor g1435(n850 ,n519 ,n271);
    nor g1436(n1347 ,n5[44] ,n1015);
    nor g1437(n586 ,n294 ,n1);
    nor g1438(n862 ,n414 ,n804);
    nor g1439(n150 ,n107 ,n149);
    nor g1440(n1932 ,n1526 ,n1288);
    nor g1441(n869 ,n417 ,n804);
    nand g1442(n2027 ,n4[40] ,n1453);
    dff g1443(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2090), .Q(n4[5]));
    nor g1444(n889 ,n447 ,n804);
    nand g1445(n2205 ,n3[53] ,n1870);
    not g1446(n1292 ,n1164);
    not g1447(n288 ,n2[5]);
    not g1448(n1656 ,n1571);
    not g1449(n292 ,n2[4]);
    nand g1450(n2280 ,n1946 ,n2248);
    nor g1451(n1513 ,n4[63] ,n1036);
    nor g1452(n479 ,n8[22] ,n2377);
    nand g1453(n1858 ,n5[42] ,n1641);
    dff g1454(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2144), .Q(n5[41]));
    not g1455(n1682 ,n1597);
    nor g1456(n1348 ,n4[16] ,n1020);
    dff g1457(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n576), .Q(n8[29]));
    nor g1458(n1902 ,n1428 ,n1264);
    nor g1459(n1529 ,n5[62] ,n1013);
    nor g1460(n1725 ,n1334 ,n1653);
    nand g1461(n2195 ,n3[63] ,n1860);
    nor g1462(n1413 ,n3[44] ,n1015);
    not g1463(n306 ,n2[57]);
    not g1464(n1710 ,n1625);
    nor g1465(n985 ,n483 ,n269);
    nor g1466(n216 ,n95 ,n215);
    xnor g1467(n126 ,n2[41] ,n2[105]);
    nand g1468(n695 ,n8[29] ,n2[29]);
    nand g1469(n2281 ,n1947 ,n2249);
    nor g1470(n1401 ,n4[45] ,n1017);
    nor g1471(n1911 ,n1435 ,n1272);
    nor g1472(n1967 ,n1356 ,n1682);
    nand g1473(n2299 ,n1857 ,n2217);
    dff g1474(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2146), .Q(n5[40]));
    nor g1475(n1542 ,n3[18] ,n1022);
    nor g1476(n1426 ,n3[35] ,n1016);
    nor g1477(n898 ,n470 ,n804);
    xnor g1478(n2334 ,n114 ,n157);
    not g1479(n807 ,n806);
    nand g1480(n1626 ,n786 ,n947);
    nand g1481(n677 ,n8[8] ,n2[40]);
    nor g1482(n2013 ,n1388 ,n1698);
    nand g1483(n1095 ,n644 ,n834);
    nor g1484(n1901 ,n1427 ,n1263);
    not g1485(n1249 ,n1121);
    nand g1486(n2163 ,n1900 ,n1898);
    nor g1487(n399 ,n8[31] ,n2354);
    nor g1488(n455 ,n8[11] ,n2366);
    nor g1489(n1810 ,n1374 ,n1677);
    nor g1490(n1916 ,n1441 ,n1276);
    nor g1491(n1427 ,n3[34] ,n1027);
    nor g1492(n564 ,n320 ,n1);
    xnor g1493(n122 ,n2[58] ,n2[122]);
    nand g1494(n618 ,n8[20] ,n2343);
    nand g1495(n72 ,n2[2] ,n2[66]);
    nor g1496(n513 ,n8[5] ,n2[5]);
    nand g1497(n1161 ,n725 ,n903);
    nor g1498(n1406 ,n3[48] ,n1020);
    dff g1499(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2263), .Q(n3[27]));
    nand g1500(n751 ,n8[20] ,n2[84]);
    nand g1501(n1982 ,n5[10] ,n1641);
    nor g1502(n505 ,n8[9] ,n2[73]);
    nor g1503(n456 ,n8[20] ,n2[20]);
    nand g1504(n2087 ,n1786 ,n1785);
    dff g1505(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2280), .Q(n3[10]));
    not g1506(n1300 ,n1172);
    nor g1507(n71 ,n2[59] ,n2[123]);
    not g1508(n1241 ,n1113);
    not g1509(n2391 ,n7[19]);
    nor g1510(n1399 ,n3[52] ,n1024);
    nor g1511(n1391 ,n3[56] ,n1029);
    nor g1512(n972 ,n362 ,n875);
    nand g1513(n1770 ,n5[26] ,n1483);
    dff g1514(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2089), .Q(n4[6]));
    nor g1515(n915 ,n438 ,n804);
    nand g1516(n700 ,n8[8] ,n2[8]);
    not g1517(n1251 ,n1123);
    dff g1518(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n566), .Q(n7[1]));
    nand g1519(n944 ,n943 ,n875);
    nand g1520(n749 ,n8[30] ,n2[94]);
    nor g1521(n2400 ,n7[31] ,n7[30]);
    dff g1522(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2269), .Q(n3[21]));
    nor g1523(n1565 ,n3[22] ,n1026);
    nand g1524(n737 ,n8[14] ,n2337);
    or g1525(n1864 ,n1064 ,n1446);
    nand g1526(n2146 ,n1782 ,n1780);
    nand g1527(n763 ,n8[29] ,n2[125]);
    not g1528(n302 ,n2[16]);
    nand g1529(n783 ,n8[25] ,n2[57]);
    nor g1530(n426 ,n2[33] ,n10[1]);
    not g1531(n1659 ,n1574);
    nor g1532(n553 ,n319 ,n1);
    dff g1533(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2283), .Q(n3[7]));
    nor g1534(n1431 ,n3[32] ,n1037);
    nand g1535(n2132 ,n1724 ,n1722);
    not g1536(n92 ,n91);
    nor g1537(n189 ,n60 ,n188);
    nand g1538(n1195 ,n778 ,n825);
    not g1539(n1323 ,n1195);
    nand g1540(n2196 ,n3[62] ,n1861);
    nor g1541(n524 ,n8[3] ,n2[99]);
    nor g1542(n1796 ,n1365 ,n1673);
    nor g1543(n1492 ,n3[11] ,n1014);
    nor g1544(n1774 ,n1414 ,n1667);
    nand g1545(n2218 ,n3[40] ,n1883);
    nand g1546(n672 ,n8[26] ,n2349);
    nor g1547(n847 ,n527 ,n271);
    nand g1548(n1018 ,n8[14] ,n877);
    nor g1549(n57 ,n2[22] ,n2[86]);
    not g1550(n1254 ,n1126);
    nand g1551(n2160 ,n1852 ,n1850);
    nor g1552(n381 ,n8[4] ,n2359);
    dff g1553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2073), .Q(n4[22]));
    nand g1554(n2251 ,n3[7] ,n1884);
    dff g1555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n580), .Q(n6[1]));
    nor g1556(n508 ,n8[15] ,n2[47]);
    nor g1557(n573 ,n304 ,n1);
    nand g1558(n1733 ,n4[23] ,n1458);
    not g1559(n1712 ,n1627);
    nor g1560(n65 ,n2[60] ,n2[124]);
    nand g1561(n617 ,n8[6] ,n2[70]);
    nor g1562(n1543 ,n5[57] ,n1031);
    nand g1563(n1075 ,n610 ,n931);
    nand g1564(n654 ,n2[32] ,n10[0]);
    nor g1565(n1073 ,n8[21] ,n876);
    nor g1566(n1923 ,n1630 ,n1279);
    dff g1567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2121), .Q(n4[38]));
    nand g1568(n2242 ,n3[16] ,n1875);
    nand g1569(n2231 ,n3[27] ,n1864);
    nand g1570(n2212 ,n3[46] ,n1877);
    nor g1571(n2061 ,n1561 ,n1713);
    nor g1572(n593 ,n332 ,n1);
    nor g1573(n221 ,n27 ,n220);
    nor g1574(n599 ,n286 ,n1);
    dff g1575(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2295), .Q(n3[37]));
    dff g1576(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n551), .Q(n8[20]));
    not g1577(n1208 ,n1080);
    nor g1578(n191 ,n63 ,n190);
    nor g1579(n865 ,n427 ,n804);
    nor g1580(n588 ,n312 ,n1);
    nor g1581(n203 ,n19 ,n202);
    nand g1582(n2164 ,n1905 ,n1902);
    dff g1583(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2290), .Q(n3[0]));
    dff g1584(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2178), .Q(n5[63]));
    nor g1585(n1899 ,n1426 ,n1261);
    nand g1586(n2307 ,n1843 ,n2209);
    xnor g1587(n2358 ,n89 ,n205);
    nand g1588(n1146 ,n702 ,n886);
    nand g1589(n1589 ,n625 ,n985);
    nand g1590(n2197 ,n3[61] ,n1862);
    nand g1591(n2319 ,n1821 ,n2197);
    nor g1592(n2427 ,n2415 ,n2426);
    nand g1593(n2175 ,n1957 ,n1955);
    nand g1594(n2201 ,n3[57] ,n1866);
    nor g1595(n209 ,n35 ,n208);
    xnor g1596(n88 ,n2[32] ,n2[96]);
    nor g1597(n509 ,n8[9] ,n2[105]);
    nor g1598(n370 ,n8[20] ,n2343);
    nand g1599(n1034 ,n8[28] ,n877);
    dff g1600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2264), .Q(n3[26]));
    dff g1601(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2159), .Q(n5[28]));
    not g1602(n290 ,n2[28]);
    nor g1603(n1056 ,n8[11] ,n876);
    not g1604(n1708 ,n1623);
    nand g1605(n2192 ,n2058 ,n2057);
    nand g1606(n2410 ,n7[5] ,n7[4]);
    nor g1607(n1062 ,n8[26] ,n876);
    nor g1608(n2055 ,n1557 ,n1711);
    nor g1609(n1562 ,n5[5] ,n1039);
    nor g1610(n884 ,n374 ,n271);
    nand g1611(n2042 ,n5[54] ,n1465);
    xnor g1612(n75 ,n2[29] ,n2[93]);
    nor g1613(n1378 ,n5[34] ,n1027);
    dff g1614(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2190), .Q(n5[54]));
    nor g1615(n846 ,n480 ,n804);
    or g1616(n1881 ,n1045 ,n1446);
    nand g1617(n2130 ,n2062 ,n2061);
    nand g1618(n2090 ,n1798 ,n1796);
    nand g1619(n604 ,n8[30] ,n2[62]);
    nand g1620(n729 ,n8[24] ,n2379);
    or g1621(n1453 ,n810 ,n1063);
    nand g1622(n1150 ,n709 ,n890);
    nand g1623(n733 ,n8[15] ,n2338);
    nor g1624(n13 ,n2[55] ,n2[119]);
    not g1625(n1671 ,n1586);
    nand g1626(n1572 ,n758 ,n1001);
    nor g1627(n2035 ,n1341 ,n1705);
    not g1628(n1267 ,n1139);
    not g1629(n275 ,n2[52]);
    not g1630(n1274 ,n1146);
    nor g1631(n1514 ,n4[62] ,n1013);
    or g1632(n1447 ,n810 ,n1045);
    not g1633(n1316 ,n1188);
    nor g1634(n1355 ,n5[41] ,n1012);
    not g1635(n1700 ,n1615);
    or g1636(n15 ,n2[1] ,n2[65]);
    dff g1637(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2074), .Q(n4[21]));
    nand g1638(n2037 ,n5[6] ,n1635);
    not g1639(n1287 ,n1159);
    nand g1640(n2314 ,n1831 ,n2202);
    nand g1641(n663 ,n8[20] ,n2[116]);
    nor g1642(n883 ,n525 ,n804);
    nor g1643(n1747 ,n1343 ,n1206);
    nor g1644(n54 ,n2[21] ,n2[85]);
    nand g1645(n1761 ,n4[15] ,n1481);
    nand g1646(n1583 ,n784 ,n991);
    nand g1647(n2155 ,n1826 ,n1827);
    nand g1648(n1090 ,n604 ,n829);
    not g1649(n315 ,n2[61]);
    nor g1650(n32 ,n2[54] ,n2[118]);
    nor g1651(n2403 ,n7[29] ,n7[28]);
    or g1652(n1870 ,n1073 ,n1446);
    nor g1653(n1373 ,n4[7] ,n1030);
    nor g1654(n1559 ,n3[21] ,n1025);
    nand g1655(n716 ,n8[18] ,n2341);
    dff g1656(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2075), .Q(n4[20]));
    nor g1657(n147 ,n22 ,n146);
    nor g1658(n849 ,n401 ,n267);
    nand g1659(n1569 ,n744 ,n1004);
    nand g1660(n2199 ,n3[59] ,n1864);
    nor g1661(n577 ,n328 ,n1);
    nand g1662(n1593 ,n636 ,n981);
    not g1663(n1264 ,n1136);
    nand g1664(n2216 ,n3[42] ,n1881);
    nand g1665(n686 ,n8[12] ,n2[76]);
    dff g1666(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n594), .Q(n7[24]));
    nand g1667(n1614 ,n679 ,n958);
    nand g1668(n631 ,n8[21] ,n2[53]);
    not g1669(n1312 ,n1184);
    xnor g1670(n2376 ,n128 ,n241);
    nor g1671(n196 ,n80 ,n195);
    nor g1672(n988 ,n355 ,n875);
    nor g1673(n894 ,n517 ,n805);
    not g1674(n1220 ,n1092);
    nand g1675(n1188 ,n738 ,n860);
    dff g1676(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n590), .Q(n7[18]));
    or g1677(n1875 ,n1050 ,n1446);
    or g1678(n1451 ,n810 ,n1062);
    nor g1679(n1935 ,n1525 ,n1290);
    nor g1680(n1764 ,n1350 ,n1664);
    nand g1681(n1138 ,n658 ,n872);
    nor g1682(n879 ,n432 ,n804);
    not g1683(n327 ,n2[31]);
    nor g1684(n1362 ,n3[2] ,n1027);
    nor g1685(n878 ,n378 ,n805);
    nor g1686(n954 ,n506 ,n269);
    dff g1687(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2176), .Q(n5[11]));
    nand g1688(n1019 ,n8[15] ,n877);
    not g1689(n1202 ,n1074);
    nor g1690(n919 ,n448 ,n267);
    nand g1691(n690 ,n8[22] ,n2345);
    xnor g1692(n86 ,n2[24] ,n2[88]);
    xnor g1693(n107 ,n2[7] ,n2[71]);
    nor g1694(n1557 ,n4[31] ,n1036);
    nand g1695(n2161 ,n1770 ,n1856);
    nand g1696(n708 ,n8[11] ,n2366);
    nand g1697(n2190 ,n2042 ,n2045);
    nand g1698(n1085 ,n745 ,n821);
    nand g1699(n1613 ,n648 ,n959);
    nor g1700(n941 ,n479 ,n805);
    nor g1701(n145 ,n70 ,n144);
    nor g1702(n860 ,n439 ,n805);
    nor g1703(n600 ,n317 ,n1);
    nand g1704(n706 ,n8[19] ,n2[115]);
    nand g1705(n1164 ,n730 ,n904);
    dff g1706(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2157), .Q(n5[30]));
    not g1707(n2394 ,n7[16]);
    nand g1708(n2021 ,n5[8] ,n1639);
    or g1709(n1459 ,n810 ,n1071);
    not g1710(n1245 ,n1117);
    not g1711(n1714 ,n1629);
    nand g1712(n1984 ,n4[54] ,n1460);
    nor g1713(n1927 ,n1559 ,n1282);
    not g1714(n1262 ,n1134);
    nor g1715(n1375 ,n5[35] ,n1016);
    nor g1716(n1814 ,n1376 ,n1678);
    dff g1717(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2168), .Q(n5[19]));
    nand g1718(n615 ,n8[28] ,n2[124]);
    nor g1719(n1931 ,n1542 ,n1286);
    nor g1720(n970 ,n386 ,n269);
    nand g1721(n668 ,n8[14] ,n2[46]);
    nor g1722(n448 ,n8[12] ,n2335);
    nor g1723(n1339 ,n5[46] ,n1018);
    nand g1724(n2290 ,n1979 ,n2210);
    nor g1725(n1502 ,n5[15] ,n1019);
    nor g1726(n2063 ,n1560 ,n1328);
    not g1727(n328 ,n2[56]);
    not g1728(n1706 ,n1621);
    nor g1729(n236 ,n109 ,n235);
    nor g1730(n484 ,n8[31] ,n2[95]);
    xnor g1731(n106 ,n2[48] ,n2[112]);
    nand g1732(n2103 ,n1977 ,n2066);
    not g1733(n1691 ,n1606);
    nor g1734(n955 ,n452 ,n875);
    nand g1735(n2420 ,n2400 ,n2403);
    nand g1736(n2267 ,n1922 ,n2235);
    not g1737(n281 ,n2[51]);
    nor g1738(n175 ,n47 ,n174);
    nor g1739(n430 ,n8[11] ,n2334);
    nand g1740(n1784 ,n5[0] ,n1457);
    nand g1741(n2077 ,n1751 ,n1750);
    dff g1742(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2274), .Q(n3[32]));
    nand g1743(n1131 ,n754 ,n868);
    nor g1744(n1552 ,n4[33] ,n1038);
    nand g1745(n1832 ,n5[31] ,n1449);
    nor g1746(n1737 ,n1337 ,n1203);
    nand g1747(n2054 ,n4[32] ,n1455);
    nand g1748(n2241 ,n3[17] ,n1890);
    dff g1749(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2158), .Q(n5[29]));
    nor g1750(n210 ,n111 ,n209);
    nand g1751(n806 ,n272 ,n803);
    xnor g1752(n2385 ,n90 ,n259);
    nor g1753(n451 ,n8[22] ,n2[22]);
    nor g1754(n17 ,n2[48] ,n2[112]);
    nand g1755(n2210 ,n3[0] ,n1859);
    not g1756(n1320 ,n1192);
    dff g1757(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n595), .Q(n8[14]));
    nand g1758(n73 ,n2[0] ,n2[64]);
    nor g1759(n1441 ,n3[26] ,n1032);
    nor g1760(n437 ,n8[6] ,n2[38]);
    dff g1761(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2108), .Q(n4[51]));
    not g1762(n1693 ,n1608);
    not g1763(n1688 ,n1603);
    not g1764(n2397 ,n7[27]);
    nand g1765(n2223 ,n3[35] ,n1888);
    nand g1766(n1618 ,n665 ,n954);
    not g1767(n1695 ,n1610);
    not g1768(n1209 ,n1081);
    nand g1769(n1132 ,n616 ,n885);
    nand g1770(n613 ,n8[12] ,n2367);
    nand g1771(n1148 ,n704 ,n887);
    nand g1772(n626 ,n2356 ,n10[1]);
    nor g1773(n488 ,n8[30] ,n2[126]);
    dff g1774(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2082), .Q(n4[13]));
    dff g1775(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2318), .Q(n3[60]));
    nor g1776(n980 ,n454 ,n269);
    or g1777(n1878 ,n1047 ,n1446);
    nor g1778(n204 ,n102 ,n203);
    nor g1779(n18 ,n2[15] ,n2[79]);
    nor g1780(n983 ,n357 ,n875);
    nand g1781(n2162 ,n2010 ,n2009);
    nor g1782(n424 ,n8[26] ,n2349);
    nand g1783(n2180 ,n2001 ,n1998);
    nand g1784(n1166 ,n732 ,n905);
    nor g1785(n563 ,n277 ,n1);
    nor g1786(n1351 ,n5[42] ,n1041);
    not g1787(n1280 ,n1152);
    nor g1788(n1956 ,n1510 ,n1307);
    or g1789(n1456 ,n810 ,n1060);
    nand g1790(n1200 ,n791 ,n939);
    nor g1791(n925 ,n416 ,n804);
    nor g1792(n1855 ,n1417 ,n1250);
    nand g1793(n1605 ,n663 ,n967);
    nand g1794(n648 ,n8[12] ,n2[108]);
    nor g1795(n347 ,n2[64] ,n10[0]);
    nand g1796(n644 ,n8[27] ,n2[59]);
    nor g1797(n174 ,n129 ,n173);
    dff g1798(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2192), .Q(n5[52]));
    nand g1799(n2296 ,n1894 ,n2220);
    nand g1800(n674 ,n8[31] ,n2[127]);
    nand g1801(n635 ,n8[3] ,n2358);
    xnor g1802(n136 ,n2[6] ,n2[70]);
    dff g1803(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2069), .Q(n4[26]));
    nor g1804(n557 ,n299 ,n1);
    nand g1805(n1126 ,n680 ,n862);
    nor g1806(n1945 ,n1492 ,n1297);
    dff g1807(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2110), .Q(n4[49]));
    nand g1808(n2104 ,n1981 ,n1980);
    nand g1809(n2038 ,n5[55] ,n1463);
    nor g1810(n472 ,n8[15] ,n2338);
    nor g1811(n936 ,n522 ,n267);
    or g1812(n1888 ,n1072 ,n1446);
    nand g1813(n2083 ,n1772 ,n1771);
    nor g1814(n377 ,n2323 ,n10[0]);
    nor g1815(n910 ,n481 ,n804);
    nor g1816(n892 ,n384 ,n805);
    dff g1817(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2289), .Q(n3[1]));
    nand g1818(n2207 ,n3[51] ,n1872);
    nand g1819(n780 ,n8[26] ,n2[90]);
    nor g1820(n551 ,n275 ,n1);
    nand g1821(n2289 ,n1966 ,n2257);
    nor g1822(n1369 ,n4[3] ,n1016);
    not g1823(n1217 ,n1089);
    not g1824(n284 ,n2[49]);
    nand g1825(n2252 ,n3[6] ,n1885);
    nor g1826(n198 ,n83 ,n197);
    not g1827(n1707 ,n1622);
    nand g1828(n1010 ,n8[8] ,n877);
    nor g1829(n1556 ,n4[32] ,n1037);
    xnor g1830(n2386 ,n74 ,n261);
    dff g1831(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n591), .Q(n8[11]));
    nor g1832(n891 ,n450 ,n804);
    nand g1833(n753 ,n8[9] ,n2[105]);
    xnor g1834(n76 ,n2[46] ,n2[110]);
    xnor g1835(n2371 ,n106 ,n231);
    nor g1836(n374 ,n8[28] ,n2[28]);
    nand g1837(n1960 ,n4[63] ,n1482);
    nor g1838(n851 ,n508 ,n271);
    nor g1839(n234 ,n98 ,n233);
    nand g1840(n2293 ,n1899 ,n2223);
    nor g1841(n993 ,n371 ,n875);
    nor g1842(n406 ,n8[14] ,n2[110]);
    nor g1843(n1430 ,n4[13] ,n1017);
    nand g1844(n709 ,n8[24] ,n2[24]);
    nand g1845(n1089 ,n619 ,n824);
    nand g1846(n697 ,n8[15] ,n2[111]);
    nor g1847(n344 ,n2[0] ,n10[0]);
    nand g1848(n1086 ,n621 ,n820);
    dff g1849(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2152), .Q(n5[35]));
    dff g1850(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2134), .Q(n5[48]));
    not g1851(n309 ,n2[10]);
    not g1852(n1297 ,n1169);
    nand g1853(n1028 ,n8[23] ,n877);
    or g1854(n1479 ,n810 ,n1048);
    nand g1855(n2113 ,n2008 ,n2007);
    nor g1856(n35 ,n2[36] ,n2[100]);
    not g1857(n1308 ,n1180);
    nand g1858(n1776 ,n5[41] ,n1640);
    nand g1859(n2147 ,n1788 ,n1787);
    nor g1860(n907 ,n474 ,n804);
    not g1861(n1221 ,n1093);
    not g1862(n331 ,n2[9]);
    nand g1863(n2093 ,n1808 ,n1806);
    nor g1864(n821 ,n485 ,n805);
    nor g1865(n384 ,n8[19] ,n2342);
    nor g1866(n887 ,n359 ,n271);
    nand g1867(n2088 ,n1790 ,n1789);
    nand g1868(n804 ,n568 ,n800);
    not g1869(n1237 ,n1109);
    not g1870(n1662 ,n1577);
    nor g1871(n393 ,n8[26] ,n2381);
    nor g1872(n880 ,n434 ,n805);
    nand g1873(n1622 ,n776 ,n950);
    nor g1874(n866 ,n389 ,n267);
    nand g1875(n703 ,n8[21] ,n2[117]);
    nor g1876(n227 ,n26 ,n226);
    nand g1877(n1606 ,n706 ,n966);
    nand g1878(n620 ,n8[20] ,n2[52]);
    nor g1879(n1389 ,n3[57] ,n1031);
    xnor g1880(n2369 ,n76 ,n227);
    nand g1881(n772 ,n8[26] ,n2381);
    nand g1882(n2159 ,n1848 ,n1845);
    xnor g1883(n2349 ,n82 ,n187);
    nand g1884(n731 ,n2355 ,n10[0]);
    not g1885(n2393 ,n7[15]);
    or g1886(n1636 ,n807 ,n1042);
    nor g1887(n404 ,n8[30] ,n2385);
    nand g1888(n723 ,n8[17] ,n2[17]);
    nand g1889(n1566 ,n779 ,n1007);
    nor g1890(n237 ,n28 ,n236);
    nand g1891(n1157 ,n719 ,n898);
    nand g1892(n607 ,n8[31] ,n2[63]);
    nand g1893(n1012 ,n8[9] ,n877);
    dff g1894(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2307), .Q(n3[49]));
    nor g1895(n439 ,n8[29] ,n2384);
    not g1896(n1243 ,n1115);
    nor g1897(n996 ,n459 ,n875);
    or g1898(n1648 ,n807 ,n1048);
    dff g1899(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2293), .Q(n3[35]));
    not g1900(n1667 ,n1582);
    not g1901(n1238 ,n1110);
    nand g1902(n705 ,n8[28] ,n2383);
    nor g1903(n1785 ,n1379 ,n1670);
    nand g1904(n2166 ,n1915 ,n1913);
    nor g1905(n1537 ,n4[47] ,n1019);
    not g1906(n1294 ,n1166);
    nand g1907(n2158 ,n1842 ,n1840);
    or g1908(n1880 ,n1056 ,n1446);
    nor g1909(n22 ,n2[5] ,n2[69]);
    dff g1910(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2101), .Q(n4[58]));
    nand g1911(n1972 ,n4[59] ,n1450);
    nand g1912(n2292 ,n1901 ,n2224);
    nor g1913(n208 ,n108 ,n207);
    dff g1914(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n592), .Q(n7[20]));
    nand g1915(n1197 ,n782 ,n936);
    dff g1916(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2180), .Q(n5[61]));
    nand g1917(n2124 ,n2044 ,n2043);
    nor g1918(n1892 ,n1421 ,n1254);
    nand g1919(n1597 ,n615 ,n976);
    nor g1920(n368 ,n8[3] ,n2[67]);
    nand g1921(n758 ,n8[21] ,n2[85]);
    nand g1922(n2029 ,n4[43] ,n1487);
    dff g1923(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2126), .Q(n4[33]));
    not g1924(n2396 ,n7[6]);
    nand g1925(n1077 ,n771 ,n812);
    nand g1926(n768 ,n8[16] ,n2[112]);
    nor g1927(n1343 ,n5[45] ,n1017);
    xnor g1928(n2337 ,n119 ,n163);
    or g1929(n1887 ,n1057 ,n1446);
    nor g1930(n967 ,n415 ,n875);
    not g1931(n307 ,n2[18]);
    xnor g1932(n111 ,n2[37] ,n2[101]);
    nand g1933(n1193 ,n777 ,n917);
    nand g1934(n2170 ,n1934 ,n1933);
    nand g1935(n1185 ,n755 ,n927);
    nor g1936(n1332 ,n4[27] ,n1033);
    xnor g1937(n83 ,n2[31] ,n2[95]);
    dff g1938(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n570), .Q(n8[4]));
    or g1939(n1478 ,n810 ,n1072);
    nor g1940(n1844 ,n1406 ,n1243);
    nor g1941(n60 ,n2[26] ,n2[90]);
    or g1942(n805 ,n569 ,n803);
    not g1943(n1689 ,n1604);
    nor g1944(n1781 ,n1359 ,n1669);
    nand g1945(n2051 ,n4[33] ,n1490);
    nand g1946(n1910 ,n5[22] ,n1465);
    nor g1947(n1435 ,n3[29] ,n1035);
    nor g1948(n2031 ,n1547 ,n1321);
    nand g1949(n1763 ,n5[43] ,n1472);
    nand g1950(n2227 ,n3[31] ,n1860);
    nor g1951(n558 ,n331 ,n1);
    nand g1952(n1934 ,n5[17] ,n1643);
    nor g1953(n1532 ,n5[17] ,n1021);
    nor g1954(n933 ,n356 ,n805);
    nor g1955(n392 ,n8[5] ,n2[101]);
    nand g1956(n2409 ,n7[23] ,n2392);
    nor g1957(n1438 ,n4[54] ,n1026);
    nor g1958(n1352 ,n5[2] ,n1027);
    xnor g1959(n101 ,n2[4] ,n2[68]);
    nor g1960(n592 ,n287 ,n1);
    not g1961(n1268 ,n1140);
    nor g1962(n207 ,n50 ,n206);
    nand g1963(n2209 ,n3[49] ,n1890);
    nor g1964(n350 ,n8[10] ,n2333);
    nand g1965(n2106 ,n1986 ,n1985);
    nor g1966(n2015 ,n1539 ,n1317);
    xnor g1967(n93 ,n2[56] ,n2[120]);
    nor g1968(n1958 ,n1512 ,n1309);
    dff g1969(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2122), .Q(n4[37]));
    or g1970(n1457 ,n807 ,n1069);
    nand g1971(n1624 ,n773 ,n949);
    nor g1972(n181 ,n57 ,n180);
    nor g1973(n64 ,n2[11] ,n2[75]);
    nor g1974(n459 ,n8[15] ,n2[79]);
    nand g1975(n1730 ,n5[48] ,n1649);
    nor g1976(n1551 ,n5[54] ,n1026);
    dff g1977(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n561), .Q(n7[28]));
    nand g1978(n1599 ,n606 ,n973);
    nand g1979(n2193 ,n2064 ,n2063);
    dff g1980(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n548), .Q(n8[10]));
    nand g1981(n2306 ,n1844 ,n2258);
    dff g1982(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2107), .Q(n4[52]));
    nor g1983(n1371 ,n4[36] ,n1040);
    nand g1984(n2220 ,n3[38] ,n1885);
    nor g1985(n1511 ,n3[15] ,n1019);
    nand g1986(n1139 ,n654 ,n874);
    nand g1987(n2039 ,n5[7] ,n1637);
    nand g1988(n2239 ,n3[19] ,n1872);
    nand g1989(n1724 ,n5[49] ,n1643);
    nand g1990(n1159 ,n720 ,n897);
    nor g1991(n249 ,n66 ,n248);
    nand g1992(n1184 ,n726 ,n928);
    nor g1993(n859 ,n435 ,n805);
    dff g1994(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2079), .Q(n4[16]));
    nor g1995(n877 ,n1 ,n808);
    nand g1996(n788 ,n8[6] ,n2[6]);
    or g1997(n1859 ,n1069 ,n1446);
    nand g1998(n1986 ,n4[53] ,n1462);
    nor g1999(n1368 ,n5[36] ,n1040);
    nor g2000(n491 ,n8[27] ,n2[59]);
    nor g2001(n1382 ,n5[33] ,n1038);
    nand g2002(n2025 ,n5[57] ,n1480);
    not g2003(n1665 ,n1580);
    not g2004(n1260 ,n1132);
    nand g2005(n1925 ,n5[19] ,n1633);
    nand g2006(n1078 ,n612 ,n813);
    nor g2007(n464 ,n8[17] ,n2[17]);
    nand g2008(n1016 ,n8[3] ,n877);
    nor g2009(n913 ,n405 ,n805);
    nand g2010(n2200 ,n3[58] ,n1865);
    dff g2011(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2317), .Q(n3[59]));
    not g2012(n1652 ,n1567);
    nor g2013(n390 ,n2355 ,n10[0]);
    nand g2014(n2153 ,n1819 ,n1818);
    not g2015(n1272 ,n1144);
    nor g2016(n26 ,n2[45] ,n2[109]);
    nor g2017(n836 ,n391 ,n804);
    nand g2018(n138 ,n73 ,n92);
    nor g2019(n1526 ,n3[17] ,n1021);
    nand g2020(n713 ,n8[23] ,n2[119]);
    nor g2021(n1845 ,n1407 ,n1242);
    nor g2022(n1403 ,n3[50] ,n1022);
    nor g2023(n969 ,n446 ,n875);
    dff g2024(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n536), .Q(n8[16]));
    nand g2025(n608 ,n8[12] ,n2335);
    nand g2026(n2305 ,n1846 ,n2211);
    nand g2027(n1081 ,n624 ,n926);
    nand g2028(n2152 ,n1815 ,n1813);
    nor g2029(n1358 ,n5[40] ,n1010);
    nor g2030(n583 ,n339 ,n1);
    nand g2031(n2413 ,n7[13] ,n7[12]);
    xnor g2032(n2363 ,n95 ,n215);
    nor g2033(n540 ,n327 ,n1);
    nand g2034(n782 ,n8[6] ,n2329);
    nor g2035(n590 ,n307 ,n1);
    not g2036(n293 ,n2[38]);
    not g2037(n1207 ,n1079);
    nor g2038(n1059 ,n8[23] ,n876);
    nor g2039(n520 ,n8[26] ,n2[90]);
    nor g2040(n1067 ,n8[30] ,n876);
    nand g2041(n2082 ,n1768 ,n1767);
    nor g2042(n405 ,n8[12] ,n2367);
    not g2043(n1247 ,n1119);
    or g2044(n1485 ,n810 ,n1047);
    nand g2045(n2102 ,n1976 ,n1975);
    not g2046(n1233 ,n1105);
    nand g2047(n1621 ,n759 ,n951);
    nor g2048(n61 ,n2[14] ,n2[78]);
    nand g2049(n1591 ,n632 ,n983);
    nand g2050(n1819 ,n5[34] ,n1489);
    nor g2051(n914 ,n442 ,n805);
    nand g2052(n671 ,n8[11] ,n2[43]);
    nor g2053(n53 ,n2[44] ,n2[108]);
    dff g2054(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2136), .Q(n5[46]));
    nand g2055(n2094 ,n1811 ,n1810);
    nor g2056(n232 ,n106 ,n231);
    nand g2057(n1079 ,n613 ,n913);
    nand g2058(n1076 ,n607 ,n827);
    nand g2059(n1124 ,n675 ,n858);
    nand g2060(n1130 ,n682 ,n865);
    nor g2061(n971 ,n478 ,n875);
    or g2062(n1872 ,n1054 ,n1446);
    xnor g2063(n96 ,n2[2] ,n2[66]);
    nor g2064(n1515 ,n5[11] ,n1014);
    nor g2065(n841 ,n394 ,n804);
    nor g2066(n469 ,n8[14] ,n2[14]);
    nand g2067(n1798 ,n4[5] ,n1470);
    nand g2068(n1033 ,n8[27] ,n877);
    nor g2069(n70 ,n2[4] ,n2[68]);
    nor g2070(n477 ,n8[28] ,n2[60]);
    nand g2071(n2121 ,n2034 ,n2033);
    nor g2072(n830 ,n387 ,n805);
    nand g2073(n609 ,n8[19] ,n2[51]);
    xnor g2074(n78 ,n2[45] ,n2[109]);
    nand g2075(n2284 ,n1952 ,n2252);
    nand g2076(n1038 ,n10[1] ,n877);
    nand g2077(n679 ,n8[11] ,n2[107]);
    nand g2078(n770 ,n8[16] ,n2371);
    nand g2079(n1183 ,n748 ,n814);
    not g2080(n1258 ,n1130);
    nand g2081(n1153 ,n714 ,n893);
    not g2082(n1698 ,n1613);
    or g2083(n1488 ,n807 ,n1066);
    or g2084(n1454 ,n810 ,n1061);
    nor g2085(n519 ,n8[16] ,n2[48]);
    dff g2086(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2309), .Q(n3[51]));
    nand g2087(n1192 ,n794 ,n933);
    nor g2088(n922 ,n498 ,n804);
    nand g2089(n2419 ,n2408 ,n2401);
    dff g2090(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2273), .Q(n3[17]));
    or g2091(n1869 ,n1058 ,n1446);
    not g2092(n1270 ,n1142);
    nor g2093(n953 ,n353 ,n269);
    not g2094(n1282 ,n1154);
    or g2095(n1487 ,n810 ,n1056);
    not g2096(n283 ,n2[27]);
    dff g2097(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n555), .Q(n8[9]));
    nor g2098(n965 ,n385 ,n875);
    nand g2099(n2286 ,n1956 ,n2254);
    nor g2100(n159 ,n64 ,n158);
    nor g2101(n1001 ,n495 ,n875);
    nand g2102(n2215 ,n3[43] ,n1880);
    nand g2103(n693 ,n8[6] ,n2[38]);
    nor g2104(n66 ,n2[56] ,n2[120]);
    nand g2105(n1125 ,n677 ,n861);
    nor g2106(n369 ,n2324 ,n10[1]);
    dff g2107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2120), .Q(n4[39]));
    nor g2108(n1922 ,n1330 ,n1280);
    nand g2109(n2219 ,n3[39] ,n1884);
    nor g2110(n917 ,n460 ,n267);
    not g2111(n802 ,n801);
    nor g2112(n911 ,n502 ,n804);
    nor g2113(n1331 ,n5[50] ,n1022);
    nor g2114(n1394 ,n5[30] ,n1013);
    nor g2115(n494 ,n8[27] ,n2[123]);
    dff g2116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2068), .Q(n4[27]));
    nand g2117(n2317 ,n1825 ,n2199);
    nor g2118(n219 ,n46 ,n218);
    nor g2119(n1437 ,n3[28] ,n1034);
    nor g2120(n1380 ,n3[62] ,n1013);
    nor g2121(n601 ,n316 ,n1);
    dff g2122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2133), .Q(n5[5]));
    xnor g2123(n2355 ,n88 ,n199);
    nor g2124(n556 ,n305 ,n1);
    not g2125(n1655 ,n1570);
    nand g2126(n1156 ,n717 ,n896);
    dff g2127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n537), .Q(n8[2]));
    not g2128(n1230 ,n1102);
    nand g2129(n2115 ,n2014 ,n2013);
    not g2130(n1672 ,n1587);
    nor g2131(n521 ,n8[17] ,n2372);
    dff g2132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2275), .Q(n3[15]));
    nand g2133(n1175 ,n659 ,n916);
    nor g2134(n567 ,n8[21] ,n2[21]);
    nand g2135(n1155 ,n716 ,n894);
    nor g2136(n1415 ,n3[43] ,n1014);
    not g2137(n1285 ,n1157);
    nor g2138(n394 ,n8[22] ,n2[54]);
    dff g2139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n546), .Q(n8[5]));
    dff g2140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2265), .Q(n3[25]));
    nor g2141(n1745 ,n1339 ,n1205);
    nand g2142(n698 ,n8[14] ,n2[110]);
    nand g2143(n634 ,n8[7] ,n2[71]);
    nor g2144(n1794 ,n1364 ,n1213);
    not g2145(n340 ,n2389);
    nor g2146(n817 ,n364 ,n805);
    not g2147(n305 ,n2[6]);
    nor g2148(n11 ,n2[47] ,n2[111]);
    nor g2149(n538 ,n309 ,n1);
    nor g2150(n962 ,n406 ,n269);
    nor g2151(n1728 ,n1540 ,n1654);
    nand g2152(n610 ,n8[15] ,n2370);
    nand g2153(n2264 ,n1916 ,n2232);
    nand g2154(n1032 ,n8[26] ,n877);
    nand g2155(n1615 ,n765 ,n957);
    xnor g2156(n135 ,n2[43] ,n2[107]);
    nor g2157(n496 ,n8[14] ,n2369);
    nor g2158(n1531 ,n4[22] ,n1026);
    nor g2159(n1497 ,n3[9] ,n1012);
    nand g2160(n2321 ,n1817 ,n2195);
    nand g2161(n1826 ,n5[32] ,n1457);
    nand g2162(n1944 ,n5[14] ,n1648);
    dff g2163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n602), .Q(n8[3]));
    nor g2164(n1517 ,n5[10] ,n1041);
    nor g2165(n1494 ,n5[14] ,n1018);
    nor g2166(n419 ,n8[24] ,n2[56]);
    nand g2167(n1190 ,n742 ,n934);
    nor g2168(n259 ,n37 ,n258);
    nor g2169(n554 ,n337 ,n1);
    nand g2170(n2100 ,n1972 ,n1970);
    nor g2171(n482 ,n8[2] ,n2[98]);
    nor g2172(n397 ,n8[12] ,n2[108]);
    not g2173(n1228 ,n1100);
    nor g2174(n1061 ,n8[25] ,n876);
    nor g2175(n930 ,n404 ,n805);
    nand g2176(n2229 ,n3[29] ,n1862);
    nand g2177(n1568 ,n775 ,n1005);
    nor g2178(n982 ,n363 ,n269);
    nand g2179(n1595 ,n676 ,n978);
    dff g2180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n564), .Q(n8[22]));
    nor g2181(n2425 ,n2416 ,n2421);
    not g2182(n1266 ,n1138);
    not g2183(n274 ,n2[25]);
    nand g2184(n2198 ,n3[60] ,n1863);
    dff g2185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2163), .Q(n5[24]));
    nor g2186(n1544 ,n4[26] ,n1032);
    nor g2187(n59 ,n2[43] ,n2[107]);
    dff g2188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2077), .Q(n4[18]));
    nor g2189(n1354 ,n4[61] ,n1035);
    nand g2190(n263 ,n6[1] ,n6[0]);
    nand g2191(n1169 ,n736 ,n908);
    not g2192(n291 ,n2[23]);
    nor g2193(n1985 ,n1506 ,n1689);
    nor g2194(n528 ,n8[15] ,n2[111]);
    nand g2195(n1014 ,n8[11] ,n877);
    nand g2196(n736 ,n8[11] ,n2[11]);
    nor g2197(n1395 ,n3[53] ,n1025);
    nor g2198(n1823 ,n1383 ,n1222);
    not g2199(n1219 ,n1091);
    or g2200(n2422 ,n2410 ,n2414);
    nor g2201(n454 ,n8[16] ,n2[112]);
    nand g2202(n1160 ,n723 ,n900);
    not g2203(n304 ,n2[59]);
    nor g2204(n1846 ,n1408 ,n1244);
    dff g2205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2071), .Q(n4[24]));
    nor g2206(n385 ,n8[18] ,n2[114]);
    nor g2207(n1407 ,n5[28] ,n1034);
    nor g2208(n867 ,n486 ,n805);
    nor g2209(n506 ,n8[7] ,n2[103]);
    nand g2210(n2285 ,n1954 ,n2253);
    nor g2211(n218 ,n126 ,n217);
    nor g2212(n261 ,n48 ,n260);
    dff g2213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2106), .Q(n4[53]));
    nor g2214(n1780 ,n1358 ,n1211);
    nor g2215(n173 ,n45 ,n172);
    nand g2216(n1036 ,n8[31] ,n877);
    not g2217(n1713 ,n1628);
    nand g2218(n1570 ,n766 ,n1003);
    nand g2219(n1127 ,n678 ,n859);
    nor g2220(n2022 ,n1496 ,n1701);
    nor g2221(n995 ,n443 ,n875);
    nand g2222(n1101 ,n649 ,n839);
    nand g2223(n1024 ,n8[20] ,n877);
    nand g2224(n1162 ,n724 ,n901);
    dff g2225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2262), .Q(n3[28]));
    nand g2226(n2052 ,n5[53] ,n1467);
    nand g2227(n734 ,n8[12] ,n2[12]);
    nor g2228(n1918 ,n1443 ,n1277);
    nand g2229(n1816 ,n4[0] ,n1455);
    nand g2230(n2144 ,n1776 ,n1773);
    nor g2231(n379 ,n8[29] ,n2[93]);
    nor g2232(n1550 ,n4[35] ,n1016);
    nand g2233(n746 ,n8[18] ,n2[82]);
    nand g2234(n764 ,n8[2] ,n2[2]);
    nand g2235(n1140 ,n757 ,n879);
    not g2236(n1314 ,n1186);
    nor g2237(n1907 ,n1432 ,n1268);
    nor g2238(n834 ,n491 ,n804);
    nor g2239(n200 ,n88 ,n199);
    xnor g2240(n127 ,n2[18] ,n2[82]);
    nand g2241(n2084 ,n1775 ,n1774);
    nor g2242(n1897 ,n1425 ,n1259);
    nor g2243(n565 ,n297 ,n1);
    nand g2244(n1616 ,n753 ,n956);
    xnor g2245(n95 ,n2[40] ,n2[104]);
    nor g2246(n1549 ,n3[20] ,n1024);
    dff g2247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2094), .Q(n4[1]));
    not g2248(n336 ,n2[13]);
    nor g2249(n542 ,n295 ,n1);
    nand g2250(n640 ,n2324 ,n10[1]);
    nor g2251(n855 ,n412 ,n804);
    nand g2252(n1610 ,n697 ,n963);
    nor g2253(n445 ,n8[12] ,n2[44]);
    dff g2254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2174), .Q(n5[13]));
    xnor g2255(n131 ,n2[42] ,n2[106]);
    not g2256(n797 ,n798);
    nor g2257(n398 ,n8[20] ,n2375);
    not g2258(n1704 ,n1619);
    nor g2259(n548 ,n333 ,n1);
    nor g2260(n1829 ,n1445 ,n1225);
    not g2261(n285 ,n2[24]);
    nor g2262(n246 ,n133 ,n245);
    nor g2263(n165 ,n61 ,n164);
    or g2264(n1876 ,n1049 ,n1446);
    nor g2265(n979 ,n400 ,n875);
    nor g2266(n151 ,n55 ,n150);
    dff g2267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2149), .Q(n5[37]));
    nor g2268(n409 ,n8[28] ,n2[92]);
    nor g2269(n50 ,n2[35] ,n2[99]);
    dff g2270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2296), .Q(n3[38]));
    nand g2271(n1629 ,n787 ,n1009);
    dff g2272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n582), .Q(n7[19]));
    nand g2273(n1117 ,n666 ,n852);
    dff g2274(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n545), .Q(n8[6]));
    nand g2275(n739 ,n8[10] ,n2[10]);
    nor g2276(n47 ,n2[19] ,n2[83]);
    nand g2277(n1738 ,n5[47] ,n1631);
    not g2278(n1301 ,n1173);
    nor g2279(n487 ,n8[3] ,n2326);
    nor g2280(n1722 ,n1333 ,n1323);
    nand g2281(n1765 ,n4[14] ,n1479);
    nor g2282(n2047 ,n1553 ,n1326);
    not g2283(n1675 ,n1590);
    nor g2284(n215 ,n38 ,n214);
    nor g2285(n51 ,n2[20] ,n2[84]);
    dff g2286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2078), .Q(n4[17]));
    nand g2287(n748 ,n8[3] ,n2326);
    not g2288(n569 ,n568);
    nor g2289(n1493 ,n3[10] ,n1041);
    not g2290(n1328 ,n1200);
    dff g2291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2118), .Q(n4[41]));
    xnor g2292(n89 ,n2[35] ,n2[99]);
    nor g2293(n857 ,n463 ,n804);
    nor g2294(n1767 ,n1430 ,n1665);
    nand g2295(n2123 ,n2041 ,n2040);
    nor g2296(n1387 ,n3[24] ,n1029);
    dff g2297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n598), .Q(n7[30]));
    nor g2298(n511 ,n8[13] ,n2368);
    nand g2299(n612 ,n8[13] ,n2368);
    nand g2300(n1198 ,n762 ,n937);
    xnor g2301(n2387 ,n6[3] ,n265);
    xnor g2302(n2347 ,n86 ,n183);
    not g2303(n1236 ,n1108);
    nor g2304(n1546 ,n4[39] ,n1030);
    nand g2305(n2428 ,n2417 ,n2427);
    dff g2306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2132), .Q(n5[49]));
    nand g2307(n1729 ,n4[24] ,n1456);
    nor g2308(n1558 ,n4[30] ,n1013);
    nand g2309(n665 ,n8[7] ,n2[103]);
    nand g2310(n1736 ,n4[22] ,n1460);
    not g2311(n1218 ,n1090);
    nor g2312(n1939 ,n1504 ,n1289);
    nor g2313(n341 ,n8[28] ,n2383);
    nor g2314(n422 ,n8[24] ,n2379);
    nor g2315(n1425 ,n3[36] ,n1040);
    nand g2316(n719 ,n8[19] ,n2[19]);
    nand g2317(n720 ,n8[17] ,n2340);
    nor g2318(n1055 ,n8[20] ,n876);
    nor g2319(n539 ,n311 ,n1);
    nand g2320(n625 ,n8[4] ,n2[68]);
    nor g2321(n365 ,n8[27] ,n2382);
    nand g2322(n1592 ,n633 ,n982);
    nor g2323(n533 ,n8[15] ,n2370);
    dff g2324(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2259), .Q(n3[31]));
    nand g2325(n752 ,n8[10] ,n2[42]);
    nor g2326(n434 ,n8[10] ,n2365);
    dff g2327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2092), .Q(n4[3]));
    not g2328(n268 ,n875);
    dff g2329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2067), .Q(n4[28]));
    nor g2330(n1381 ,n3[61] ,n1035);
    nand g2331(n2265 ,n1918 ,n2233);
    nand g2332(n2156 ,n1832 ,n1828);
    nor g2333(n255 ,n71 ,n254);
    nor g2334(n45 ,n2[18] ,n2[82]);
    nor g2335(n1350 ,n4[14] ,n1018);
    nor g2336(n356 ,n8[25] ,n2380);
    nand g2337(n2318 ,n1823 ,n2198);
    nand g2338(n2138 ,n1752 ,n1747);
    nand g2339(n691 ,n8[13] ,n2[77]);
    nand g2340(n1974 ,n4[58] ,n1451);
    dff g2341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2299), .Q(n3[41]));
    nor g2342(n1540 ,n4[24] ,n1029);
    nand g2343(n2020 ,n4[42] ,n1447);
    nand g2344(n2237 ,n3[21] ,n1870);
    nand g2345(n1609 ,n768 ,n980);
    or g2346(n1466 ,n807 ,n1068);
    or g2347(n1871 ,n1055 ,n1446);
    nand g2348(n1093 ,n626 ,n830);
    not g2349(n300 ,n2[63]);
    nand g2350(n2062 ,n4[29] ,n1632);
    nor g2351(n1353 ,n4[12] ,n1015);
    nand g2352(n766 ,n8[23] ,n2[87]);
    nor g2353(n1422 ,n3[38] ,n1011);
    nand g2354(n650 ,n8[23] ,n2[55]);
    nor g2355(n543 ,n336 ,n1);
    nor g2356(n257 ,n65 ,n256);
    nor g2357(n1507 ,n3[5] ,n1039);
    nor g2358(n584 ,n291 ,n1);
    dff g2359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2286), .Q(n3[4]));
    nor g2360(n1356 ,n4[60] ,n1034);
    xnor g2361(n130 ,n2[20] ,n2[84]);
    nor g2362(n868 ,n441 ,n271);
    nor g2363(n1337 ,n5[47] ,n1019);
    nor g2364(n492 ,n2[96] ,n10[0]);
    xnor g2365(n113 ,n2[61] ,n2[125]);
    nor g2366(n947 ,n484 ,n875);
    not g2367(n295 ,n2[62]);
    nor g2368(n1367 ,n5[37] ,n1039);
    not g2369(n279 ,n2[12]);
    nand g2370(n2089 ,n1793 ,n1792);
    nand g2371(n1788 ,n5[39] ,n1637);
    nor g2372(n497 ,n2[97] ,n10[1]);
    dff g2373(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2086), .Q(n4[9]));
    nand g2374(n765 ,n8[10] ,n2[106]);
    dff g2375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n554), .Q(n7[17]));
    nor g2376(n1926 ,n1555 ,n1283);
    dff g2377(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2261), .Q(n3[29]));
    nor g2378(n1333 ,n5[49] ,n1021);
    nor g2379(n427 ,n8[5] ,n2[37]);
    not g2380(n1273 ,n1145);
    nand g2381(n1179 ,n643 ,n922);
    nand g2382(n809 ,n273 ,n801);
    nor g2383(n1050 ,n8[16] ,n876);
    not g2384(n1681 ,n1596);
    nand g2385(n1809 ,n5[36] ,n1642);
    nand g2386(n778 ,n8[17] ,n2372);
    xnor g2387(n2329 ,n136 ,n147);
    dff g2388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2171), .Q(n5[16]));
    nand g2389(n2243 ,n3[15] ,n1876);
    nand g2390(n1013 ,n8[30] ,n877);
    nor g2391(n483 ,n8[4] ,n2[68]);
    nand g2392(n742 ,n8[4] ,n2327);
    dff g2393(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n587), .Q(n7[29]));
    nor g2394(n1411 ,n5[27] ,n1033);
    nand g2395(n1754 ,n4[17] ,n1473);
    nand g2396(n670 ,n8[11] ,n2[75]);
    nand g2397(n621 ,n8[5] ,n2360);
    nor g2398(n2026 ,n1442 ,n1702);
    nor g2399(n1946 ,n1493 ,n1298);
    nor g2400(n1068 ,n10[1] ,n876);
    nand g2401(n636 ,n2[64] ,n10[0]);
    not g2402(n325 ,n2[39]);
    not g2403(n286 ,n2[33]);
    xnor g2404(n2388 ,n6[2] ,n263);
    dff g2405(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n547), .Q(n8[8]));
    nor g2406(n853 ,n366 ,n271);
    nand g2407(n702 ,n8[27] ,n2[27]);
    nand g2408(n1790 ,n4[7] ,n1459);
    nand g2409(n2238 ,n3[20] ,n1871);
    dff g2410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2137), .Q(n5[4]));
    nor g2411(n499 ,n8[21] ,n2376);
    dff g2412(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2151), .Q(n5[36]));
    nand g2413(n2117 ,n2020 ,n2019);
    not g2414(n1222 ,n1094);
    nor g2415(n522 ,n8[6] ,n2329);
    nor g2416(n1564 ,n4[28] ,n1034);
    not g2417(n1653 ,n1568);
    dff g2418(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n552), .Q(n8[12]));
    nor g2419(n1820 ,n1380 ,n1218);
    nand g2420(n651 ,n8[12] ,n2[44]);
    dff g2421(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2135), .Q(n5[47]));
    dff g2422(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n540), .Q(n7[31]));
    nor g2423(n1048 ,n8[14] ,n876);
    nor g2424(n38 ,n2[39] ,n2[103]);
    nor g2425(n462 ,n8[17] ,n2340);
    nand g2426(n2322 ,n1935 ,n2242);
    nor g2427(n2404 ,n2397 ,n7[26]);
    nand g2428(n1579 ,n701 ,n995);
    nor g2429(n358 ,n8[20] ,n2[52]);
    nand g2430(n2236 ,n3[22] ,n1869);
    nor g2431(n21 ,n2[34] ,n2[98]);
    nor g2432(n460 ,n8[7] ,n2330);
    nor g2433(n16 ,n2[16] ,n2[80]);
    nor g2434(n1436 ,n5[21] ,n1025);
    nor g2435(n220 ,n131 ,n219);
    xnor g2436(n2359 ,n108 ,n207);
    nor g2437(n363 ,n2[65] ,n10[1]);
    dff g2438(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n380), .Q(n6[0]));
    nand g2439(n762 ,n8[21] ,n2376);
    or g2440(n1879 ,n1046 ,n1446);
    nor g2441(n212 ,n116 ,n211);
    nor g2442(n858 ,n410 ,n804);
    nor g2443(n1769 ,n1351 ,n1265);
    nor g2444(n1821 ,n1381 ,n1220);
    xnor g2445(n2384 ,n113 ,n257);
    nand g2446(n2415 ,n2404 ,n2412);
    nand g2447(n1026 ,n8[22] ,n877);
    nor g2448(n348 ,n8[29] ,n2352);
    dff g2449(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2160), .Q(n5[27]));
    nor g2450(n46 ,n2[41] ,n2[105]);
    nand g2451(n1571 ,n760 ,n1002);
    nand g2452(n1080 ,n708 ,n815);
    nor g2453(n1501 ,n3[7] ,n1030);
    nand g2454(n726 ,n2[0] ,n10[0]);
    nor g2455(n571 ,n306 ,n1);
    nor g2456(n440 ,n8[27] ,n2[27]);
    xnor g2457(n97 ,n2[33] ,n2[97]);
    or g2458(n1449 ,n807 ,n1044);
    nand g2459(n1623 ,n774 ,n961);
    nand g2460(n1037 ,n10[0] ,n877);
    not g2461(n280 ,n2[44]);
    or g2462(n1465 ,n807 ,n1058);
    nor g2463(n1831 ,n1391 ,n1229);
    nor g2464(n400 ,n8[31] ,n2[127]);
    nand g2465(n2275 ,n1937 ,n2243);
    nand g2466(n1977 ,n4[56] ,n1456);
    nand g2467(n1930 ,n5[18] ,n1638);
    nor g2468(n2033 ,n1370 ,n1704);
    nand g2469(n2303 ,n1849 ,n2213);
    nor g2470(n537 ,n318 ,n1);
    nor g2471(n362 ,n8[25] ,n2[121]);
    nor g2472(n1363 ,n4[6] ,n1011);
    nor g2473(n823 ,n351 ,n805);
    nor g2474(n2045 ,n1551 ,n1322);
    nand g2475(n2110 ,n2000 ,n1999);
    nor g2476(n1397 ,n4[43] ,n1014);
    xnor g2477(n2367 ,n84 ,n223);
    nor g2478(n994 ,n367 ,n875);
    nand g2479(n2142 ,n1777 ,n1766);
    nand g2480(n2080 ,n1761 ,n1760);
    nor g2481(n501 ,n8[7] ,n2[7]);
    not g2482(n1670 ,n1585);
    nor g2483(n1757 ,n1348 ,n1662);
    dff g2484(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2081), .Q(n4[14]));
    xnor g2485(n104 ,n2[5] ,n2[69]);
    nor g2486(n934 ,n458 ,n267);
    nand g2487(n2258 ,n3[48] ,n1875);
    nor g2488(n193 ,n49 ,n192);
    nor g2489(n1512 ,n3[3] ,n1016);
    nor g2490(n839 ,n419 ,n271);
    nor g2491(n568 ,n9[0] ,n1);
    nor g2492(n1508 ,n5[12] ,n1015);
    nand g2493(n2176 ,n1969 ,n1963);
    nor g2494(n24 ,n2[49] ,n2[113]);
    nor g2495(n840 ,n473 ,n271);
    or g2496(n10[1] ,n8[1] ,n2429);
    nor g2497(n950 ,n524 ,n875);
    nand g2498(n743 ,n8[28] ,n2[60]);
    xnor g2499(n90 ,n2[62] ,n2[126]);
    nor g2500(n935 ,n422 ,n267);
    dff g2501(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2279), .Q(n3[11]));
    dff g2502(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2096), .Q(n4[63]));
    nor g2503(n170 ,n124 ,n169);
    or g2504(n1448 ,n807 ,n1064);
    nand g2505(n1573 ,n751 ,n974);
    nand g2506(n1199 ,n785 ,n938);
    nand g2507(n714 ,n8[22] ,n2[22]);
    nor g2508(n1954 ,n1507 ,n1305);
    nor g2509(n229 ,n56 ,n228);
    nor g2510(n163 ,n34 ,n162);
    nand g2511(n1116 ,n664 ,n851);
    nor g2512(n800 ,n9[1] ,n797);
    nand g2513(n1112 ,n603 ,n929);
    nor g2514(n976 ,n461 ,n875);
    nor g2515(n260 ,n90 ,n259);
    nand g2516(n2067 ,n1978 ,n2065);
    nand g2517(n1102 ,n650 ,n840);
    dff g2518(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2267), .Q(n3[23]));
    nor g2519(n1822 ,n1382 ,n1221);
    nor g2520(n157 ,n29 ,n156);
    nor g2521(n1949 ,n1499 ,n1301);
    dff g2522(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n558), .Q(n7[9]));
    nand g2523(n1812 ,n4[39] ,n1459);
    nor g2524(n433 ,n2[1] ,n10[1]);
    or g2525(n1882 ,n1051 ,n1446);
    not g2526(n1657 ,n1572);
    nand g2527(n725 ,n8[16] ,n2339);
    dff g2528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2321), .Q(n3[63]));
    nand g2529(n2277 ,n1938 ,n2244);
    nand g2530(n722 ,n8[16] ,n2[80]);
    nand g2531(n647 ,n8[31] ,n2354);
    or g2532(n1467 ,n807 ,n1073);
    dff g2533(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2300), .Q(n3[42]));
    nand g2534(n1585 ,n642 ,n989);
    nor g2535(n874 ,n429 ,n804);
    not g2536(n1302 ,n1174);
    nand g2537(n741 ,n8[24] ,n2[120]);
    nand g2538(n683 ,n8[24] ,n2347);
    not g2539(n1299 ,n1171);
    nor g2540(n40 ,n2[25] ,n2[89]);
    not g2541(n1658 ,n1573);
    dff g2542(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2184), .Q(n5[59]));
    nor g2543(n1789 ,n1373 ,n1671);
    nor g2544(n182 ,n137 ,n181);
    nand g2545(n1718 ,n4[27] ,n1450);
    nor g2546(n901 ,n466 ,n804);
    nand g2547(n1173 ,n700 ,n915);
    nand g2548(n771 ,n8[14] ,n2369);
    nor g2549(n1743 ,n1519 ,n1658);
    nor g2550(n1755 ,n1347 ,n1207);
    xnor g2551(n120 ,n2[39] ,n2[103]);
    dff g2552(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n589), .Q(n7[0]));
    xnor g2553(n2331 ,n125 ,n151);
    not g2554(n303 ,n2[7]);
    nor g2555(n391 ,n8[26] ,n2[58]);
    nor g2556(n346 ,n8[2] ,n2357);
    nand g2557(n2282 ,n1949 ,n2250);
    or g2558(n1640 ,n807 ,n1051);
    nand g2559(n1900 ,n5[24] ,n1461);
    nand g2560(n777 ,n8[7] ,n2330);
    xnor g2561(n2366 ,n135 ,n221);
    or g2562(n1486 ,n810 ,n1070);
    nand g2563(n1022 ,n8[18] ,n877);
    nand g2564(n1040 ,n8[4] ,n877);
    nor g2565(n991 ,n402 ,n875);
    nand g2566(n2320 ,n1820 ,n2196);
    dff g2567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2148), .Q(n5[38]));
    dff g2568(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n573), .Q(n8[27]));
    nand g2569(n682 ,n8[5] ,n2[37]);
    xnor g2570(n2373 ,n109 ,n235);
    nand g2571(n2032 ,n5[56] ,n1461);
    nand g2572(n721 ,n8[18] ,n2[18]);
    nand g2573(n1588 ,n622 ,n986);
    nor g2574(n1996 ,n1509 ,n1692);
    xnor g2575(n100 ,n2[59] ,n2[123]);
    nor g2576(n357 ,n8[2] ,n2[66]);
    nor g2577(n1057 ,n8[4] ,n876);
    not g2578(n322 ,n2[50]);
    nor g2579(n251 ,n33 ,n250);
    nor g2580(n842 ,n375 ,n805);
    nor g2581(n1813 ,n1375 ,n1216);
    nor g2582(n1525 ,n3[16] ,n1020);
    nor g2583(n1971 ,n1517 ,n1313);
    not g2584(n314 ,n2[45]);
    not g2585(n1687 ,n1602);
    xnor g2586(n2381 ,n122 ,n251);
    nor g2587(n1748 ,n1342 ,n1659);
    nor g2588(n1419 ,n5[25] ,n1031);
    nor g2589(n816 ,n358 ,n804);
    nor g2590(n360 ,n8[14] ,n2337);
    nor g2591(n383 ,n8[30] ,n2[30]);
    nor g2592(n1894 ,n1422 ,n1256);
    nor g2593(n1418 ,n3[41] ,n1012);
    nand g2594(n1177 ,n689 ,n920);
    nor g2595(n927 ,n350 ,n267);
    nand g2596(n1187 ,n646 ,n864);
    nand g2597(n2003 ,n5[9] ,n1640);
    nor g2598(n1335 ,n5[48] ,n1020);
    dff g2599(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2142), .Q(n5[2]));
    or g2600(n1463 ,n807 ,n1059);
    nand g2601(n2278 ,n1942 ,n2246);
    nand g2602(n1740 ,n5[4] ,n1642);
    nor g2603(n1771 ,n1353 ,n1666);
    or g2604(n1641 ,n807 ,n1045);
    nor g2605(n546 ,n276 ,n1);
    nor g2606(n478 ,n8[24] ,n2[120]);
    nand g2607(n1141 ,n690 ,n873);
    dff g2608(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2085), .Q(n4[10]));
    nor g2609(n1903 ,n1429 ,n1266);
    nor g2610(n149 ,n23 ,n148);
    nor g2611(n2399 ,n7[11] ,n7[10]);
    dff g2612(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n565), .Q(n7[3]));
    nand g2613(n2304 ,n1847 ,n2212);
    nand g2614(n678 ,n8[25] ,n2348);
    nor g2615(n233 ,n17 ,n232);
    nor g2616(n1046 ,n8[12] ,n876);
    nand g2617(n681 ,n8[18] ,n2[114]);
    nor g2618(n597 ,n283 ,n1);
    not g2619(n1232 ,n1104);
    nor g2620(n1346 ,n4[17] ,n1021);
    xnor g2621(n87 ,n2[25] ,n2[89]);
    or g2622(n1490 ,n810 ,n1068);
    nor g2623(n248 ,n93 ,n247);
    nor g2624(n978 ,n488 ,n269);
    nor g2625(n187 ,n40 ,n186);
    nor g2626(n1443 ,n3[25] ,n1031);
    nor g2627(n408 ,n8[6] ,n2[70]);
    nand g2628(n1108 ,n609 ,n845);
    nor g2629(n870 ,n421 ,n805);
    nor g2630(n1072 ,n8[3] ,n876);
    nor g2631(n576 ,n315 ,n1);
    nor g2632(n1950 ,n1501 ,n1303);
    dff g2633(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2129), .Q(n4[30]));
    not g2634(n324 ,n2[48]);
    nand g2635(n1171 ,n737 ,n909);
    nand g2636(n792 ,n8[17] ,n2[49]);
    nor g2637(n1933 ,n1532 ,n1287);
    dff g2638(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n577), .Q(n8[24]));
    nand g2639(n1941 ,n5[16] ,n1649);
    nor g2640(n515 ,n8[25] ,n2[89]);
    nand g2641(n2072 ,n1733 ,n1732);
    nand g2642(n619 ,n2323 ,n10[0]);
    nor g2643(n152 ,n125 ,n151);
    not g2644(n1283 ,n1155);
    nand g2645(n1181 ,n728 ,n924);
    nor g2646(n824 ,n377 ,n805);
    nand g2647(n1988 ,n5[63] ,n1449);
    nor g2648(n1064 ,n8[27] ,n876);
    nor g2649(n1802 ,n1369 ,n1675);
    or g2650(n1646 ,n807 ,n1047);
    nor g2651(n1336 ,n4[23] ,n1028);
    nor g2652(n1049 ,n8[15] ,n876);
    dff g2653(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2116), .Q(n4[43]));
    nor g2654(n530 ,n8[19] ,n2374);
    nor g2655(n2411 ,n2394 ,n7[17]);
    nor g2656(n20 ,n2[40] ,n2[104]);
    not g2657(n1215 ,n1087);
    nor g2658(n1432 ,n3[31] ,n1036);
    nand g2659(n2001 ,n5[61] ,n1488);
    nand g2660(n685 ,n8[3] ,n2[35]);
    nor g2661(n2005 ,n1536 ,n1262);
    nor g2662(n37 ,n2[61] ,n2[125]);
    dff g2663(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2189), .Q(n5[55]));
    nor g2664(n245 ,n32 ,n244);
    nand g2665(n1015 ,n8[12] ,n877);
    not g2666(n277 ,n2[55]);
    nor g2667(n172 ,n127 ,n171);
    not g2668(n1261 ,n1133);
    nor g2669(n2406 ,n7[9] ,n7[8]);
    nor g2670(n33 ,n2[57] ,n2[121]);
    xnor g2671(n74 ,n2[63] ,n2[127]);
    nor g2672(n1390 ,n5[31] ,n1036);
    nor g2673(n1959 ,n1513 ,n1679);
    nor g2674(n1787 ,n1360 ,n1219);
    nand g2675(n1082 ,n764 ,n826);
    dff g2676(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n593), .Q(n7[26]));
    nand g2677(n1029 ,n8[24] ,n877);
    nand g2678(n2131 ,n1715 ,n1717);
    not g2679(n1205 ,n1077);
    nand g2680(n667 ,n8[17] ,n2[113]);
    nor g2681(n820 ,n372 ,n805);
    nor g2682(n153 ,n25 ,n152);
endmodule
